��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~%���4������ҝ�?$����S�zܟGd�<�٠s]����[� ۙ`���J�շo��(P��?
=-5���R,6܀�w�e��qKd'Em��;��~�'8�M��G�Q�	Acr�q���Q~��]���h �ϰh��&}D=8�#��IO��p��m�����4���4V W�R���1�(�ո� ����R�V5X*3b���j˥`c\��dy�]M͝��vB�?���ܻ�uVe��u�@�E?����c(����U>Э����ءtp��X�ō����T;�
{�2�m�h�(�Hԡ({�Z��E���g��1��j]{oG#�N�����%��јV�d�A9��9{u����M>�s�b���C) ����/��G��&���=��QQc¦��wC�I�����lȹz:-3Կt�cO��M����I��h��t����&�Z���d���(�<M(gV���R�%�� ���=陌���ȆK#�.\�!D]����F�����%$��mB�x�ԯB���\)%�c�U�g��>#�?v�20�o���<|3�״>u��?N ��$���H�&�?�DGS����itp���s��$����:Ēzy�C4)����"A
�).l#0s�+��G�1�1��p�֗��`������������!ę�Ҁ�=v7b;~���!-���#��lnV��(��$�܃"�n��a�s_�,�!���:r�8��.fVc���l�������SF' a����3�%VZMh�)�$��,K�ܾ���K���B������X��8���G���.��� �y�O��˥m�ޒ(h���FM��W�o���X�BG�/�r�@��,)-��Z^;� n&��S3��vf�x��ݟ�Y@ذi�MܿfQ�N����7�.n�m��x;���MC�R�#P`k�Mg%���w�5�-�v�����?dM����`�Z��gr�G7r�J������i�܁��A�ۻ��*�cҰ��Io��	������4�jG-�y$!8��e���TBN�	���U���l�L�uv��X���x��%G�y=�9fb���C,l���������t9.[���K�w�"wC�:�Hr����q䮖����2+քL\�*M2�4ž��::c��8h�����H*�Lk̠�9��,�D���m����*Ȩ#	d��Q* �rWU��H�s��e�uo�j��nhrޚ�<S֠�D�f���T�D��@�֢���0`����cV��<.帤�=}+,��`�	����=]N����ʕh�������2!j���<����}��D��&����=7W������������"��5Y�V���k�H�;�I�:�~���n��s��X	ϝcu���c�Y��ؙ�ض�	��ǯ[��^x��`�+8��G6�K&>�)bJ�����t�}�`ڣ�m��+7ca$sD#��X>�8���8���ʦ-�&Gz��	�|��o|"��T��fb9�?�jC�����c���e�����l�K͑�J�`��	K#�v��Ԓ����0�FVnQ�)K�+lQ��n� ���ƶh�h6�8~(R1b� aM�r���~	$�'L�7��tWm�v�;��n�,~���lK��Y��?�z�V{דn���Z�K�b�O1�}�k~�"];��C|��c?<�JY�%��2�BT�@:U"����y$�
%ېu{���2�|���u]VUר���N�FXQu.���ܪā_`.sT�{�ݕPX�+l������F��]kvD܂Z(����|� �/�5%�&���R��'��ې�)O�ֈ����L�j|��ch�G4�%��7St��`6]|���������gЈ�/��w��C4�{�0c�5^e~��ė��y@���H�$��͙I/��I�y��TB��lDƢw4�h�'�A>�ܞ%|!$�α���ֱJ�s�BU���j޶`n�����(`�A��i�Uu���)W;�*�jMӧI;�	enx{�BВボ��.�}"��đa�e���O��1(`�L�|��N!Eyx�0��%����ן��f}���đ��g����~����@
{����h�c:d�,�MIN;-���@����9�5i���<��dxD���k�LN\z�'��A��z����gk#�q[꓎��X\�#�;i!3{3/�z�&�H���R��S*)=�	��/1�Q�g�f�P}���ȩ�ZZh\ז��M ������j�ey+Vn�D�N��.� /LQ _���ް*Zq���)��;%3�Q>;4-l܂��R�O���w��a[��sq5 y����J����ʽ��/J��	Fz\Ve����n��|һ�����8e9�����p=��:��մ=|SC�2^/ەI
~��zU�����?�F=)7�2{���z��H<��M��&�����eOkQ���RI���4�ئ���l*�2��'�&>���P5n�Y��1�4L�4^��r�� �ƊWnb��_�Vx�qq�mD�kG�
"��3|���q���7�5j��}���-:���������)���`V�!Ì�SjU��DV��?��W�P�a��9��~w�L#�Ů���RhƖRw��Ƚ�������Ȩ�� ���Cy�2ʫ{Rk���Nb�F�?kL�R�k�*���&LԥN����Ӧ�x�	����>�1�\w��I��
��u�U?����������fy�9�
���=
ԅ�i�W�4��8U��1yG�`�_�\�2 ��&G=ֺ`��sF��yNB�c�$�KN!RH��)��J��^<���k�齨��7|VB�ࡨK��v|"zA8����{_�Tp25�&~�����c����/�2�ZX�
H&�a�u^{����vV����t���:=i����rZpZ��� Pʿ|J�����\���0te�Ku/��4�y܏�偷5��q_�{EmW-Q�rNR_ҪC���&��b��C������sow�j�6�
��A�ܽж�3:k��{��xMax���_k'#υ�0�|����w��;���!�NH��e�jYbw�-���4y�;-��X��7��W%P�����W[�!QIym%�"��'LВ�n�	]���Ϳr��4i�{����%����"�d����� 4�ކ����g�,eA뼕/>z�ֲ�:	�O��x�\��EG��!7�^���@�L^rus�`���c�:KKU 3�!����RŻ%5�7Ŝ���yx!��A3��j;\���t�+)O�da����&��T����T��E2��yĒ.DŭNj��6��V�OV�&�Q�iB��BV�
[�nyv��sx�/W�����(��J�vH��@���5������o	��Y�m?G��`��U��K=��h��8q>ҏ�5N�KX:�ԣ��Ys(��	�����4�D�N�ŗH��d�R#����ZƤ��'J�GbA��+������cC���q|t^}�?߭�j����{W��t�1�ހј�T�}�Ho6'":! ��8�ʹ�˖d+A,����y�`�i�W���F��\؂�c�[���h�}���Z@�h,�@���3:�)��H���\
֓H?�Ι���4��"32�q	��3�� 3:�D+�^��fk3[�nMC_����pX%��Q��:���H���u�(�]���e۵�4���҂L7��I�_�ng���Y�T���½�*�q��PQ�F�����t4��˙���B���� �x<"«Ґ�k��@����V�5��o��Zf���~i,��
��9���"P�i�>j	z�qT8�+���B���h�����#r����h}����Kׯ�S����hM|�pG�/4Ә��R�t���N���G}uJ)ފSX�)�20���6.Z����yM�,����F\�	�	��@��S]|�}�ш�+��ρȜ��[�%�3Ӱ38,�7�r�Q}�����6��]c Id6G.���N���#s��x�����C�Ќ�/���%4��+	���-ZX�OGA�2�a�cT:tNG���j��zΔ�п���+a9�V"ʐ~x��\Cֵi�z�c6�5��=>P����.&����S0d�^g�Da������;�	W�WVz�P �X� ��W��{�z/�qÑ3��ؙ�"�K"_(�B�@��͉db��Q�G��/��6����)����'R�1������X��^�mD�)C���>��� ��_i�}ێ�0nRy��D@� �cRl/~�v����)�?Zf�sd�����1��Gҏ�פ?���&@�Mꮬ�I����_Dr�<})Β�.�c<�Tl�|?� Dpq�؜�CM$P�=cTh��z����Ɨ4�	�����Qq�j��D9O�H�q¢^A�ˁ��;Hf�!��֌��5+�Ă�s"�5M�2N�lBU��yߦ�^C_*����憭�S?T�ؔ��<�
g��k����|+�;%hK�9�ju|h�])�X�\#�K	H[�1�/�D�%ѫ2��+EA��i�pn�C�@��'��s�w����5Aϐ*�7�nԜ��&�dj�ˁ�S��y�E쭭�}�IqEN�5=�zW�`!{tJ�H%��{�/�L{���d��R���Y��wV�K�HS��� [r�ĕ��c�M��K�+w�G����C��_b�QLmD�~��@ܢ,3
8��t���h��T�����
O*���vA�B������B��N���o���������9<_!��7<l�脫�Ԑ�AQ5�]��'S�ȍ~7D���~p7=��-:M#:�8�w�{ʍ��aa�D������b� b!>�uv"���}Nٝ���SЦ��މW������A�UH]�Sa�l uɄo&@.���Z^3W���1���UY��=��wkI��wG�N����Fh��K[����^���Fnkc��F��D�� �E
��Z�:o�?YP�j*�W�YԱÂ0��|+�b`3970ޛ�ǹ�:3J��U#uN7;1�n�Of��μ"�Q���٘B�7S<!%N�����֣�kb���X�^4$��䙛c(0�#�p�����u�z�3vu�Zۆ2����#1r��P�XJK���8:.��h�zl�.?�~�#L�WA��&7��ģ���
�7H�
�$:�t�n8�G˩ϯ�,B���k+��B��-`��o�`���
m�#=�(���CS?���FR`-T��sGi�`�t���GN7a��lT����ȕwc?��e��1�Bу;��`!��/%ۮ+�F߫�_5������]A�}.�QL�u7�w�R�m�)rD�-5e	g
�@7��-�I�_U��{�|!`j%�F��p�L�bg�\z�䭣t�����Vb7�<�Ӏŋ�閶 n2���u�-7�棗���e�B�y�B�Q'�"ۢ���f)Btߴ̐]�Q9xBw@ �;�$̂��>�����0���r��|�:�hǼ���"��%��MӯD�~#_F�{z��]"&hG��Y~��#9F����g!a��#է�V����2VA�&/n��^WYeza�b2fLV~���h�i�P��^9	�׽g��5R��H���k�9-��k�3��BJ�)�o�Moeӌ�A�9]#�L�I<(�W�H*�`�i���sU(�t�[o;���u�<R��Ō��i�fϥ[�"��`���i���%K��H�L����<bfu�ݚ�+�k�+KJ�����u��hr�R�:Ϝ�����K*�lĤk�~BG�yøW#����C��E�oSk4_I����uD�����e򄳯�������~��Y�rY�x��b�l������s[e�7{�Y�4M�~?,u��MEv�&�P�6��ߵH�}��!��=��PG��(fKB|/m5��de[�2)�_B��/�d��~�7�[���̈́Ɍ)5l4���,��y���(l�E���74�Y�n=uQB�����(��c�G�~�VGa� _��G���$��Fp�F:��X��1}x-)V�XS�v�Z�C�#-��Y�9�m9K��5�؜�,����	JUp�"����+�
�2_��뫧N�[�L.�:�ĵ�G���2zu�d?���q�) d8��z�F*����6�c���8��������ß���sSw��#�lC��l'~���h���dl����k���6@�h�����O��1��ȝӶx�
��x���|��e��BHmrp��.����n���Ӓ;q͙���|��
���p�ő����>.�M�_a�d�:�
e�YS36c�HY=E�܃��u�0@��9^�(T��/�]��<ֵ�����᏶3��#��ɮ��R̓�?�1��U8`QFN嗰V3c�B�!�r���9�������?1f-{#�+�F���BuD��$��Z�[=����=t��*_�	�A����w6��xB#=�KѫxU��v"F2׍^��7�csE���ӭ{>
��*x��I@TI�n�}ծ+b�f9+Ok��%3�ӓ=�Ѷ�p�nU<��+��ju3���ޙ�&Wլ��s�wiJ���5�b��p�s������~S>�C�u��yQ��?۸�do_�ͭ�C�,���@���1�4�F���Eo�b�/�ԏ�������7��5.��]�T{{���J������y�Aϑ��Q�qY
�)�bg�:B�CX*@lS��TeN�F;7���� ��0)�۳'|n�<�2CYda7�V9�*=WasY$V@J.��`�u��3�z�0-x�λ��7~��#�Ke����6t��	�����dz�,�I��F	�|������q������� Hy����9QȞ�m�b��8�a�D~��čw�	��Wրk1V�<����dÍ��c�Ύ�k��`{�}  |�$��U3�� [�&.ؑ��*b9����w�k�xY4yJsDU��γK��rsx�Q�����T\f���f<�hǗ$n����V����)���\����� Gp!=�r�{U�C�5�����W���k3m�\Au��(��mp|�?��=G�u�n�-^��+o��� 6�������!��Y��3��1���;֮ۓt��y�:V�$͔r�@#�L�%�%�F��
��:	=�?m+��Z�����: ����p<���&�G̳/*.��j��E�Lߟk�%�ˊ��6?�DsCi(&[7��K�/Kn�V�fa�w��a@;�� �+�tP�$�h�6�n��>��e��,��l�X��I��8e���94a�������rv�/��7�pw�d�>K�}��}��2�0;�����~��y۠-���[A*���_������^�N)�<�о�+�;ܾ�ϳ�˚'{���Y�k��U�\������x�*�EU� S=b��jqg�ļpǚa�?PM	fZL��e�D��&�`2�yo�-��<���������w��va�#�n��KDlM����*HJ��q-���dNG-���9ZA��J�.��ˤl���ň���f�
u�Ci&��)�:�@�΄���~�|��ᎍ:��V�7��lS8�
+��~�����[+}-��{ y�C\�vKԹt�d?�>����D������=z���6��.��}Yy,��Qdܤ�d��Tr��|����X�}:p��f�M;��~A#���e�����\a7s��e�#���w�L�h��3+z���%����!�j��N2,�����w'%^�#2�d��aZ󘨚�oa�=G1U�CZ��v���tCWk��F��m�TR�������s����S���R���|�&�j�XD�$�N�26amW��=��V��S�Ď�=��gz��YE��[`m�R���xfU}���:Q�a�}�F�ǩ��'�Lx�l�?�Q���m�	��9���1��W��5�̑q�}���i�1��LRT�Y�{i����v���'q�E�\�?ٜ��ϪI|I���a��!5�ɦ1sk��UB�X4}�b_���E�.V�hbp�����`�� %/� �
`�����xlL#�+�(�"������Fp���k�x[�n��7>�Zb �D>�/�r��ι!�&`�	T#�-(Q2t����%���H`c���Il<Rj71T�uG��|���J�8VϜ��/V!��@�F&���|����{ܥ��n���:�&G��(�;�{���N�<�F*��cJi����y���ޙ홃���8�����#�A��H����C�<x�����ڐ��}�/�� �M��_3�KH>����O���#,��M�O�ap �x� 2�b]��r�,0���Uu�	�[�Ǚփ���՜�K21�p�L5Q����մf��F�4�b-�pL$���-Q���_�!��BBix����/s��g͌��3/"7d����ї��S�/��1� �%�Tm�B����3��-���[�gz9��L�NhEڢ4}n:��`R������
�0�+��b�"g[E*ܮ$y>��+������*ɤ��c?i���D��|����$��\�Uz�|T/��|-�[R��e"P~��kiʚb /�ѥt�g�9��3l+�`u���?1�_�����q\���ǐ��q����a�0#b	�o��23u��]jݰ��3Ԙ��.��b��QL��TlS�Y�����KB�Zn��X|�qo��%��Q&V:F�09/�5E76��G����qd���x�N��@ír���xkh�Q��Ge��Ť;�G�(g�x���������4~�T�ϝ���sT�z�cN��D���'?=�l��h����d�f ���66�E�A1%ҽ��R�qS��Q�U2�	;����}]�~���՜�C~/^�˸�:��GX�D[b�� 𥣪M���kL��E�~Yź�����+�F�2��ur��/�ҨH˰��ݸ�7k�gp�#��]U�^/e�Z�T���/(��4�.�d�9�x�����U�4��H�-��{�{8�v�B�B���yq�����?rAHdq�zi�^�	���.#��� ��b�\^\A?|0i@o��ܜqE�\k�®�ٲ�1=`h�[�L��>JǷí�^��H�y\��l`�'<�]��C���1;sX�=i�i����#���%L��o�ޮ��n�jN���`۴�M8�RD�d��	���$�ɇ/�񌿂d�7��$���A����`s!���Ք��r[�p��7��*�dﰝm�&"jש��]���hTf���VX��������Ȟ��R�:�"���	�R��g�2,�ak�q��ؔ�� \g	*ǣHg'?�%�-d� ��o �'�֏'��hH�{\g�w��"=�Ug;K�ZuZ�6od��Q��>�6��9�	�E@sHQR'C\�Zꆊ�y�P�"�3K3m�3���V��>gZ����{�N��F�mvZ���li��8uơ��)N<���zu�Yݒ�g{�` LW��j��z��g8�?tWvmCc� ��)��l�27���i{� L�g�ͧ�:v�@�j�\?w�9BY	���xr����{"��q��M7/~kK�n%�x�9���"�X���j���[���m�T�]�/}a`���>J��b3����c ձo�ƚ�kK��d�ZǚMx��%XG"���KP�'ѱ��ѳ��&mwq��Uc�	�f�4쎀��[5U�%?� �`!�%����{|ڄ��/��?��J�&X�k��G1�Ҷ��r<EA�W��SU�x������,>H���J��hM�q�9��dG/%T��i�t���/�t.�� `Q�p
��}4��C�&���I�SL���P,'K2�b=���z���Ä���,�YAEkLV��5����
���y��o@��%����p�l�u���K��{��ʧ���"H t<���U��:"�(��>x'>i�e5��dh�%A ��O=O
��!�16R.�0�Dz�Tn�8t�&	Љ�N��g��C�Uf�������C0��\GX
� �K��m8�,{�� g@M|�~*����8ok!=������D(1��Z�0��OH����+=��)��	u�;��t��Yj�,D���ըS��5���~)����
�h��z9�)=��)A�54�����d�|W&P���l���\��U�T[ZQ缵�w]V�?
<�QGe6���H�nK*n��c�O�2��O`�Z1T�� B��������ā5Im��ɔx�Ѯ3�.S�����o	�v �o/|�/�E;���y��{:K9��̰E��_N�'y����UX��G���۠/S��� �v�A���<�"���i�5��Qmѧ�Z�9����ݼr�)��U�
u��w�GN�����'���&�ۖq(U.Su�-�5ڢs�DTƋ����(+P�����V�p��5���PkQ�/���X�0!P,�>y��ds��q�֢���2-P��B��l� �UΫ4{J�'.G���߈�'t�"5c�`��47��P���/���Ϊ�*hSda�É�Y.4�0��ϥ��p����>��[/������F�� ��R�h��uq�&M��ro�pcs���U����/��J
F��=��ۥ��ʳ�n탸��'8p�م���@;���B@R'<Y�p�`���sQ}ѕ%8�7��3��ߧ���쨪�`���jq��;Wh��΃��.'^Z���Y�L�;��ŕ[�P����vH�Q�R����@�5�-�M��\�œ����~e����s�J*w{%���|@ta�,YYx��cF՛y��.�r��}�n������&��)�<A�T��a�^b�՗m�$;)�>�e:k�Y�ZfK8�B�ە����?d+�y�4:����X<��I��u[Gl���U�>b]���4��l"I�������x$s{>�"^Eh$�k���-�_���aq"���QQ?C%�)s2���I J
H��%�f6(�Ә������i)�'��0 n��d�k)��e�ݍTo�,G+�����A�a�J�2���sj%Op ����(�g�a1[�NN���s�0�������YBJ�D�T��"X�8`H�s����;��%i�Y#P��9:1cyƕ0�2���k05o.�|=�v��HRɬ�N�ΕE��ș��nH���(Ԭs�Pv~��D>-�����j������Y�������֊���Q���;D���VgU�ꓟ�5�Y�rf��bh{���%�8�����]�*i�K!!���2�nr� "�u2e{�K���Mh}�"u+�<�O��Zzض���������[�R��{�������ם2hf媝PaP�5�f[���	�K��Xͧ�K�)a<7�ע���H�&���:�,��5ߒ���B��gF�Y�H�"9��_�)a�@OM뗢g�*��?O�|U�6uic>� `ZaǠ���-�;�
�}�ԃ��wj ^�}�!�0����nXqzwB�HbT����_Tg�ݩ��L��]�u���ָ �M�_�f�MF��{�]ߋ�*5}��)�oĕ�{��Im�'��c.�O2�鏀(�,�l��S�#B>�Vj���kL�a�EW�1@Ž�՜Ǹͯ�bXσ'�C#&;�����G)K��z���y��^�5l��?[�X*�q�q�dX�X� ؘ�{A;���v)[P��$�`��%��çQ����:�������"� �KF SN�!�"�w+=�J�<[��]�Sx�2�a��lt�f���%� �q�E�7y�C�b~<�_��X�)q��1���Ӻ���f�:�j��8ѳ��ur���W4��iq'��?����%2œS�kG��4F~��,���?��j����A2Y��΃Q3#�L;��	;dW�pq>����W3�t����`��`
��ߟ� �f��n׻�J�.q3�3{*�v�圵��h��`��7TD� ���Z��V�R0?�{ɯqɀͯX:w/�6�	�Xv�P5��f!F���K�0�+d�`���.��Q jn��o�8�.�df<�W+�1��T\�_m��b3単0���Nr!k�=ٜ�%����2#�P!���{u���K	��U�P��5���F�1��ī�,��'�\e���oϦ1�2�Խ�'���ie*{��<�2���9S<��B�b�x�(r���{Y�X�ɶ�'��T@����.�bZ:��!��y�82'��m�B�
�:�|4��<0%~7L��?�����W��Q�X}��	�2�Ƈ6)*��F���Z��\��G�B\[�I�Y��AGY�v������x.WB
iZ��ţ��J�䲷0�X	���1ϗ�y5̀�\��!1��_t�����/������Kq8k��|��q�+ϻ�28ޅN��QM�<y8����c�c66�I(/���~��M&���>5�9t/N1\ɕڼ�vK��g�A��y����'yk������zC�Uհ�]g�ĝh��k�K"HD�n\��O�2*����Ռ�&N�#'���s�RA��^ Z]PG'wYX�p�q	-_�'�/-}6ae����hJޑؽ�4�Q���˘RV�﹠��/�z{�V\`�f����W���˿tO?4Kw������av
K�����-����bo%��d{���jtIyHe�g�a��G쭌Zm%!y�Zܑ`܁��Hp�[r홧Ca�rY8u��X�šg���h��M�m@h}��˸��z��v�r���Ntǆv��70HQ�s�|1/�����Ubմ�ɞ��ʀ���?4����@�V��m�C�5}���IL�Oe�+������ߪ��k��VϘ`��B�U��O����.�4�NF�TP���=�#q�CD�����y�u_މ���h�/Vlp
���X�j�+���_�ݳ�>�>n]�3�r�1W���o6�`�_󷴶�?�l��l q���t_������j�vS��pUB?Dqc�J������q-w�6Y����m��2��kO\��^p|�%�v��X��BH�f-�s�V�V3�:��ߥh~!5�� ��?����h4��;n��6¸��a6�]�WF�f��N�^���A�Sʆy]6�`�S�����D�?�V�;� ��B`�m1�m�X�􀭱lؙ��e�0��Z|H�������qB?� 9�Pe�T�(c�_Z_�p�lJ��Hyx��< �2���n�u\�Eڱ������ �si�Vcy�M&��YV˺��F�N2�M���i�R���.t$L�Wv�+v�dP 
���麊����El���/����^���_:����bE��4��Wxk�W�ՠT��p�P�j��)i�Xx~��',�`�V�?;�"�R�N���0q���F�S<��@��V�c�Ⱥ���z����\�D��ՎZ[�#}���|���V.�&o��� �#�U(������Usk�l>�8U��J*8|F�d7�ɝ�˾�W�8I�|>Yك^�-~H���KN��������j��"��v[)9�7��t��#�;�>)s���V�I�u_���ϡ���rC2晽����D��â~/&d��Y�-�[�Vϔm(��?k�3bq�ˉ���,}Z�����p�ڣq؟�a�s<o�8���#�H]]���VF���8�yRn�����h����-:�'dWz��w�j�	���sc��?�;��h1�C��el���L]Un��X\��a�մ�4��?5,��a NP������D\��lT���\m�:
��ܬ&�s��rt�<�9��<;\�t��y�'`W0Ò���W��6���z W2\���d����e��T�)��2?�C���əV~���<H��lx�ĕO�|��uN|X�����]H�'y�vut�c��6�s�~�y���\ ��v<W�y���c���czǭlf�AO�JdT�IC�VbD �/1Em����∶�Xs桥��=�J��[�'�
n��ځ��mꟛ֘Z�����/����
E~�g��k9H��!�\/u�ͦ%JV�2���͑4F���WIX��T�t�z�yX�@H�!��}S'�Tߒ����k����z�q��xX�o�Q�V&R{��̲jq4��9q�f �0�۳�Ӂ�kbk+	��8�l���OEW��&���<�HV��z	ɠ�<�G^��S�5bygLk�{?~�f��$l_	���w�� ���+	6	�ϯQщ�L������L>3�#�x<�����i=�F'��(�"�d����`.�W$�S�S��>�;G�"f���[��&��HSo��:v��h��=���g�h�l����[�h�0I���2�$����g�CF�]��(Ƹ��އśeG:w,xF��-^��hK$��ב�Cb��g�X�1���B��c&�Y�6�&%�j��s���\���3�N^�t�D����+�M��*�$��Ī�$�Zn��z8����Br�t����KAm�;�{�������&���>/6 7��?��`@1��E��-�v5SjT��vD�zd�teM�����S5��i�D��p���/�i9�O����(��R��C+uI�7�X�8�63�4���o���S���X*���T;v	�͸��Q��u�u�Q�/���p,�Mdr ��TU�ܯ(��	@�ɴR!>�����f>1`���b'���n.����cp�=>:e��h��.Cyx�/k�Q��{�u[ڋ��Ds���Tu�CX��>@��}��u���YA�n)�Ư� �0LfK��]Lmr���}�-�����3�l���$ݕ��3��B?v�QG�V|�c��k�fM?p��]���"[��`����S���p�Φ���E���+�)�"�)x� �;)R�*�w2!���èy.�a�A,9��"պc� :�N���	U�z#$U	��3�u�<J	�C�Cs.���6�[H-�Q����Ϣ*����$���}ջ��*�$���(�� !`L�$���e�Ab��kU���<� �AF�s�|N:q���B?`h�z�w�PJ1�HV���[W�a;\���g���~�$/U��t��T�� ���?�&k4U0{�rV�R@&P�pc:4�s
�=e4�q��T;˫�q��btJ��A�|sn����9�_A�eA]lǊs�.��)�x��x�:�1~�0*��⼭�:�����q��>S���N�l ��Ľ�R��srGۤ�S {z�vV�9��,D1��9ތ��5=��:�y)�S_qzʤ<8�:�(g�8b�MM��"����]2�H�L�Y������(@b��`������g��Hp��N/杄ƕ4�������[0̟b��4�򳡸�wg�E嶶'��#5���+�I�S��-�J	��!E�}����q��j��]f����%��1_9t7�$,I(XO�v���B$F1z���^IrN =�*��YZ��������i��K��jU�z�
��0���3��=*�Y\0��"�8���pW�{�>�>��˶�╱�q�"�{�=�k������Hĳ����9K�? 4e��N�n�����	cz�(�p�*�_�hb�}����73L��KN�7b%�I
��Ȅ��-z
��;6���%p�C�Q��1H4��G��`��b�N��ɮ�T�vs���7��_ T~���
��tc��e���.��(��b��+���Ew&��6�j^f��ӷ��o�Ԏ�.�%C���ͫ�ļ�QQF�8�lw%��h��Q�h=�r#�Z�����~����R�~?�k�|�Q����ѧ�&�,�S�6���#�����I���d'���u�>������i_��l���Ð���"f��ì��j���),�!�'���K�P{%	���;fO����c-pu�Z�ane��2����#���%�jP���I���b�5�F�����i�x[���)��S��s��?w��g���H�h���ݱˎ�Jw|$�c�)�)�걠-{��0ʵ�`j�)�|x�hj#�E=�#.�%(M�'!���,����0'T}�$��$B�oS�`�����bu׽w���r�)V�10^� <��b��q�&�&9�H�=s��h����ƪ��~�7�kI�b���^9Q�������*���rQ`�X����,5�P�M뤪�4>�p�t�q��ίq�T�+ж��jNl��RMG�yAƊ�`? ���@�0�j�ٝbd.���f�9j�w�(�8�Il���FM!���J �:C��s�Q�Q�m��^�#7��˒�JS��	<w0T" ϧ�QMJpZq(j�{�4̱�M���	�xw�	B%�q)[*��Z�Iw�W�=���)�X���y2�D�n� ߄｜��L`�J��"(�;*�q�
�L�G���윅����ˌ��$`�R�V×��^��$�N���4.0>�/�2��e�J�����C+ �&�zGyJ��f�~ϾOQ-\����~0�G3��+㼊~��pՄGL���4q�9mp���Og$��)��6ʓ����Z��4Ѯ�̜Q�QD��W��]T���0�@=#�d�K%_�<T��g��#�5�����<$d��
T�w̻�ӹ��Gf��;�N�ٺ�wv�t>h&"���V�tJ����`lj�'֬#�=\���n<G�"��*名&6�����E!ѩ6V{İ/1�@����v4}�s�e�:Gv�E��J
���d�8*>�#�l��"�(��aB|��ӠAe#���0d1�SIҒGE����w�|w��6��Cl�r*}��jص���\�L�Pwyi,:P����5$>�����\����F8��-�͡C3�)��xxl+���������&�/���Ǆ2��ћҰ��+�v��NR�v0�-��t-cz�8pu�AH��9����	b\�@���ӔN_����WKk<�$(/5��~��8�Ӡ�����D��Fb3�dO�Nۋ$��\�6�U� t��%�����ā��c��b�g��X����j,	2�b2��)�޳�J�9;����xb�rm�V/���;�(�}�o�X=�ׂ��LI�4E�xW�O��k�:-G�ɛq*�&Z�/&�	6�Ql}�� ��Ʊɛ�+~c�^��A�j$#�/�h�ʧ�y:u��{�u3�|�^BybA�ㇽqI�1� lV��%{+��Zd�p���@����PsĜD�����(��t� ��ڀ���	0$��~��As�w��E��U#�ɒ���&n�0�@�!pիWO���s�)��iR�����yN�����?��-I[�=�Bn[f�����X�s�I��*���">��ٸ��it���?"��ͻΔBS[���{Q�k�ՄI�)?��+[��4F�c�̇���?+Md��9G��إ�#��4a�u?i,�F�3V_���H�Ú�ޱ+A����)��C�)����;ؗ�WF��n�}5�L�����ߔ��);
L]3<���f��/L�2�r靳h��(�J�'k��6C�=,Df+��0Y��Q?�x��@�as^�|-����*k]i<����ݲꫫ���?`O�����L�a���h[,��%�Zu k�,���w�ogy�?N��a�����6��LP工L�Wjd4�5���%V���|�/�el���7�S�:I���
uN�{�|���U���G6���Vw�"�W|t�=��p�]~�O�c�������)h��t.!��^{�����}yd�d�a�q�ѩB̓�z2� (u��[��1E��xv��-1ҁ��nk��/><�
�"���l�^�$Ϭ�@����V��,��bm�MO[D;��`���C��5����gs$V�ƵՃ����j�r�Ȃ2�r_}�dR�H�������PD׎a�	5k2}֩�,�^�ɜ�E��7d���b0y��қ��z��Ee'�"�B�@\�RO&�y���!�d�<�g�.�qƥ��0Ʃ��!��^�i��q(f���MND�������@C�Qn&O��E�Ĥ�>�/g=�`3O��Y9��'@gT�&g|*�Z�����}؍]~�O�t(�<�l�l}V�z�m��׊y5ɩ�%�E��R*�q��E+P�e!6���Yֶ�xØ�Qm���ZK�(����=�*��897��
N�{P~[Y�%��Ar޶��?\s�ж����p��{&��1V��:�����*͋���%�#���;���_�Z.):	�R�+wBu0>��� �l����/��&�a�K5X����{��r����jt�?�!�,]P��FDLeTB��5+В�b��+U�k(��C�le�s g��+�+RV��������̢"R<借�~�N�g�D>V)���]��|��;��Қ�o��{Qe���F����Tr�e����Xx�)�����$�;G#F��D�qA�ј�ct��H���y!�� �&�3�H����j�v�`�`E��cјWG��N4�_f���s�=�愂}md��]*ѿ�M��H{_r�\]b��w����^FxIMV��Z�����ȖL/;��,f���sNMx�r*�~�BNX�Fs˕�-㇚�F>ן��=3���Ƈ�֠xRK�rDk����,���|�5�ͱ���N��`+�\t�e���6S��7���a�y٧�U���.%�I�z�@��a��&{ '�B�bN[t�*�׍����]Hǟ�l
8���e��a�tx�Qh��P���.H��2L�]J��Iw;��n���!�i�{f��ҹ�K�R�����露�;��7A3Ɖ��.E�ـrQ�QA�Xû3�IWv�c�n����ĳ�F�LsܿGIT4���y����>�hOSO2�w�h�Fg���#��o�#1:h�#dLq?����������1��Xiʴ�;�)���-�W�@ȸ=C�_i�>e������u����"28u0۵��i,bE�����|����?/><�XY��ŕZ�I��d�)o��߇bN	��ě¾I��#��Y�v峎yCTt �R�}���6��ã�&�`#��DIYJi�xp����3�Ѓ��`VZܛ�l%8b�` bd��ЏCӼ0v�����96��n`��~պ�F��Զl�4fΏ�Bᔪ Z����v7O�O�3]Ͱ�wc���r��qMh��f�[�����MF�ݓ�LR�Yk�����C��#b\��'�n ��"$�f�˫��K��swgvQ��xV<+�Φ����ՐR��03D�����^�.����
/k̺!�X3��߳�� ��3h�6w:éT�����j� ����k@eO���?�-dBp�.�y��"_����b�A���	��B�H@�Q�FC(�����&l�G����e�i����3��5�Ns�܊��b��|Q�!K�(�,��1��\t���:%�a��~�[��`;n��۵�գ�(��#u8C����&���'��l�-[��5}���9n����5����B��D�H�ɱ\R�J#�} �E���V�c�����F��������b\��f3y�lǾ�8l�v̷;�}�UMe-��N���x)���e:O��o Ϟ�y/yY
�h#��D�zy�r(;M�����'I<�ȥ���b1kX�)�/�uR!��7�h�W?4t�̵��(f'd��&��w")}
"ى��-To���DN�u��R�/�;�P���qb5yA��p�F��
�y��ô��i����&M��'������f��l��w] Eu��b��9�CL�Ž�iCY��L]n5�t_�;=V�����o��=
K�]��ƪ"�#��Jq�ǎ�髾�{��}��1(�\�8�L�&�x �6�]�
���?Ug�&y(�<��UYY- ��cC-E �E� <5��2{�$��Ύ�f�v��4���J�����%�aO#2`����ID,��ϼ����ma��P�Nn��"]tsS�ЛW1�wy>��j��5�@��y��P�U��)�5����^�3�6�7R��؆��Ĉ �R*�+q���D$F�i�%/qzK?�43/�P� �j���c�����:*Z5V�x��8�C��JpF����g�N����@��HQ�ٞ�O����ث��;jw�請��)�P\Z&D�����k ���u���Z'�/'UVDb7PWB2�!8`�$^,rb��=?�4�OT���{�����be)._�C��$�k��!兌�T~�.���Y �>�th�s�"]������Z��'�.A�Mc%{n��S.��Zg�����y�ٻ��0O[**C:>GeU�a�>�=7��#f�Q9P�F��E���&�B�À{�@{�4��}d��5��F��K��+�.
��%ӞI�W4�����<0�B�n��m���l�9'�~]���Z!�;9��)��K��I������!�
ՂXNW
���������j�rB��Nt��
ԡ�1rH.����ʎD)W�����7����hk!���8���R�R֩�0I���~*� 蚗���ܿq�2�κB����������}�'lk�����Ldޔ��{�4���?��
o��%�Z�sdhP�rҾ���K� ���Ԩ8���l�10��q^��h9s����OZV�
�>4F����&�L�?�x�W<���C8m��1�#�gx���u��f�a�9��� �û-��X�aT4��x��ZPg��h�~=A���h�hh'�/���p�c��I�t39!BQ��vb e=���̪l�V=��F�]!y\f����ab��p��Ӫ^�{�O�\m����%�'֠~P�)��ɽ}�Ҽ2	�Ůb�'S-D�E����j����P%c]��jQA5j��,���e��m
��&�0�|+ޣ��1
� 
m^���$R*Q:�\,(yӺ,*�3t�w��v�}�����mG|ȝ�X�!E�F��L�HWFJ��L��xJ/Xwe�th5ұ-G�➜|��|U�{�ܥ����#�8�j /�3��=�f⁖�v��T�/������M��^�l�A��Mp��вSgN�~Y���J�R6[�`�g9�W*
�vC]	��9a�Fw�Pi��Ð��Å���) ������3gi�̢���t��90���[�$M���Z�����גy��B7�&Ij��Mنݼ�od��(x��1ZL}|�Q5�Ķ�E���%��-K&�ٲ�o%u�Mx8���o��� ���TC59�ֆ��w�/y���*�5Iጙ��_�B�T��Kq'�䮯��x�ծ�r�C;��V�L��i�zG�q מ(&f�w��$5��_��f��N�!�UzpH��?��gڐ�,���2�"����eY��q����>TCͦD$�����������\΋c��Xt�h��e�@��&@y��V1a#)��Jk��;!"�l���4��D�mN�R��p��C�j���w� ��Hs��U�LJS��A@�2M��^���E�goFć4�����U��o\��D���48u�qʆ��Fa�u��x��/�`Kn {FS_������^��M��(����^c��F���T�c�@M�o� ;`�.0+�;�"ࠋ�%����0}ML-�����S���}���n�3���nn�<R�|�C�U	��փ�!��lV�Z�~2g�azH����>�2��=�EJՏ����+�U���yg�b�]�^�����̂Mj������ox@��!a�G ӎыa톏Y���t��������Xu���=�C�!ߚε" D}'�b���)�J�L�c��ɆM����O1Ea�[լ5a�~�� 
J3=R�D��6R*Lj��*��p�#ӇU=�����0W�bhS�R�Az�����m�?z���k#�����/����O�=��3
�����Q{n��łg�Y�J6��H�QT`�!cY�Qe8/�r�e��T��Pc�mH�@��Qs�#�ɬa/W�o~1�4����BTb�y�0����3YQHW�y�G����/;�zۂЄEIg6��}]�}}#�k�}־�� Dq��B���8n��1Z�
�����6�4�A}]�f�q����R}sp?���YT+�,���(����!.U����@�u��Գ��k�Kg�n3�1����3{e��pj{�"7�a�rSX�����[�a��U�Z^�*�s����4U�$�w[��J�X��������}E7�$�4ǿ�ſ��B(�z�˻�]6�ITm7g�� z���Z������$gv�T��x�1�[%�x,��^�6�bދ��Ns�R'{Z����*��
�Ϲ��ŀ+c�Ӓ��Ycm9���p&=���wЄƝA��e{v��t�������ܨ'�k��������$�e��ۻ����j����$�&�i�7���#E=`l�P�X���� U��Ԫ$@y�+b�9�z8��u�Q^9#��d��*[#[3؆���C�E3�sJ8���S�xk�7��|W�Y���թ��9x-����1��!"�Q��"��$R��ʸ�y���'�"Y�w�-ruY��ޡ�UA���zD]� ��\$d�'v}���
����%.Ѳ��s?Q��_���qX�j�Ĉ&>��������X�0�[4c�W�K��O�(W�/��Q�uA�	Ͱ�ױ� ��4 ��䭛�ǣ� |��l!�D�d�xA*M�^�&�0����k��@uM��=(₩��cn�+��=L�$7%������-�!�������G�y�Ujn�yk�5b��PZ���G'�3�"]O��Ӫje���~�y1���Ԝ�{��D��u�04�S�ͥo�w�v�� z�%:+۔WǪ�/�t 2���0c�1ـ�tA�~-��M,���o�8�8�\�@5�S�~�=kԉv\�Ϳ����ِ�aog���-Y%nL����Tᬣq�����a"��v1�R號�`C�?�#ߙ�0��������T��,qܸ�͔ɲ>O�^�
��&Nu�f��e���
�>��x���T�.�si�����E9L�J�X���j�g�ߪ����Y]oD�[w䕵i9��*�@��o0ӧ���,:ιf��P����e3M�V�f��"����r�������k�u��h�^E��g��w��=�(-���"�i����e�m_�X���RE�����B(:�i�cp���sq *�D��1:j�������k|T{�Og@��?5qlK�q�<V���_%�_�t,l����p1zi�K}sG���,�n��x��K��FG=���s!�L�Ђ�'_dN��M�n�W�����|JS��"v��Hi��7���+���Pl'��*?�9׈,�s+���!�����5e[=�<;����h����O�ހ���냉�>��*��yi`�g�}ec�n=y7k���T�V�$x��fS����J���dl	�e����B[�^�ߨ��,�T��1�7a��D&t`�-?ژ�c�UK�y#�]f~�Cq��]`!��
�DʒDs`ڿs���M�R�������M�<$]D��ô��=����?���j��]TH��������1��/cP���ND��l��+g$��ѐ��PRya�bL+cSH���K;��%g�sIl�l ��
V`՜�
}_��t�(d0�uD���^�2"Ź.C҄V5��ڸj�b�dv�t^yo� ��3�g}/�0��}�[�p���5
=�l��½9	��u�+�~�Y%�u�ĸY{���Yʩ��w�8��m�>U���	�W�z^���\$��7�&;�lֲ�.R�/y�Y�CK�񖛕xc�ږ�ѾXB;�e��^����}?c��}�H�2 �i��y�9�c��*�|�o�0y�צ6�ܢ?�[���VZ6W�x5��5�`�ZHM���f���˻��a��@��R��k|�0����:Mn�,�R9I+?�_��?�m� �@y���vd�tC_�gKF&Uϐ6+�w�v��C�bL0ΰ�7?�E����A�3D�17] 3���6�� �\(ޅvU� ��ފ�e3޹R�
��A��� �;m覍��E兀�A��mrss�Ȃ/O�:^<���;ͪvq�s�	�l��뇚��|��IZܹZ��A�D	5�b؁���
Ɏ/D7�8{?[g����m����S*[���՞����N��&�[������jL[r�{r�tҀY#|T�Uh�Pojz�*�M�0���Cx"٩ohn�4��Y�d��y���/����]0&���_2���,�~D��|�$"������~��H��If0�!��E��sv}.�}�!A���R�D�ne-ph�/�Ռ�����S���L]��\1��ʋ�1�d`"�>G��]��k(���\?u��%����x�م�yM�U8	�>)U�$�aü��Huk�x'D���\�2�j�K(��S�<?J�o�~�Amw`��4E�I�Fov"�ڜ���3tX���:�?E��BM�|xp@ C�$�m�����ˌ��l���i�)��Y�{�d�n@x�r$��SE3�sͳ�ֽ�h��:��r���v���p���S�v��i)�Ҙ=#�S���2|��L����x���lS��&l�H(������
c������6���0[Q*)�C#p�����S�Y���c������=�d�V"�:�&z�V���)
*��h��Vſd�й)ߧ��U�o�h	�Ǆ���1&� ���cA�۫0��� ���{\���Q�:c���؍�eQRǝ����"�������������4G�!(�j�$�_��{�{�e��w����p4��L]v�"�)�62��9`�X�@�MN_��}��������Ͳ8|���{�S��o$k�B:��e��ӎ����('�\���n%�8���F\9K�?�k*>�[���+r��kvu�K���~k`|��t��!��c �Z=�������sqȌ�����9�x ���P'�R�*��b}P��Qp%�m��&r���dc�X�ڳ1L8�y�W�Ư�4���ٝ��ى]l\�u4K�b��y%q�Cs"���B�EbU��W��4!��`?��e��-��{^���ɼ3
f߭Z?>����WYO&M�Q�]�{�V�J��A��Z"e1<�����9�X�l������H��@b���b�'����ĵ�E�!�����x���v�3��� ����d㡑^_}�׆�7��q^��I��FͰAl�e�n�7���S�_�`bo�vY��W�G{2 "�)�V%�V�S��s,
U�#�3��Ҙ�Ͼ�����"yꮊ�y�o�~d,琊M�x� 8Բ������*c��A��-��aL�,�LB7��_��`e�ٕWK����%�d91c��u�g4j*�?P_�ou$�m��V{j���&?�u��B2|��N�|�^��[��r��U�O}�������X!zQ��9z�����6�����ZϏ�QTբ�X���]�y@-/o2�M��I�o���]�
"-ZzG+G���7���+�<�Kb涶$ |]�\IX�/�s.$���рa��ivE_�qD�R�|��?�u p��\�=j3=�}�V�ي����
�yv*O����>G9;6�?��X
mn��tY�+X;����P��f?MS��zԧ�Y<n�B����D}A܈�	�E4<�r1�6ftՐ+���.��BLm�[מ��7�@�N+n����S�C^`y�D�1ߺin�J�-�K	;�/�9~�UYY�\U�a�/��K8����~Oٹ���C\��PD��[�$n�=q����w�j�*�:]��$�����K����{ǀ�������"�e���� V�p�"<?�V�!1��P����zj�����0�pS��W~� X��>�])��x&���Ƨ��!}r��F�!�z����¿�7k$�S�z(����*�p��
�|�*�@S���CsCݐ�f��ާ�u�ɨsl��pb�e��b[����qD��6>ĨW1J�MbԚ�x�	l��Rx�ݬ��0[M�zl�ܫ@=�=Z�Qrβq�)���'�Nf
H^�L�W��%��v�qm�&�M��τ��$p���A]Ydu��;�p�ӽ����8�[Y�h�Y����KFzĞ>� 5��I�TE��;�c��]����_rU��'�GH-16��"��f�@L�D�I���.ܶ2�t��5vu�;�i�g���/���/�z�HT�<�G�Or$a��q�{kI�bb� �*��
��zw
Q@�\��z)/ ���]�;Kʣ�XЏ`�1��r^&J�t��q���X�LWb������@4k�����ɧ�-���x�;����+p�41���� -�!]�5J���Z�˩0��`k;��i)�+�]�����F��X6EYQ�K'�c1E�S�q��Z.5�H!��ʁ�aA{lfwP��׍>r ���g���y�ƅ�m��¤����c�^�y��V�VOSzY��3��6V�M��L=5���N�ڜ��8�����
�%��*�DJfﻒ}�_zU��Y�ȭ��+��7݊��H�6K$�����NZ�8�*9ǅI�S0%��ϗ��Q��{������:%�Z�B�*�ٜ?JT��I��ȍ3�s�� �ds9��Rg�1��?�?��{8�����8R��œssp������ZܘB��y���k������V���,�,Ҥ�;Yl��E�EZ=-iJmH����P�<T��䄊�[za�1U�S����q￹zT�;���n-���p� ~��&�������s��_> V�va됦�==$�9WVh��^^��� B����$W�q�b�V-��w9�p�L�z�Fxz���i�mZ�K��3]���o~!��'��ѶHR����^]'r���iZ0U\Ǚ�4%�4���T�a9�?��lޝ��jeA�9�#. �Mc<>�1���F��n�>L�������<:�����FR3�!n�";#���P�T$Z�ľ���ƚ飯�7�&�nj�iXe:j��A]�[�1��$�ܕy�$\gK���}��	��?'�Ms{���W�{gﻣP�'D��Hk+�MH�7��R��Pk���)N�cI��F�|�Q��!Y��,���w��?0tw��v�,���
��r�$x#��~ �#~k�irr>��$?�������@X�o�꟔�f( �;bi%�6U]3N������|ѕ;��B�%�A��Ф�-ƽ��T��$��B.:��4q�P�7��|5N�Ɗ�Cz��i�"ޮ���̧^'���(�O^g��a_sC��%��q����$�wyx���祝4l��&i-�(�� 5v�H��^��������\'�
B���ĵr<�%p�}˻F�*?#��$ϣ}�T/X� |�5z��p�X�@���!�P�T�K@Fށ��}��:q!�-�њN��b
;J�zu-yUV�#�yY�0d�[?TXtѐ��m�@+n�����͌������z&��ˈrހ��A>kѡ��2ܲ�SDb8�����_VM�Y2��-�)�пʊϖ�gL22����cO��Y�J��B=�C{�dx<++�q���P>����V�'��՗l���RB�1�ҕ���	��_�o�D���ɡ^'��h���Z|����	���3��;bǠ���@e�ـѫ�/�i��ʡ�A;�,������Z�غ��Cjk	@W�IH�����+N�=���]�W�o��ݶo�7�""�Ao�1:���ZUKI���EN����Ľh}\��ص����w�y���m���&��Ř@Õ	�+_G�x������g�~a7���v@(a�l�*�!�[P0/�}P%E��|�Dk򽿕`��K���%w\���Em�}��C� "ʘ.����pB��8���Y�a��h�D�*�-(	>3-)�&́��^A|�* )x����-lLP���RZ��� ��A��n��fM�j=����Y�j�����(�B��P�~��@���(L��B|�C�zΊ(?��9�#ҷ�p`c�nN}��g������ �|�U
�1��)ItiY�$N��-���	T���7����\%�1��١y����r�� ��Eָ}�r7�;�{2��\^��x�g�j�uՍ�/��TB����A<S��v�t s�;zjiq؜"�wJ���A�����Yu8�̚ځR1�~�L���ݤ��.d,�4L��^��E�z���Ī
P����־�w�i?�H�o�a����.��v��w3�����a� E��/|�#�&�@e%喒�@�P��C䥬���&���f;8 ��p6S���0�OU9.�CX��23^��ps�����0Pz�:z �_�ʃ�^��� Kg	+>#&��ύ ����]�Т�T~�����`��z��&/�wQ�e8�rV4\��;�\�z<���JyL;���T1��<��my@ְ_m��X܅+$T����*z�a����]���AP)V��b$|�r�}Zs�֣P���ɦ`��]O�E&�iͦ:�_����`8�sU�:vD ���_"E͒x����XӾ�= 䎸�o�H+X��+��]�3�����]a<�1�gFo:ש�BA3�]=���yB}@��;�ﵒ+}�Ct���c��ju��Ж�'1�P͸{!��F9�&��Cl�޻����i�d��� �wˇ�ƨ2�CU|�%�W���P�؏ڕ�V���5�gژ�d Y�)(����d�,y�_��y���-�ˎN^&�eJ�e3��<6^Opв�ƚ�6�pp���Ý�H	>�d#�xar���o�Y؁��i��Qܗ�~Ͻ`8n���_4�W�ϣW�³0��O:	q�|O�a�A�8ׄ�����o��G�/;�ٗ����:����T�P��/��-���8�v�D�C%��t0Q� ���T�|@K�s$�(�߿�}�Y!���P�5qP{��S�Ya�u�7o��_�Qѕ�̂�4���K�;��&ɺ��H���۹mA�]����'ǥ�! A7���  <4`d�͕�Ҽ�m�N��q0R�ō�(�S�_/��R+)�(��o'F����$�N6�g�*���aD����Ȑ@#~|���{��^�i�5�/ϗ���a�>�v�i�ynQ��Ϣ%9��BS��xl9w\7cf�r�l��;P�U�m`#�۪�P�6&_����&8��յ�a������|]r�kG�8w�:i�ġ^�-�����\��]sp��i?9X�wkb?͹�^҆w��d�J�[�W}�yz��)����ã����w�. ���a	 �Sr
YCQ�L$MC��;�Ș ��T���2�M%REe����"*����~"W+��
ˊ�<*Ҡf�u�7���F�Ec"#����惼2ѵ3�ӽ�*&%�}��O�q3rǩ���dm#�.�a[�h���f�,���  ڳ�6�a���G'X�9����I&Soyk�v��¢��i�j�;Y�g{@Td�W��"�`F��Ta=e�yc,=�Q����i��N��<J<�L@��>��<���͝��ߦ���˚�i��1����Jq�iQ�h�b�3�k�ܖU������� �d���\�A]3��Oe� �Y�t��=Y��4+���l-.����?y�8T-��v_�N�[�=�enؠ�4���qq-�?J�dJ-1 NV�7�ك*Y������3}��{M��zX6f�eN���hqk$�NQ�� ϣf �T�~�Ĺ8<�}�&i��CX9�Nė<�@[� �����2��<ku�{�u�N�9A�p�|$l�^8e���e�\U-���H+w	H�>6^Si�\w�	n�}}��w'Y���E���<5L�c�AZ��B� �J�,�t���WO2]$�xIC�,��e@�~���m��	w�M,������J�C{ܕ�g�)Sg�w�
e= ��޶��7ه9����d�h�Pj9�Dƕ��X�Q�ӷ@��`��>���_�AO����3��w7g�4^�������&�M�h�/���0�F���n"yv�K��(~�:���A�o��2Yi���ұ��m;����W	mDH�f�/�{gh�+�c�0�_�wM�	��©.!a#��tg5ݙ�=��bEQ.�/���>�
�%0%�J��t��jx�ǸS�����������sT$P�D�5V�s����l!�!�hTX��mh��:�2}�^9�N�­���;oK�jF�^��;�+��R:	?�	���~PX�S�lW��("�Vކ,�Ϛ�靉�E�r8�
����+s}ؘ@[$8�ѵ�O��|�LJ%��A|�1��d��7�L����l%�9;�M�%�Ab���m�l,���	Rb2�6�����V�O�]׏8���@i�LM�X���#{��FڠC������;�I���1� ������R��ʟ�9i���b�5
��yh����N��95i��`I��2C�}��
���&�#&���gs]m�҈�Pzgn٢[�zd\D-6��v�p�4:G�\�� �<��Ʀz���Q�G�>��K�镘b��l+�K �}��>î8<Uو�t�b����2���6�>��owL����	Id{����UȏQ!d���If��ty�Ef�GX�@K�7�o������:�,.�����s�a~́���e��uZ(\�մ�7{$���H���Mޡ}$G�4�� T$����ԄC�1�%��1�)a;��*��C�q����6&>;5wΉ����)3�Ki���vc�U& W,T�J��Y���YAVQ��f�`ޞH$���~����b��`�b0H�IP����(X�	iΨ,�G�$�TI�`��*�o�c��Q����u0R����;w���Sq[����;�3�W�����i,�?}Pb)�`�eҎ�]B~H��85K�_-�:=m�LFt��?�����u^;�{��ǍK���j�'�$F�p�:�m �4CZ.�)����ď�]�N�z��?�L�}��7��LJ�+
��qlDR2������%��U�6�9�R�2F��PI��J8�i~O�ژB�G�(�_t�M���/o�^�������G��X�����_�o��+!�����8�H�:����j �GH*$e�v�7�Q~�0T��N�$���zJHn2��!��@[�;�u��DP^ȶ�K���bE�>&{���0;%�w���;0�ӥ�Z�H�t8�l��X��\'���x�4�,��6�����g⡏�G*���J�d����I�#��+m 2��#��±dZl~��ә�W����)m4�q�#�����o-�L��F˚��Ӓ����w�u�[₞��=JQe_xd���ݞ�X�ݵ� ��q�ه��yF>�Z�!��M��d��M��fE��r�k[ ��(1M�J�	(u�)C�"H.9�P�UP_WS0��O�{l�wA��G�����$����Q�����#%,�g��B�aGvp�*_�{4\~ 5'x�ǝ���I/�'l����ڦ�̷��+�i\��>�ba7[&
"R�O���)��Q�'��DÈ��#� ��e.o�橭"2ZܩM��mVZK�Nj~ ���:�l�g	���z��=eâ���z���-m��|m��Wp�6�K�����w��X���-�����Vo��[��v�O2SdQm�� ���&�^�6	LR\�����%Ç���3�E�Р]�Ш@���j"�X��8��
�s����ɺ����c|.2K	�n�җ�. ���{���ژ�#���d1�c��������6C6Tq�E9r��T��	}DW�W\�Ԭ�����V��d,Ta�]�FGU�X^�5n�S|�p��,MŤ^;�� �ؖ�os�5(~�/݉`G��N�׭�"�b�
��?]�ۘ)�G�����x^F�2��1Kd}-7��X;�c3�{�알=�(�r@*��u,�}Ŋ�*��QƘ�[sʕ�6���Kŭ%��V��n�ՙJ5���h0�`�O�O���Mu��p6� �L�� `���}�-z-ٺi^����֞d t����Ҏ]�>Z�$���a6�jW)��~׵�(Hػp�V�±���)��%�~�Ѫ`�:N����8f�u"3�m��A�x!�K�3v� �֤��8�i�*�����#���%��W+�T}"�'Gt���
Z& W_a�/qj�~�J����a�]_����y�xY�y�ktd̜T�C���&�=�����(��#  I��7��KӶ�3d�3�r�Om������}��t����.�_�HI���`V�}|�B`J��D��cN�W���aϊ&�O��5�$�2�P_6�/��j�ņ&��ۨ��my�O���m�bީT�m����#n����D{
���2G)�5����] ��.=�2��J�jE6s� 	۬�\�RXE�p��S�Zr��aVWe���̗a�K�'˙�Ń�,�3��n�x��b�p,*"���
���~j-g��ޮ�e��]"��L���c�j��JU$���c��gH}~vg�بQ���k����d���z�r�n\p�+��p.M�+һ �(=��߾ʚ��ϵh��i�RV+c��T�ܬo�:}�uH�Q�����)P��q��������f{��E��teB7T�k/���YbU0(���Á�� ""?@
��>�=�S�1�����gi6Km�%6�sJ�ZB�ͼ�i�
4���xN�igGx�M,�:%aJ֩yV�X�/Rx���H�p����~�x��#s���G�M	 �n��s0j7�w§�ݲ��|��/�1^[H��|�H���C�ƨ���� ����4A@$G��U�P�'6cXV��u�Vkz�;��[wb��C�K��QǧӓMo�
������J�W�܆��y�����Lˁ
�#�e����A��K��IA
�]�x	�\T �Wx�)�T���C�7y�s/�1C��+�RȄ���w��xB����~R����������m�Y�+�M�$~ƚ؛�y�����+&�c�Ӿl�������J_���Y΃\�`�7�i]v4� �v��t;�ϺYke�{g������-�p�����j��<S�)7�T��[�������|~1ڧD ��nG�A+$z�-* al��������+s�*�w^ܖn3�#���TX�����wؠ���]��%xRR�)#f1�|~l��5��w��57���aś����
�M�z�B���c��\�"���h�d�c�y�h�"W̈ٲ��5п��qR6��wі���Q�V�9�8"��\�lp��B��rǂ^\N�>�����ȹ1[%Agά��B�������Vj_�p�3ة����d�Uw�q��	[����Y!�v��7>�Ƿ�M��1�Q�ƚ�J��$��T��]�Ի����J�F������D!ZU)Uª��K=�K&��f�^Ir�E�ԡc]+S6W;y&Y�a��*�DE ���ӡ�QڥJ�N&?8�� ����D����=���+��������aoE}{l��	�UQJ�o��<H�5�q��\�tQ��*H���9K&^k�9�{��ܶ���*�d7�>g�z�W8����+U�ŷk�����?u4_��W�Q���P�L��[2��5���W഻��m]�L�\��!����"�K��H-v���-AG�c��4!�4u�В���l�ýg~NS����T��æL{W���.� ��(��3 ���W�l�M�҃�f�%����Z��ᳬ��*��#��e�����؃��Pmj��Z2c��B��Z�0�����U#��	N~(��E<N�l=��c�M����L�s���\���^W5U��ޫsn���o������vˊ�@�e+��g���qG�hv�h���X�~W��W��=���X��l;�_U𽔪��&<I�� ڱ���vqC �t�����lbT�g�x��!u��'E��(>5���"��J�2�2���RyF�=Jn=Z�lB���-=��ƆP> ����/H��jW?&į�&������u�� ��Vz�"�J�?
l��#_PdX�U��k{�W��n�sxuBÆ�}#�=Q^������%���Dqf���. ��ײ�9z���rrpE�a�x�����S�4(�k�I�6��Lk�JZY������?K���oa�}_�`*���}W�t�meG�̅��jLڻ�9	WL��d�֍G?�I:��I�ËR�6�F�C�v�%U�yCg���E�{�D�j��R�2�{�XN�V��nK���>�f�%9q��LR>m��T[�yO4�G$p��UJ�TYUN&Ce�U�*�@�;�q`�`�h����Am��o��	��b�:\�Y��Urg�9�T}���E�dk1fHrZO�2�Wg2�9����� ��[�Y�>�5�w���G���*d�7��� �a{����2?U�Ȧ�Bt��I�]�޶���7J8���E�,�p��B�A2=�ͦ�},��+C�H�UT������3f���!�D�]���L�x�rc6�`�H��R��!�V*ɏ~�r�G�b���i��S���Urq��H��刂�����9��V��.-�E��!�p<�}[|��jW���R�� �&�T^)�v�����"�0,�#�,��������v+x<��ơ��KP���7�TP��lHE�5��|��ߴl��_:����`H^B�����=j5`�,�Z&���Aj�skd�)�̀G�f���/|Yc� ����!��
{_��`]�AB���q�YI��P�1|�O�;�v��l_e�tK��=�&��7=�E�3ʖ���^9im(���x��[Q�)PQfIk� u-c�_* y�Ǻ]��b���09	��qO�M�k�}s
����<��!0h)��	�*!��c��=͡J��ԋe���z1�d]��j��m��]� ��03��4@3G��>?D��b�0%{�!�D�+ԟ�5��^_#�Lh��&6�����qh���?~-r5Ǯ�z�hj���(�-�t�A����G ��R_�����w��ּ��Yg�S�t�يb_���d2�aj�ײ%0"8̱/������r�:�(�p�|4it��LC���iRt�	�C�/���C�S�c��9�S�S�08�k�A��HLKrt�����P��y+�Xo}��������K)YA��Yuem�}`>��(��G�D&��Lyj��;S�1c�}!I7�x�&���t��o�z�� jI�5M��y��epF���թ7���8f���<�i�CJ�iz3��o�y�Z�D��B�y�#�}O1x�υ�.���n瞟�eLo�� �H`��rW��e{�g6��y��}
��-	�/=��滢�3ۮ^Sٮ��'�^#�I�c�~2���	C�z�lН�!���L���m�¡c�ԣ��l􃳋'��qP�p8Z�l�@��A��}�G���~��X�����n7}H��Pb��ȟ������7�C�Ĉ�/ި��?����CpMM~���j��V��@gƱ���+�CF@;��p��Ũ���^:�Ǔo\�V��xz���;�P��0:&��V���6�G7����<`<g�̌|�It3y~h�uo�u�@�
���֓m�QE�{3)l=��kƜ�{
��Z�L> [QRK�Z�{QL�6P�`#��������D�W]���=(� �Jln)!����F8hu4�@����K��EG�����T��=��K��M�B~�}�r�`�^��i�(t��Z�@Ӻ�]:�{���0s	.ndSEn`rBpC�gH�8MΟ�H�A�igX'vb�`��lђ������z����s�f��4V�f�p�.�'��l�,�Ea\2W���E�e 0JFBw�0��v�f9A�k@�-��,H_���2�:�#�p��Oc���V��u�k��y���6K[K0xgC�><"?���Jq�������J�4��2��n�uVEL�Z�%�� 1����{]���f�CJ�G-�
i�]���������3$�e�gC�|-��t�-�(���f��?���\��2]!~�̷���E-Y�۹U|W�4��Ro"
r^?��9�O�� ������"���(��3��ٸKn����:6ŷA_'8&-�)L��g0��|����?`ȗUD��'��7�f�F�+qWs4%9�&6�����h��(M��s���r�nÙn�c��$9������'8 �)ِ/��)R*�|��J�N�G�($.��2&��Ԩ`e jY�n]BB:	h�F���F��,C�IE���:�����Y$��@a݆�j���o�)"׼����������_"���-�ʜ��A0�8퓆��RM9��
q1n'�NK��w��95��8>�r)[���v����<��*��>%/�S���ş�P����{���mp��L��o�m�<h����U�����l6mk`�]<�c�`�Ky�A�A��O �/\Qa�0�XX�'�*R�e��A�Yյ���l�Yx����0b򙭸B�Ka��췸�H���wȯs�>�H�M��l�ߓ�B�%�,����3bo��@'^S�P�j�S�mO�l�9ך����>��b�#,����U��2�/m��E�s_����Gh���d�����O�sC���_PJ��hWFO�Q���<����y~����{�kqߨ�m�Y\d�������&H���摎�>h		��8���`�����n	i�zT��c:ݝ�l=0�.��A��L@MOX� ���+��@Rvգ�(��;�8���54�QJ�Z���M5U�b��� !���	�in�q���ᴻaC��U�7��SI����]�m[���_"�C�Pm��Q�
����&C�����s?w3g(��k��6E����|s�ҏO5a�Z��/���:��V}4۩�������[��.n뭙��r��1�ss�.�.�u+L]C����}:T\�"#u��k5�ρ�˳<�I�߸)_~Vh��[��C�Y9k	�W�An�B�/:Õ�xW��o�Φ�uW�C6��T;�v;�Tj1�}l�=���Wo�!��%@���M�l���4��s3��]�2Aב���A�ݍ#��������72�B�"q��U$\ǰ��t~9eV�b�-@�o?+nC��񳃣$��"JMM���q� s-�n���W�*���r{U,�H���8���^���§mq����7�. ��`��_xKZpA~�cͭ�+ ��eM�P\
���a]���t�<��C?/��+sD�+�;�议���NK�	���Lz��
�_?:���V�u`��ߤ�W�m����/��b�9��5�k�q/,#�61�����p���Y!����Fk���E�ŉzCI�܇�t!��(�!��A��r�+�C󆒈hR�$�2�����Dg�lis�)s�c�R�r�zA��=�$���TQ2���u_�������ʶ��x,j���g"Ej��h�����Yp'�VǶ�� ��ۇDQ��ɜ�gm �_Ȓ�D$�V��E�5_�Qc>�����쵀vE�\�z��R_��z�b���
[�M?���p��0퓖�n��R�߀��1��/�����e�4�c7Mв*��C��ʹ����ڵ�@������ۓf.�$�Q.xC��Kݓ�a
%��߁x�$
핧�/��R�`��d��B�X�_��UW��k.-!�L����ʰ��5�,Ո��[��i��hL<U�W�B�{v5:�"n�ʯh�b��=_�����u,���~��t��g,��-KD�;��*=�,FT@XpCX <�	�
�@�|}��鼙�XP�F6��8�VЪ؅�L?4��K�r�|�����ۃ-�L���0 ͖��HM8��6��d��F�+�׽x���weza��opb��j�y"�R��~��f�c$��E�����@q`?�Fg3��iF��l�������5~c��::�,��`��bU�*pU)me�u�#�pp	⫯+<����Wa���S�-u{�	�F-hP�V��q��NM..����Iw�HP-�
�:��x?E	��j/�lq�+'j}@=�-N?��Q=�F:F� I�rs��>�Ĥ.�m���'��n$\�p�WS:�EQ�m���)�޾_�_q-��5�˷�������ǰ(�e��Y���~&���k�̲�Y|�AأɃM9r�����+=\�������=���^�qF^����dF0>Y�ݮN�zT.�{��Ȟ�����d��A&���g���9�R����Dw�O1�~�{X)��'I;�v�&�*ғ7���:�4�n�X�:�E��=�oqZᥲ�e��lˎ)���R.�Ҵ��yS��ĤwxJ���X+��L#/�vp���Y�|�=���3�{������nl�8�$讣�׏Ɠ�ʿ�^� ��q��������n ��/�q���.�7�~���~yꙙ67ʕ���NV=D�J�u����W�g�#G�^�n�6*f��I1�&Μ��=h���nE��fH�6<9�8�NCk΅Fo��l��B8X�QZ�oy�,�jp#�R�|��M��������䶆����3L|�$��X�#������K�&4��^�
��I>�!7eR��{r�np��=ݦ��$@��{I3ole;i�G����s݈k ��@b���W���w�Q�h�d<ǻqPfܑ(Q��Gh�k�_y֟�s�o9o+qR
�g�F���^�����b����hNJ��������6%���t��Qf����g�s����y�@D�r�{	 ���KU'aj�ݑg���u?���,F~M�Ӯ�r��l��5RJ�C-h��G��[�9�ΦsP6{�Ϋ���泪d(����d��GO]�'�!Q�v���%:��;���A(�"��16�m��	C]�঎8�-� �R2q}�lԿ�F�}%k@�ʚ������tJ�.j���؃yXh�L��]jKhE��Ԩ^F	�O�*�5�҇�Z��`x\#������>�t����&�Sn��W���Z��*+���*Ф=J��!����Z���HyJ���Z������3rd��&�+��M �P���6�n�3������$�����.��S������O�ϼ+�+I�4e��ŜЈ'I�\�!�ބ[1�̠��k���Kz���|���o��Z����9��1��,!-3�h+|:i�!��"6������1��|S A��f���?,�H��<eyٜ�[[��jK�$��Mj�Z^�f�FZ���e7.��@��E��'Gm+����צD:�Ex$Y�z^�SN*"5 z?,5x�����nK�K('Va����t��\ʵ���|����b�)��L۽>PH���mI8��[���=�H �}�*ba�T?"����S�^�2A�S��$I+av`��KUP�$}�`����ͩ��G8 w:l=��+���ʱ�K�8�.�K{H�b�P�W���h<�@uRЭG���Uk����]����|pG�8�78���gv����/�Uͪ�QK�k�#���8_'�/���_�Z�5R��D�rd����r> �q�_${���������} 1�t3��wb������rnp���vЉr�cL��I��SX����!j�?g���E��f�N���ܳd ߳p��_`�� �l3?����2�ї�#�!��<��_T�怘�,-�W)7j�uJ��ȇ_Nh�:�,��)�$h����H^����	����S^�f��	��jb�Ŋh��9� �T��E��c��۸͏Y�:p%��>>H�8�oP��������Y�T��[Ʊi��YH_J<�VU�c��V�S��!��[���qq���x�w���p��g�s�>�� c1��G��\��M&9<"�W�}t"]#}�OS�a�'��R�c�#�-��gc,�(�D�X+0L�Ik��#ۚ��,������&i3��3�Bzd<��Y�%!ou{>x�ۿW�)s�������������+*�Rj���o'�g	_�n�.�A!�^^ �T��^��Y���x�R��_�E���ˬ�`Nu-�횿�;��Y7Yk
�\�)!^g�W�eJsdY�����p+�Y$b�j����x�?!�Py�8\&>f��DWm	¢}&����cb=�cK�rk~�U�?��ͨ��N_�2�B;o���T����>0mEci��i�N�z�N�r��u�6�k���qD�K��k��C�g�L�� �|N�W��O�AL� 4_���M�T�m�j��D�s�P	���rg���@��W*t��.���J� �옄��ک����.�I�3�Gu5F4>e���'�l�� ���F�h4W�&�FM�qh���t�}��JT�>3��h�٭�
%��AH�/�:K��6����l����iO�8�5"�x�R6��%+�u[�~�G�k���A@��2�

���!�9�z�#|�HQ�����k3v-���M]��:2������\�ޤ�����1���3�K(�*-R�?�.�hƙ�A�"<��5C��v5���$W��G&d��Swy�����\�8щ�|�4�]�W���*b�Qu���Z��,�*%�W'P���I�N��Ƴ��N����&�Ku7����Y��@!��޼���	1�"g��N��G0��ՄhJ�h�~B�pK --θ����Vא#j:x�M��_ْ��9�C�i�Sp����G�Dx��z����Cfz�Q�x��d����cȔو����UBx�k�:_~�@�����@��L]��&<�)��aF3�c�<�W2kH�����3}���"�03���*Ν#�S��i�d�z���T[?�8w�Q�] �n�}�F4l�6�I\f���oXg	���1�s��0qgy�9��W V�]M��y���� R�H>��d	�Myh��P"0���ߗq&s&m���o�M\U��t7h����������Y�����j�i?��-|YF��^���'` �#��0pT�X����F�J���2r��Z�a�����^�����%e(Li5n��	C�+Zk�>{�X���ޑݟ;�Wg)����� �Z�D���
,cw��=�Z>aC(Hۿ
1��,w�;�k'�;��q���͕���S�@���GL}�T��q�8p�w���l�3<�q�٨�bXI�&�CO�X����@��y&���\�S��}����?�S�p�C��I0B?r�HsB��/ !���!�<"�����K����鏜�������;V��[˴rh�ɑ3az�;��|���R����;/�]��ǒZv	�L�VAc���\�=R���M�����r7ǩln�=�:�X���l9���u�:���'���\b^��Ⱥ����������A�,��ݢ}7�K�-�w@|����H5�f�~x_��h�`܈�}i�eS?#���+R�l9�|���  �M��Y榒,E��q��������Pq��/���3��}�\�7�_fM՚B�>������8�O]�\m�]Ǡ����1�����(�)̠�8��찕Є������eet`��!z>@���m�Q1J^�ٖ\��������E� �?y_ѥ�V]�����CP��j��a�6Gb���򿏘������3L�/�V�->��\��J@k�~��=w�6\�UC�b�I��cf�o�$g��?��J�Ԍ"Kd��m�a+�\���n%'Og�p�p<�i�/�����d�w�@�����N#�e���������]�!Ϭi�k���+�a.�U(��R�D*괴E�`�U>�h%���+�֊�weBg�<-���(O>�$���GJQ
q��~��5�&�;�2�x��m��+��[�����q�?�srJ9�I%{:)��b�!�DAf����T����f��2��Ǝw[13�*;���`��a�Ϻd�>�w�ԉt� t���!�}Ee
T!�ƉB1"HV���@���1��� ?9��`���&��m�q+����є����1�J-��!���ޯ+�;��u�_Y���I��>ޚ6i�9��/h�إ��P�&�޺���Kz��E�-~�O����~���}P��K�1/��N��Ya��o�����kD~N�;j���[��c	�9�n����%.bHq��,4�D%64F��'��C��~jt��K��ŝ�K�2���_Ϭ�X?:�,�n?��,��0��as�x�;�;H����#��Q�\.X���ZTB� �{AC0!��u��	�����b,��
�^{/y�#ɷ���A�To�W�?�{�X�ٴ�fhw �̹z6�ا=Tm�߲$��ae�L�N.d�Ge둥���v�b�z#�;��^P���U;�,��E�PBGz��H��b 5W!X�
v��Z���?��Ya�C}������w.�Hg,u�i~ez[�3\_�"��e����[<?E8'Z�B�~8X�[������j������Z��7#A.J_� �n���k^ j���Ģ��v��%v�܇.%�J���
��b����l �d���E��Q6!�O�4�%:�2��3����_/�I��"t;M҈L��6r��9Kyy�$����Ȕ�{�zH�-����
K$E,(�ܚZV-�����*��Vn��t����+�����1b9��L�"��Q>���=F'�7��-����A;��_� {�u&��8�e�Z̛�Cw���!}���+��o�	�0CA��a���[������� ���'��f����Y�C"���nCu���y�hCY�f�a�	{!�a�r��!
`��8����^1�t�����%����B�M��,��4��6���V�8�����(J­g�{�Մ�����~[%>Ѓ�ѩ��G���ɹD����i#b ��E�uw*�B�l@S�W2���h�f�>��C��ZcG|,����Ҙ*ە>K��T@'"̱r �.�Y�oVЋvZaFu��
��P�4�h]� ����\�4$&|���%�/d�Y��I�Q����^���жE���Q����������%6]��Q̅ߢd���i�+�:񫑟S��c.��+>_�Y�1k,.+�����u ���J�!���X%~�S�V�:�E���p��t��=��נ��ѹ?�Cul{eZX��c��֬!���0�p�- �W�+�@xu�͛���A��!�	�s"Ȯ����m�MΞ[��C��w�6��y��k�=��ns#����o&�[�G��=�E��_��/*�sg,Qu���PJ�r�Ӊ�L,I
���HE�s��� ��]�]8� �L��ʢ::/Wk���	�mO��_�O�A�Y.��[��?A(�V�ˌ�j	�1�~�X=ʾ�h��&x*��Z�i���+T�TT7�\�zM6�]���VEi�xC1��F��	�$����;�������sT�W��/Ʉ��
p� U�w���\i��bVk����&�\�"q�Ul�e�� D�LV�$ң'��
��g�"��(:��ǵ�V�~�������<X�T�/�:b:6�%}J���i�$� �-<��&\|����Vz�.|9�?�~y���(�!dߗ�PW�U���k�Ԛ��cx~�ƾ���yV�tՅ�����f��[4S��M3�|��y�����~a9V��xa�i���i�p�)h�T��GV���ݬHqX&��g �}�O0 ���3x+��2q(�G��@ʏ��`�o��������[���n�,+垞�2�[f�Y(@pđ�t]�犫[K�싑Jx_6 q�Q9|yE�7B�����5FU�K!l��: �����4��+_{�����+���>>���+V��K�-}Hi�(��'�G*1Z`�)������'V��,},��=�? fךeB��x��W=��Y9:#����7�O�k唕�!���@�����t5�
1�[�1+���i��+�d�=���!/0��Y�S�Q�ֵ�䎲+]68純�H�f/B)5K�IH� WY�� Q9]�@.*u߶��2f���#��-��1]��� �X�}x�q�C o]�˙��>Pv{�Ո\�4IE����o�n��z"�X��lgR�jk��U�"w��d�x?���4	(�����8�'G�Y�c�W�����W�6������R��e��0B�*��C6������Ϋ�'Ρc� _q��(�|��cc��s��@:&Iՠ�ʄ0����t���ݯ��jn�c��&�Ϯ���"^t?,�+
����oQ=��$�7Ƹ$�Q�	�B���[�2A#/=Y49Y��h��l�{��Q/x�bD5�I��"�P�֧������Sm.�}݄�F����>�e�|�ʃC�y��Y��~��=#���X��E��$��9U�h���cG�4-���t��[��ٲ[��ק��]fz<T��ܓ-��	yϲ���9�j�-���n"r�Ћ�Yv�4�m�w��
=y������긭|�K�G����e
�J_&�:��>�^/���6R*�j���b�u�z�Piy�'�3Zq��E�U��u�*�
�<�6h�����H
�ۖR��B���Sј�	�!��'���9�և>n�Ğgv�Ϥ�x��L�v�<f���jt������<���5�K^�^RB�D�;��%��;I�7������{�ӞK���<��׫�s����C�d\Uy�-�t��a�g���M�l_�No���^������Ã��f��Dƪ�`@(m����C�r-�~)~�!҅����%ct)�Hųd����0bR��k_-n%��B�������/�C ��m���,@=��!mDr�uRc����7�S�宻�#���t��I�C��*���X@��`���bw�����dU�œ�T���*��yx(U}t7��Y����n�#
7��l��\T��uL��D%H6��9k���j^�q�/��*��n��2`�1T�UJw ���u^��Gt�
��������6�y�6Q��
��������� ߆s5*d��8Z�	����}$��ʅPț���FP�����GBMD��jV� 
Y�;]Õv��w��p3βn��8��,��t9v��YYs���+�'���MpG5L�W)^,w�1Q�#ǚ���g�יavuF��E��aƫ�y��Gȴ|�D���n��2u�F�ì�ƀ��̬�rq�S������VҚb�mb�����l���RD�@���!�nn7����
�lh�7�vP�Y]cA/�%B��
Z��X���.���r�	b��h�Q����⺰�y����pb`�W�MF�K\T0��4�ꁢ�Nȣy�e����"��&7Ӱ ��@_0j	D^�g"D��E�&�/�Z0L,;��*���~"rXĊ�_�_v�.+��H���򅇺%AF1[���s�w��;��X��{�X��5�l�=:n,��=�}�����rHN��.���l�f��������	z�E�MW�_�\@;iW���q�6w/D�3a�@�Ms]�E�?���-y�+4T�D?H����)���]�:�]��\u.` �*3.G)K6ͨ%��L4�l��@I�6��&�7�� ��G YLf#��ߨ����:��r�u���� 	�%y��ϔ�i&��_���c��d�4Jq�#x�	���� 'v�J��`�D!�Mix��[l·�U�/0����g�����\8 �2�D+kV�m���'Ȣ�/6/_��]<��HC^���B�7�-�?�B��28m^�@��|�b���4����]T%ݬ��X[��9扆Ʊ����Vo2⺍�E�1�)-�&�&X�^y��7@P(<�Mv���.�]ĚlG�n�?tg+�p	�8>RK����Q!z������ 7[N 155D�&ʷ���b���kw\��ig����ӊy��j���&�_�x����/ѕE+J;ܷ��Ԥ��%8EDv�Y��\v��^��c�y���=di��_� y�����Xv4���"��-�ht����(� o$�㛭�q�Ï����Y���xg�Z��ւPPT��R�fq�e�@�ǘ@��4�������(���CNK`uvtIF�nL�'�ZD�,�łV�qBR�a����
�k�-q�@D�h/��"�G�����Ҹ{�-n�0���M��0����U���*U�x�t��d�
irؿ<�����R'	�ȅ�@١�@t�8�`�̴�V7��	]L8��=��(��B9a�^��0*��kql@FXK;B�$��eU��έ�-�>�xQ^�#��RTȿ��f;��������u<gc��Yh[(O�t�M;�������fpo���OI�t�m���u@���:� JPn�!z�|�GF�O���{���+$T��hp��%"�EI��ư�֠�#�5(���"��%�cNf�fkm�zx�����Ca����盀g�}z-;ۻ��-{X�[�WF �v�P�VY����P�р{�����Œ�=VBl0Ջ����8�Y6�Q~�٪٘[!FM&֭��e�҄�x?L�>������eq �
*���o��XW"uJ��k��yi�t���8����䝩�R��~��lb����������|����0�|!�$�T���kHtҦ�/=+3�]v�S|�
o��a�7���'WmV�����_�rZ�
�$"	@���_E���'�-PE�G�q�*|h�r�w<�hYH����9ȮQ��49(�cWAPV��?/.Z�b{	mgR�GN�6u'�X�k�u3k6ɫn�P�0��S��ͺk M���Y��+��p�]=z��O��S�[��Kx�r�k�'Ɓ����z���@�I)eL�6l����؊D;Nf���u��߾��P흰�a��9�,�.T2����=��bk|6'K)Y���j^w{��_)R��VV�a��Xs�i��Ezuz#��w�1]d2�_c�D���ls�w�z%L\����g�81�K
�VgWA�֛���^��: �j!.���)�ǌ��[0�>~��
L͟3-uɟ�^�ksLc�i�8?l[��6��蓣�?������NR�ί���E�2췛�9#&��l}Q�����?ݲ%�����Eس������2��\�e�����!���&s�WX!G.H�V̮	�T��'�i�5�`A��Qx!J�D��֡r)v���� ;�s>�`�Hj�M�p��h��]{G�xS����<O����a��n]x/�~����lA2|�9R�<��u�40hw6�[���	�n&�M�	x&y�D��Y�s@�J^�Q݌w��-"\-�ʛp�I
�����G��C�lc�i��\�zQ��MS��PM?j%Y��/�%b+�+<��25�ռz;�v�~%T�>D�O+���;���r�Î	8\�
Xn�1�_�it��%�6�� ��ޏ �X���[<O�����feCr��EP��W�g���.��p��"Ah���S����|V��Y����#�&�?˸�8��bDwr�Μ"m��
9|�_s�l��k_�!|(^-x���ݴ���z�� ?���KBX������)���\���<���wڑۻ�rS�*���˗�7Bͥ8��;qL���@w����Fmj��QT��-w�0����x�>%��!4^�z��*6ᩑA�q"/o
��(�u&��/Y���+���3���=i��W����2A����o2OCccx��d5�wJ�Xurg�=��[Fu�r�ӴK���ɮ{]^��?�����8�����k��"���J�^�Zs�V�7��^1�{s�lLBnA�S.��۠���ޘrfg��o3�_]ɸ
}M�����4�}�)/ʟ�]��b�t5�r�`S��l%*����s�SLvr{��n�I��^f��G��7l��`%Cm��i�0GY��O�O��D�3~���'�݈�.��Q��ǿ��&/���؅z錦�8z��NЛ�0`܃1��>����7oK6��f\8*�*��n�K�����1bb���j�y�u��~T9Ĥ��h=�P�:g~%�~�t�g�¡`�nz*�s+=���2Ǟvl)����đ��L��}#<!�?��7�-�n
򵔧+��pf�x>Gz
yT
���ޱ��y��\�7��)o��sMNҀ:"�������}v7uf�3T�F�r	~`��ͪ��������Q���O!��$�X��m��Q�ޡrF��i�v�cg��Y6�/{�R1ډi!Ջ������X;O;!-���n�x��e��+�D���Vė�i�Ǘ��
��β�QvR8n��x��lR��Ռ	m�g[+���ޣ��kEɑ�S=[2^_����b��M� G�}�Ǯ�UuQ�es�<\!d]�S����uu�j'F�po4𱑕�Rrx�vs��YT���(0;��]]DQ
�2�,U�C��s'*V^��do��m@G�\�r���[�#- �� 	;ﶥD���-a�~f�-�/�|h�F��hY����N.� ��\��/�.t"���2/)!�o^4#=�,��K�}��!͐b�+�7��7��:�L��1��z��l`L�\Fa�un��^3ݸ1��2hχkZ-����g�)�k��V��I�N�W�����N�LJ.Ct�K<����Z�KvrЕ`�I�J�Ӹ+��Xw�pr|��ѕ&@�W�`O띙����s�vc?�h�r��q���-�s1����P�u�j�p�S�ڦ�pys6�K|���z`��OyE����L<z��
9I�R���|�#׶9?E#�x֧�@��(Ht�goǢ=��x��?8M�u��[���{B��j\�h�[I3K�PX�LUg˚����d}}�����4���L���(���kH��-�Y��A�X{+$�����)rI�u1��RЗ�D��)�*�	�
9˭���Kf�<b]��A��Z�.�v9AEҽͬ�����/T�|a�@�Y�fe�S:ܔ�;~8���]!)��8�K��`��c���B8ԣ�Éi6�B~+$�2�c8n�;î�t��rr�P/�ʷi]�glp	2���HtG(�~*HA���Jt�]z�ղ-�8�� 6DGk.+`��xc4
��v��X8.��F��"���9Pr��sE㥰���Ͼ/�|M�1ZĻ������!��TY2>�X�w�[�i�_��"�.j���F��j���M��mI�:s	���f��H��{F$k������5��{e5��ۂ]H@N�.���:��A���|����Xy{�^�U�$��]�a�)��ͱ��"�z5������g�d�`��A6�C��������)ܖޭ���ʺL�	�[4�ؖ��E����I9��d1=8�35w��� ��q��RN��V߀L��์����p#OFȹ[�Yd�:j�8<:΍���?�|�U
�CȘ��>�Z5��`��pܡVˎ�owf�t��e(��6*�K�*����o�)Z�Ʊ^J��&?���<�jʚ��u~���^p�s:���0�ݺ������Z�,DkfL�4��]|��R�HΒ%�I9� lG�Y�J�P�4\x�� ;���������K�U�'�s7Gb�h
��N��կ�}��%!��,���¿�c�ḧU|�X:��
��BH�ޱv�x��R���0�}�<C���ET�*�U(6$��(|����
C��s՘�]c!�xgr�u����O��5�����-�j�p���g�̳{MM�sQ�4�KI8Z�"F�wD�=k%ϲ �4;i���G�6�lO+4�j5%m�c3^$5LQ4�$��H�к��I�.?ӱ��e������cD!5v�~`m�ۇ�L-\�'�E�t�;4~�	V��g	3w��Y�;��g��� �N�9wʒ��k�le�L��x|饽��"R�ϴ��3��h��a�#o26�x8Ž����.�s������-�%��W�F���$�<[�itޏ�p��aQ]��r�GuM��E���vY�F}����,L�
3��N��Bqp!*�C�,P\����S����t��aVՎW��
66������X|��N�F-��r�Ӡ��E,`�dRq�~lE�3��~�}l!��g��٧F��J&~�hg��IMK"K+�T
lg�s�~�F�0#�iM
JH9G�z[G7�������u2_�U~N2]�N�W��t�V�P�M�J�����X2��b���'P�)��rՃ�̆��vOi���j�-W���Q��Ӝ��y�E�>��f=��Q���W)�T]���˲��.�T�*Xkx~v���6*�ʯ�mEX�F���8��c���Ȣ,�PN���b7ZB��vl��o�;d3)t"�La�[o?���`����.�W�$ �x;s#�q2J�lD�.(�#üL&�KbrO=�'ֹ:���f�Mp� �ș��vhǰ��y!\y�Q�5S��>-��Aq#��_���ٜ��/F\n�AR���"�ӏ_���As�7��~{�w\lˌ+���Uv�F�'��z�����A^&rM�o��p`�<��L�+\6��K,���,�*+w��~d� $�X��*?�@ʻp��w�J~]vHX U��DO�p4��$s��Ͼ��\���,@y;�̂Zam����3/َ_�(:L��+�ؗ�S6T�m?��@�ߝ}R�T�u�
g��u4a({�} fA�^V�K�	EC��x@}�Mխ �F�Ƹyv.M��Ǳ�x���Ϋ��$��i{�:�gb�jw򦻟V�2J����ǩ���K��I�T�4�h�j
�?�s>�G�`>���e�+��~}�`�C,����6�
�Ձ�U�M����Q�M�v�D�zD~C3`.T����C/5r-�d+�{����� �T���px5��}zf�A����,��^жP!�K�~l���:�f}�C��;fy���ձ/!��r=����U��������ƌ�;M�i���Մ7�{p�J]L~�.>������W�ut���N-��#�q��u�ƞI"g��3p���7�8�IM�R��:���r��!F�?���m�1�+�$Cv%U���ʩ��J2DrM��`����٦�O$�E�DB��n�������ؐ�����_qW{�J's���{Y<Z-9���$��C>�߳n�L�տ�p�.�7'Pg����>�	�>���6�D���-��r�(�BN8�6�����f�ibVTJ�e�ٜ����W�~���Ƃ�FT�vN ?�Ȝ�����xmtJo������5����`�
�[uYo"�^� �����{�p���H{ͦV�Ns�&��T�mn���ۄ���g�������{�'���?w,h��lf��#���q0y��Bs������[/���_؁?���4��a��{NΜ��,��F��Fa���(��P])Kk{X೔<�ۏs5���d�?�(qH�x�ɡ������І�X���i��U��-�V*@G\T9� ;���MG��"ʄ�T ڥ�~�tw�#�i�J3Ϸ�Z3vy����$'����MZ�K����s��V^�D�������=����'V(1���fԢ�m��U��M�y�d�A~$��tm~���:�v�ɱǄ�}����.�)N9�!MfQ,��8�[.ׯU�U�Y�;��r5���H�!�#h�'�$϶�]�EUIl���A�z����ϨA���70tH�������]U�l�7����AXuoT�Z���*�<�& ��b��F�1]��2�g�fʼ����;y��Q~�Y�(Rq��ڇǗfeF,���>�4&#�� =����5��L��j+4��&
gEք&��uȌ�7���;���sFx��XT�^���8z膵]@D�>��r������$���iK{~���;�Yc�Mo0�����b�D��_�/���7��]�ƻ��:B;r�[Z2�`����#W�Ÿc˨Z�	i��������c��y��|��ҞA�3h�$� 1��Z��4|e��^sg��no~j�6���&wsg��a�q�}��LVf4�a����M�c}I��v���쓰>��ʻ8�zv�Ύ��:P=[��EI�
�������jsz��H�O���5�1�kuB��BP0�ŝ�J����X���OL��*⸾��R�b�Ĝ&qɶ� .XQ�W���z�t/� 3�ʾ�!^ɀ����c��/�C8j��>���)�[���3_�yCO*N��ZӡE�9R7�/����|R�2���ۜ���|�afS�#��Dȿ�y��}���VE0O�\��OP��Ҝz���m��ɤ��+P�¼�J�h�M�l�2��K��fWQ�т�Hl~�9�����Ō��*��BZ��W�D<z�wO3!�#CH�KD��'I*�A���|��W�"� x���ɓңi�lJ�ͫˠı
�ҳ�)�S�u8`I�&��3�zO���G)>W[���~�h	�O����C����8���z��rH��n?xR8��|�
�46�<��/�/}P�ȸL;� W1'�i�����R��x�c��^��Ҿ�NMQ�֟S�hm��x9�o��֙ r#h{H��(��
/M�iK� �i%�b���1�+�^�e�cb��{ _�=>�k�wv�1���������'�S<�m�6%s���cw]��]*ԛ��"N��3��uu\n{���M���}�T'2�N�� �����O��uXC���wkY�A1x-t~z�e��O�%X�鳁¦�QzZ$�M��M҇��/�����=�Ӕl�w
!D�CF�풽�EzY�:����3S��s5�Ց�=<�h1E�ћj����5r�J(��S���%[_�	ڈ=F#qյ^��I�l@�׹�x5 �4�����P���eřnA�;q����g�ʂpS3���^z+��G��em�a�R�>���Q�P���.P*����;p�wO7����1�} ��
QB�F��4��9T.��+֧6�]�ƻ�x�s4L>݆$)�8��+"Om�`����6
������3՟%<r�il���bʝ{]j�[L�j�3O�{dm}��﫾N�V��R�yu��i�S����g�*X��Y���蛲dl)e�������;�y-��$~��Hĸ1������a�M�&�/�'yLck��7u����R��(c 5����de[�����={���gV9԰�0��]H?�K���!�œ�W�*<�N0�褚ٿ� ��O�^�����{*�n�����H2GS���SSx��#~��T2Vi����I29<�.�s �-��s��i�Ze��Q���^y���%�3��.�s���g����\�':�VV��D�ˏ��R�F�S`��؃��)X/�g�SZ�_E���ai���S�����8��.\:3��������ٷ�@H#ک��'U���u$: �ɑ�pۻ�=*��"`K��8��E��%R���EB�����â�=732��'�KrE/��W1�A�+B�b�U�eJ�c��a�Eb<�I�4�L��o�Qcr �sO
SG��y�U�j:��yЫ��.�`f`E�!S�����$�D�� ������vFZC����0�¤?((��T�힘�>���Z�o*�O�C��`��~�e=
�` ��GLE����ŕ��&��Ȍ�OM�6���v�%1�5;N̑a3�� �0>����ޅ]���6," ��GQ��B'9�f1W�ս��[o��-��*��+�R.!�t
�~�꽒�;)�)���
.�_:-��C������"��g�:��`x�-k�Nl:j���&���?��lua�.�Y<���";v�u�gs\�=�ſ+����ɫe
3�RmC�iMH���*���R\Hsż����R�x���^��Gj�c�4���M��G��g��ĉ=�x<��Ӹ���\�!��˙�\�ߑ��ֵ���槓��>npm�=���b%��cIl�L��jK~�o��H)�:b�D�/c9/�w]��?C�=����Hή��*��q#}U�]@�K}"�0ؒ�q����7g�i�#i����aZ0�!���D�Q��	`����|��9�罕b@ه��!�6;3�᱉�� ��ެv	hLgc;I2��&� POc�z�Lae9�ҝGO"P�ȉz�'�!��1m�{�![��ė-��1�\a��������w5�-n���${Z��׶:����E�����sy%w�b�ʶ��GV��Ջ��X���x������^7���v�A���o��A���Ϳ��.�,��W)4%��޲L��2�5�:�U9,{��5��c��FM����&�<�ٗ\,���1��X]P�H��W�wu3�H$�V�7
��|�oe������n��>�,���)��? o�|)_�y`���h{��
��ב_���{��̌��,�������D���GqE�mvL�!M>� f��m
��4F���0aSX��.��� ��kH��]�bދIh��O/�Tk*�8yy��^ ��$y����V�*A{�\]�;f��+f��Wi������?�Y~�Mu6�ށOц����
��vȕ�j��(n�� �#��+�w�B�F�7��Tæ��Z�F��`���o�D��R,I㸩L*8Ao����+1�
��+��$�*�	�~{:>���E��
��'��1�*t���8�M�f��B�4p������6Z~XQ��00���d?>ʡF��FLF˫'@kFRB����V����M(��>�~�����(�;�{�3@i<U�Y���s���	�ER��d䄵0@|(g]�ku4����8+��~��w�mi����YНz�Y��[SR_��i�j�m���`���ϗ'� �&$����@31����־t��l0�2M�_^tS�d�Ț�0�"��
!����b!3q
��8��Q'��43�I�I�q��=��k�	-�+�a�H̿�&���]ɳ��7x�?��Gw�E7:
@UVdz��%�Խt=�	$sۥ�Fs��%���G������u��:�����B���ϣ�����%����6$Xd��hG"�\3�E)���Rj��9�o�/4�Y����B5A�#�q�4i�����a����y�w�0䑀�W��R�1�
����Hy����b���f`I��e�C[﬈:U�J"P��z�щ�<'���R���w����AG����Ċ������8�����K�d�J��|�MYⰆ��1k�}����y��̩+�������"~�{zd�/!��Tm{C�B8��|>���+L�I=[}�l��ZC-Cz�I8��$nUq�������l�����_6!��~�ʔ�A�+�V��wf�)\���۩�J�����?�R�S�@��F�zD��7P�*}����N��`7l�]���ݴ{QtU�v� Pҙ4��:�H�V���ۑ�Xm;�_nt���&����ߤ�l��g�g;>Xf'V�&	��($��y���2�/�"������
^�%C�%�� ���`�-"j<���I���e)�z~�>|���*H0���UDO{�ټ�I �Й�H�Y&f�>;s����b?��8����j�!�
��v���DA~�[�*ݭ�u�A��@�F�|=cd6&U���rC��mI�d/�ar�q����7�*QP�媽����ZC�)�&����Ĥ=�x*�%�A�r_L�
H$>���K|����C��(������m����K�r-&Q�3�f�7��f,ˢ��IY&���������a����g��+���z�,Ú���ϳ�;�:�a���E�1�񅊚�2�
7=Z@dz�,4ղX"���o�����R;o� ��{��J��Q�Ѹ��+>�K`����C����m����U��(�0^f�:$����DA�J�����#39�ƙp�|�$��>�M�Cg��Ԝ���CAi\F8O��T�q.Zb�z3
6v:b��v��C4|�����r3x� r�0�Wj�F\hX���@�ĴaU�Pt����J��T�X*ᚷ۬W���mތ��6���1%��#�i�FXI�vq��#�Ē���]��3:�M�%X6���	�!~�h�	�����o��j:5�;���{(����K�o�(n ��˓h� 3��ל��e�� �4(ʒ�Xl�y���2~���=jv%6..lu��s��?�i&b��e�5)�c��yecggOK��Ȗ�_c�iٿ~&����S��bz��/�G9ή�-݇��D��l��|9����8. W�
Q@�[��G9A����	2AC�z��#{&J*�c9LH���>� W`������#�Π�JI���r,�u~�t`�ʙ!���\���t^aځ���fd���j붦��WwI���8Hϕ��F`+��	w�fz"�3e�_4�:aQ�i��,�d�x}6�x���{Q�m �W V17W|�O[�)�?��mWw��� `xѠ%���4��51)üM14��@vF7�gNf=�H�I`6~�j�%�����b���_`�?���
�M�8��Ƥȓ��Pl���{]�-�8��\Qe�Їsg}��qA���	f�`�f���Ocj�*�F0"~JS�͠G���WE�U�|Y3T��ڭ,�N�U�'�-���{���1Z���mK��0��D����	C�BEjW��iw= 1����^k?7ƅ�~�5U�����C���'�ێ���f�>�P�\�a�����o�����Σ�ʇ[}Kwr��%+	��%�Z��j�Pn�gԓ���n�4��z����S,�~D��0@1dm�`ͺ�M�j�	ᩮ��� C���q��nŃ�XcU���'d1Jf�����>�HĠ��q.��\�/�~1��%[�J|��JE~(ۻ�-c�:<�U�~�$:�<�2��������է,�-����#it����!��|8=lxr�c"oÅKy�R<SpG��
���T�S\�B�
4B�v���!��ܿ5�c��.�_@��E\Zl�?�����3�̨���Uc�m�wN��yM�4&�aJL4�&g"Y��;f�q��(���Y1Ǝ�h���cT�̴��J�aIM��V4����Ǧ��ٔ���x�X��������Mv�8a��.\rV8ܫ�%'7���nF�����D
��2{�Ԉ]���y[��A�*�+�����L��t:�}1ÿǲx�jma�����8�e�#�J��j���f�v΀�Nk�&��?�$!��^�:k2��ڛ�\Zu�<��(�C���6����"(bˇ�'�U�$`��^$^�or(��3T��Ʋ�nl0g�%�Yr�<�+��f)J���`��S�}�U	��Z��Fw�I�(4�F+�#��7'�>KZ��a�����!Dk�A!��S�F0�V(P�XtT�+�/�������ԯ��ۚ���G-�@�E۷��/�U!�:eDxw����H����G=����Hu(��K`�d�U^^a�
��U�xy1r���۩��VQ,���c[��mV���بJ������3�{N�Y嘄w���s�h�[�P_�I�ds�D���%�v��<@���e�+��*��h,�-l"����QX�/R0��L,F87���,RMǖ|�_�9̖k(}M-��k���iPыa�e����At&Z�v�
��8}6O�$�o�Ȳܓ��b���/F�BO�9݃��YC�@�3�1u�������%{h�u�wc�y����x�n�*_H�m��OO��1�u�|J�/E�a���]��	�Խ̫���G����[Żt;�#*i�W#4x2 ���Vԙ�
��)����"�_>�Ag�cD�Lh������z���{:���\5��Y[��������E��lD��b��X��=�:f�Wm�>��Fr��:	մ~�M-A$E�s/�K��Q�Z��ߍ�鶘��ʡ�>�#px�����A�j�a����>�Q�G�3�:�����g��	®W�zh�Ӓ��9�'�IJ;��
�B�f�v��� ?*�A��]��E=��zgmP��WW-?ql g,$�7z1� ��߳����ʌ�>K�Q�#7J�H�	P>^�Y���%p�yv�#Aj�x���x��yFV6�@��TB��F;�2�0�X� �d�qikD�㳢��Ds�NoVƐ��O�����F�j�[���"n����Gک�1r��3�%m��
�e�����h^�n������s�܈�sf`"��a�71���(�J�p
�g����\A�u2Ds�Hn4�]u$��T_͹Ŝ�٥9(ƺ�"@9�D��a����_J
���oe��{����������-l-���Ҽ��տMN2(�u߿}�27Χ���d�����"�aq�P^����j������;�?��1y�.�Kt��n=��0����l�Ƃ��?ezp�D=b������QjKt6-���oMfO��{0" �\~�m5_h��˔޼|;d���Lp����?N�VS�^���W�$��&��v�)��v��Za�iU��np�j�hV����0!^��i;xeǲj��0;�x�ebvDa�K���u�f���v���	�SJ����Ĉ��%�I7m��^��� e���@�'���K�jQk�NWê��e�l�:��)Po�G�Q��ٍ5�\�I�Ț��B�|���ŒG��=�eݗ�d���x�ũ�DG�h3��S���B V3΃�PÛ��0�&
W�X���QS>!����0�Θ(?XINп6��7R!�s��(�l�k�,J-��{��:�ː�H��KL��`p�~Qv���f�����2=C/?xo�I_�����J��Y�����ǰƼ��}<�a(��e��;L���Z��J��}��S�U:Q2^�m�}<j�Rfr`wm,L-yMÆ?�=�j���d�X�]�aL<0��g���ہ�B�EP�Y�k~�b��C����.��Sb�s;!�f�Ga.����	�c�-b,1�P1-�y��D��|^�"�{֨1q}�JD%'{N��XzY��U�tq|e�t�5�p����2��Lu?�'��[(���;G-C?q]�|�2��2>�XUFݿ/�,�~�Q0�S�CB�м1��wO�W��EBi~�#��ʎ6"�	���C����J�Çc�<E��fl��(�0� �"�{S������i�s��*�BT��	4���a\?�&q4+}�]�H���_�?�%���g".�
9���E�
C6;t��A���Cǚ��sm�h]+I�w�=�Y���$'�����G��������d�3`�IV�cz���\RϔX�4�Cf��]����}�o��|m��F��bd�	�j����v�pѶE�y�J��ׯ545f�$	��sa|�nJ����ui�W�����ܜ�Z��M�8ג�,t	�j^J��P ϑ Sih�c,D�̙砦&
Tdai+�:򶯂�/�8Xz#�阹�}�G�a�(REYvĮG3e�c^�6p�a���pT1��*;�4�#w���x\6ّ��N}��g���4����ylW���ߴ�T7���"te��CX��4	&)�]�ᩥ2�4�Or�Aę
�T��`�씷���[l�]�Ȳ��)�n�^^���"������[�rʽ�̋i��n�ah`A����A��O�>����d�y�.�-.J?�K��j2�D���;��Qu�\Z"���V'W.J��Ҕ�.N�~��������9�YD+Y��������CE��Z�-8P�]ì�e���+%�����ܡU��i5�0&�t����C���>Y_-P��[�h}Sp����2�.�r�ֈ���ua������%Z�Zȣj<�&Ғi2F�\��q�W��Z?P��D�S�>���n�f!Y_�(�{Y	g�,,��W�����!/�1�9`~k��O8t!��%����9�i�-�c��HsFM����Jѽ����*�5�`�]ۖBa<52IM��J=&i���s@���U�i�)N���6n�*����E��8Gp�˴(<��LB��q�i��r����=~Z�*��߁^�P�Kǅ���)%��P.�S��1O8
-6;x�By�Nf�\���iꛇ5�.UǁfG�]��.
͘(�PS��
�8׀�W����8�hSx1�˃�\ErN#�.Ǫ�ǘݴ_�c�' e�X�tS��s�1V 5Z�`e�Cka�0ZS�F;$�,�k$��\�H7�^�ht7���'A;�Ϙ}��R�WXҿ�pX��]�S��O9���$�e��Q��e���ws�j��{D`�&~'^�:��%
Y�P(���R&�im�&kK��ypEVs�iB5��@����l��i��3v�5��yzRf��/Ɉ���I��s�S�>i.�>�?�8�Y�v�����NǇ�i�QL���H*�Ӈ��v�Ɵ@k��_Ĺ���BSl_�KfF�݁}Ќi�CB��F̥�&��xS(/�Z֑k�,t�����C�[^�L�)/8�������/�9��
��@�xٗЉ���Km��uX-���@�R_uS����	�!nVA}4�{Kg@43o��������a��vHxڭD*!X�������U��P&��y�5��y��4/��+��u�K�Ԝ{�����` ��Cv)k������e����.=��z�l��]���f���&���wv.|�䴡 B�,�������$6� �~�5`�N�W� �u�qu���S�J;Xዃ���+B���tq�����K��᱿�>���W�7:@`8��˷��M�V<`��w'G]8&��gT��o���_zf�4�~ŬCk�C�Sh��"l75?],�*<J?M��iEe؈c���������f����%5pPh�c��	�/�~)y�,��������x?��+0�+wZ��^��4z��O�,�O�Q��[X���(v�]t�����u�A�'�	n��5t�Y>3dILL_#������!����?J�cz�7X��)qo��0��Mk�!͇�I���O;�
,=�h���p*��٥����8z�r���&gP���e���pg6����q<ْ=���3P^{g���
���u��] `~9�Lr'^k�
r#[��N�3�B�j`��A�%�Œ�[�A����|� (h4��vϿ��M��<��W����uK�V{�z��0�, {�:�B4���{�j&Ea5�oj^�>�d�1+_+�~�;��_�����iC>w��W}s�����qpNjy)#+_�[���۬Ȣ�S���Њ��������$�<�#:ƶyz���K�7���^�W�_�qLj��M-�b�W����U�~.�_)�Β���$3���`95
�z���R5�k����K}��w�c��ϫ:=^�:l?h�Ք���\@Fu��m��ZIrULy�P�77��`;@6/GȟY����{��L"�ާ�
��ϸ5�*Sń�{������ً�!��6�����0s������6P���Abz:u��`�mx��d~�s��d�ďP�;�jw�9�^v^�O���D�3���ncO>yF��G�w�_���`(�(���H�0 ��TV�6���uaT�4�U/���>`�nO��Q��jY�P�OxI993S�a�չ��B��"�au�*�C�
���g=������Q'k��u@AՇ�&���aþ4C$�o%f�U{� ��N��@�s�G-�~�4���Kf��=��@;|��Q��i�u)��Õ�~�t!��J4#z�[~�c��Nkb�p�X�f����p_���J��8R���t�%$U��/�_��t��u��L���f#zĤ��(e_JvU��h=��$�Ңvۧb4����vD��O���OeK=�@$እ��I@���?ȅ���r�l��v�#�Z75NU����I�"F��V�q�y�������(�ہ������,l�*� }ʫ2�$'z�/���ia�E 'N�l�Lt�����@P�a���~���&s����s��^A��}�Aش ���
��=FC\�_��Z��:�������p����ɐϣ��G��SZ8q�¡��7���Y7%K��z�����-� dC���ve��z�R��~ьL��S�Nd�%aUUNc�9"�.U��.F�L<��x�6k�3S;��Z�PP�z��H�o����ګ�ytUg^^��_ 8S	E:��!f�,� �}�S�V{m(��{*0��cv��Q�;�Z����9f���hw�)�Xî/���F���]Omz�A�Jf%k�:+R����pP��/⦞hk�:B��M�^�Tʒ@�������D��+�PIs���]�UR������?��Y�nno���(�uu��26nq�v��]$!ho{)+C��{�\�p�+���/*�4�i���J��!��w	K�0eYq��s�73��=�Z����Gh�d�@׭̇��Xl��<o��D:�~�����82�������į��tJ���Þy�L��+����Uҩ]�AUŢ��ִD�j��r��q�h��5mpM�`%,7�L�^߰�5��L��=Es�L2gj�.n��J���ïҪ[$p/X�JR��}U�xNIZ#i��(�tAN��<.�����V�
�U�KT|hׯʜ�W�KԻ*�rR*���z#?������j�fp����}�/9����k�+�(<����)�TÛNT�&ݛ6����
��Q�)�F�T����'�V-����;v����b�$9�s�p�j$�����H�<�i2v�~D�����k�=��O׺캦�@g �gf߇w�����_"�԰eg\$Lo3���x�j���t�ۗ�d<">A��SS�T�0@�Q��P��f��G�j�6º�Ҏ�)�X�"7M���)_��Z?v�J�S�P]�/��I�.S�c�%h���q�nAq��2�tPC�06xYO��͜AtӦt;�c�zbu�ǃ��A��%�W-��C%b8F�B��@��cz�y�n�������S"=2�Z�=_�n�]��p�+� .�m}�I���_v���~����	x�?'3�)%�W�ú�4p&V�����yu�t� <g���N;���RzR36���4�D�I/��btr^��٦r�5���#�px�6���UQ��O3�l�ܱ��.P]0�@?t	2�~�U� МIq#w�!b[d`���]�#�_��@ .0� �锄y�KM/�x咧q>��U�B�)��M�L��-R��n\�i�6V*i�68A� �z�X�~D	�dτ����h���;V���0�8�h��c`�`��=�"�#���4�>l������E�/C=��xF�|�fQRX'��5���|f��8�U>-;�VK�?L��'J���� E�����䌬]T$�e��p���a������`�.�%XZ��~��W�W�W�d��[��׾dZ�����"m3K�޺n�ܠg����W�mw����R��y]��Y~�LQ3�B����R:�л�㵎��,�-���K��{�r������6�:T@��= ������T���g�+x��ێh`2�*�#�?#UR�?���i�o�xaFn����Th�ʵ����7�Ql���:���u�4w$��,͐�a�?��e^H0���u�� V���C[A������O̔��$��š��T;�]��b��Ь��zS�p���e���7]�I]e|d�s�e�9����jX�4����@Q�ˈ��8\|o��'Z�s��B�F�ۻb+���(�ֵ@���xϼ�K\S���*�~�[�H��D3Y	=����m*���u��n`lW&w�캌gdŌ�n+�l1_�=V`�"\n����B2	�xk�^�Ƀhg��,&�U�����K}���� �
S m�	$��C���>#z�#��b�@�^��9���m>d�\�qTN�$�  �TϽ�	���߸_IW��U���/�0��)��{.z��z!�J�.k�R�w��4o%L�I�揟ıx���f�C�Q!����	=����{a�G�E� a��l^��n���M��ϑ0�w1_e7�]��b+J]��m��IhA�F>�;�D{��s�l���b��#g�Bz�bs}��`#mY����J#绊n{,���%�Te���O�ם�3�~y��݁nz�ޱ�16����:��ؘ��G%4]-���]�0Z������zh�2H7��fy}w�	��(w׶���>isS��Mo٢�8��4�"�$�G���-�k�uY�T>�#�"یs�u�>����zK���g�y
��q4�&��i%����Z�}bU�{��N��a�{�����}�^F�6�����PS���;�b@�9��^[�T�U��wL�'Q��Sj���Cv�e��eZ���HW̮R˶Ie/'��"�9��O9I��=J�� ��4���$��[mE��SŎ����E9�:���U%�Z���H�@��e�آ(����6��Q�~�)F��yb��o���ʹ�r����~�l��k��I�Ǝ��)�t���q6��4��P �o����#BT��hl�B+�!��,�F�&*�c~q��UV�X���<��a�_�~���H'*������G����J$E� k�W)a�
]���c<�e�s�軥G��1��k��H�U����DG6���rLݟ�I�Z��d��+j�"ە�U��3ٸ��Z+�n�'د)�f'�zC!U #9�+{ψ�a���g�t�,@��>�c�����L�SRYW��K��!�������_�W3�����ۖ�����b�0���ː�skh^Jc%�&�a���3���6�� 僻z��UPnM ������q+��5�6�v�f<��sp�W�6�
�����G�E��>�#;t����p�e���q���� :
Ӱ`�G����肴|I���@�����p|��J\hY��@iIWvF�Onx�����ˀ����m'��hCș�r�E��R|�%1~�X����`�L������heJ����A�m�XX	�c�p�L�ш6b�Zʄ���r5{RuK�}=`T�����@Rr|�U��=�Ȓ�;~3�H�]%�)�Ԝ6�aT���f��T��6컵�����Ь�淌�S�'j�+�� ���	B�H�3̖[��)�!ɭ�7��T��%�4��Ĳ�R%g�3($V&��(xJW�8�,y�%�������J���s��}3�����3��L~����d���}"�u���/���RHH��R��,G�{�ǵM���qE�x�T��1-��3��F����� 0/�I���(�c�5�j��Jx����Ph����?ttWM�6����w�����n6�Zz�s�d�[ U�B�<�>W�毷���t7d=o����}];.�<�sB���G��vf�}D�޼5}��������-BE:Rw��#MV��@�`xJ[ b�`�P)¯T3��o �;	Jqیiz0��nNa��3�"��n�_BJ@�?�X]ȻLM�n#�-{�\�]<�0r�� ���lz{sr(l�i�t�"���T���0kK긶�\t�D)y_��KC�7W�dd�jB1�D�6�7�1[�X�?���m�<b�G��^Sd1N��bT�Fb 
����
^�Az�n3<Vvz:�Ƣ˧mм�v�0�:)9�Ҝ۟��ˌ�������T���V��A?7���i�n��cjz��<e�S$�nU3d������$��܌�����>��ýf�Qr����o#K�����WL�������*uz�*<��l�W�>ԪB5������h
?m���4F�Y�x"C`|�p��`��*Q.���N8qD�f����7e?�����f|=~k��#tjsh����`�&c�^ �d���Ù7X�a��-��B��LE��ޣ���p2;�4�[h�YxV0@��(�%�^�xh�K�� �(�;5$����;Ѿ����)&
^w��֫�����Q�����o;� ��A���xt꣤���_��hٸ��?kp�,�7��=�:'/�t�`#�a�E:�qTo���ͳ�ʎ�:�"w�(�S�P0�DZ���0/-Q3jÂ�c�o�j�8#\ݩ����f:��@��#���.D_�.�����"�'	�)��R��@R��fDwi�����֚j[�=ecd��`� %I���
��1������ ���ڎ�,�>���y_.͚p�@�J�ܐ2�D�jU�O��Kwa6e����
��*��b�k�;03�<JqoLv$��������n8fyu:}����o].�G��8Z-����a0x�T�t��.>���"1���$�Wdgg�+��'Ø[*���4�%�A�7|���^av⃷��{[����M�~>�T���B	H��3�tc2a4]"�Eh�m�e�Pp}�_���p |Pu�=B޳h����sfM2�p�u�aDbo��
��K|�δ��������B�P�#���{es@��ҜZ����	ʴ_�k�{P��:���a�lO�t�/EQc����4U^gvm�����6A�k�+�NZ��7�������R�  
�k�ٛɹ
t6�ջcH�_�'	{u�V
_!��'1j��*^ۓ����D���ߜ�IG�w��Ֆ?]��^�m5��k	u:gw[�ע)������aSc�n�qP�]��TBj�&`�F)�m��@ƍh;�3k.#�(�����5�'"#,���~gB���!�ĝ���@,~I�����`� bg�ZLj�-@s��ăn�+T�4w��4��GI4���j��X��waK����`��'�Vf����u0�q�kq����"����ܜ��w�nO�F��g�}ʮ�N�zw��$����ut���Bt1�! �� M�P��'��R�F=o��:`r���a���i��]�s���DH��V���5�Lᖞ
�
�D�P��y��,`��[dY� 5��h����z�;��q�]m��qe�8�fzO�Д*J.�m-�ߝc�t+�ک�5�!��sC���t��7R���M4@��k�(ůu�\�	�������ѹ��0R�f�jh�(��Pϴ
�Ѭ���t���^$�y����E��j.B�<r�����%g]�c��D<������{H��E�>��	�@�a:,+XG��t�����Uu��h�}�	���!x�`������0�R��׹G��j�\&�=	W;�A͉�i��Ѥ���f�h��3�3�d8N�d��u[�mf�I�5$PQ쥀uXB7�����Ԏ<��a�Ǡiڲ��i"���p5�����ɲג^6�W���U�c'��:Smn}� �ݕ)u�S�e_�s;����� ɺqw��h�t����+����w��q�X�Rf
���J��<]W�@�MKy�Ť�'�]zeVY�tт[F����~�(B?�g�jʪc���i�ɗC���_�p�+�bIP��j��gD�G����>*���vp���F$	���D��-7>�,���I���]Q�d�[��,�=u�6�M_aX�fRw�T>����GE�;�w�kH���U|$�E�`6|��M�r�ܛ��H�
LP��06���wH+��5B:U{8�Ħ�~![�F�	�M+A4[<�9���ڂ�� ���S�Ь���?K_{d�k�f���I���m1�I�I *��M�0��������x]�;�}ջl},�ߢJy�6��C��i��g�Q�ΘJm6r���x�~Z겍������D�+R��`��)���x�|u��_vʏܳ!$�"�����.���iϦ�|���t#��\pLS��.$f4H�w�ɀ����4��L�'��9��@�H�~��4�4�D��o'P2���ǧ�B�����8I)�[�c��K�����c�$`���^���3@HZ:+YD�����0&D����v����kez�����$�<��׍"'��7����`�Bk��$1�џ	�"h��`q��|/V&Rc�g3��DMI�ib��*�ӷ6,�a�,�	Y��Z�}��k��z���aǪ������]�4?����Q��H;N,�4��2�K��㉧�U$E1$�o��e���T���L��l�7X{��$U3�|
V��4�ؤ����\e�43!80�G�s����E[��������N�{CnWdګ�����ı�� o�b	TM�:�[֩���qT��<�G�t~e�hR�9�����&F^Ud���R	��;�R?��e�{������Ӽ; �-we�Ћ���8�6Ek��������Cg�fT+2���ߛ�����Tk�n��.sy���'Q��ǳ� 9{c��Ƈޏ�\� �Z�#ko�wz���wE���A�/���es��vL����h;\8Cc$�6�~Bs��+�L�u��V$MF��F�䂊�/�(f����W����[��ɐ��г/m7�]�g&h��6�;����#J��\��L��' X����"��O>�(��b���t+{�����N�{���g���X���dt�����*<�ͬQ����v���������caA�#_���:+޼�;�v�녷?��uW>9?��p�6lY�ԫx�����^�s6\���E��ibŁ)���4?QGj�����}|��|����Qo������?�=��\±��AZ*~IX5$۽#��j������f� �<ǣ�<�!t}m�S�Rd��b�������b꟮���ս
&O�֦w���A�TՇ����L2�ͱl��8���Fb�
/�N��e��%�v��_lT;��������F����h�@��1�Fa ��ffӚ+�g� �Y�)�A_��a��s�]SP��[�Y)p���7�@��E�e�5W�	��ҏQ	Q�����k�g澔{^��h�[r�6��Ju���n�EO��Q���x�Pi��S��6�Ă#7\_���G)kzg#�\�&�K� �0������T��Z�2��!�%���h4�Ӱ�1U=�<��+�����-oq=z/��A���ſ�{Pa%Kb	���:E�eb�S�!�cM���L��v���H(Ȉ���x��+�X��)#i���m��h03ݒ�=�%f�@S�i����X��Ζ6��#���9aJ,:"xE2���/���Bs;2��Ä����j&az�� Y_�WO�����z��k?j�Fc�}]��S]=]�>��1�x6���3�+���k�ۧ�J�(9W������E���>g������~�C��z4�'�j�4�����h�JK裖��>�����婘MT�	�.�����td
JC����<P���R�G�>d�Z�^����]��Y�9t)]���vz���o/�,r�ȚK�@/cD #ÔW����u'�5�^��ɏ��k���S�����;چn�	(�8��9?7؋�q
�
ZtueM����d,8�]���&��E"(����.��k��E�B�|����:�n(���+�RY�l4�AIAw��m��	��+D���s�S|`�5��W�H���a�o��Fo>�A	����D���vua�w�Ai�
r!�⥵ɉ�Y�Ĕȳ|����4�q�X��tb�p��>�K�zԷ6�֜e����)�0bؚ�fa��=_�C<Q�X�R��_����W#l@��AMj�3�����̀TP�u��ҵ�j��\�XRXx�������c�w��߁ˑ��q���;̫�Q�c��޴�a���ԋ�0��O���[�NP�00�rDQx��М_�{����}�;�p���aq�>MUs��e���/���g&ߒ�d>+���.@;m38��F�N�6c��!!mY�7�7��`�?������J�dha�?�.ڞ�C��ӗ���];N�3���δ�7֞����B�S���[�=8��#0�H�]��%��2f�A+�H�F6:�6���W�Xq)�{_�>Q���=-0�(�qS6�����F��z����v�#G9B��X��g�7�ڼ��!p�M˪zK�I�{9���xB�f��(n ��[iǲ� ޑ`�b ��"�g�w���i~�Q�ZI�[Y���qtflD.F�VK��ظ4�U�8B(qkAo�2d��@���v���>��	"8��c��p�D���K�c�Mߓ��J[���f����̊�J�g�o5�X:��+ ܰ���(�̜J1�S.�c)Qʜ!�!���Ā���M�.?�0C�-K`��y�u�wɽ�׆�t������@������-�R;	p<3�n�d!���{�R�S]RJ`J�m-7v#֮�	�n�Dz���@���v0y����k�F�Z!&՞d��	�ձĲ�����^��;��&q^U�D|��B�nl
Kt�V�	�"��pH����e@`���N��h��0�H�����`�`�{����eq�B��� �B>������n�v�[�y
v�;迍-���TXA����F�=���U�o\�jڬ9�V�e���k�2ۑh�R%��Y`Ԗċh�s;�y*��Y@�ǛfL�y�(p<٬� ȴi[k(+�������**��{TL%&��qL��{�@�y3��l�y+13��Fu�͆�}�0SH��(�)��T��]K;����������>���%ڢ��ؗ ��)�0�9��ۛ�ƅ����X��e��Fj��6����zv�}��j�g���i a��:b��S,?L�^Y��ca'�#�*9,�C��hW�f�d�6~�� !�vS�X[	ĄlK^�u��x�'����T�,��5�1+sJ�,_!�l��NB���o�kb,$�秮�A`s�Y�+ѶH��D�&�5�D@F�r�^��y��痢�Z��k��.��w���JFB[U�5�l���&`.��ÕU+�H�E�:�� ����R��j�rw�6��C�7��6J��Z3࿦��q���N ��1u��~"���F�A��uM�!���.cN�:��H�7$�]�!���Y�7��Ѧ�Y����!�zH<U�ٲ m��Gq?f��#"?\�����)�P(�](����&p�Dl}ƶp(�5T[l�C��V:a\�;�\��X��a8�B*�)Ua-��0�A)��ekLh��UY�����d��h�ꦜY�C���L�$���*���!��8yXn�U���)_��~C�z�B*�6�Wy>�;E�pw�7>�����(��1��74�f��ap���(l%�Y����jD=������5��l�v"v��r��Ȇ\o؃�k���o���;M�$�<8�0�Q�<�~S��3�an#z�_}!"Vj��.�l�r����J��G4�+�q]"L�_\����yp;�T!�m#;Ω͙f�u�u��^�PaV��&6N�Þ���ҥ��6����1��3 �*C5_ZY?FZ�� �M��t`/z��o鷲�[�L"�F��C���m�!��
��r�� �`M�PY3�[�z(K��S ��hV��yY9&�٥��da�EO>��l��6y
Tŧ�3���n�3x�ꗍ6?�����������5���i#s˻%���/��;�^�H~����Af�a��w�����bܪ���ĉY���V�;qs}(<��\0��6�)�'�P���gs�=z�X �:;�B8]�u�5����9�Bn����Թ���ŷ�w��fu7����z�j8�v�Ŏ�9T��sVi3St��X���� 6�K��@&&���+`FLo1�ܿa�nB��*�\�p��p���ǩ�u/_�-�4,7�s�.�ڮdY':َS������Sh#�������.��|�|��cu�=;��7|�z��r*V�ө���9C�LU!�;�"�E#U���G�`�FCA�����d7̚��+� �H�V�����i���d8�N��U��� a�}�D�qy*�Q�v�m#� #ͅI�N��V���#��P҇p�S�ޭ�n�ӾZ����aQ�A�,�tT���� p�3�}�QtJZ<(j縆1�<�е;;+�h��������!n�7r�pZD4�!��]���W����P������?�ȧQ+�Be�R7���E;���,�k.���V{�_�=k�
�j�v1���\�[}<��=&��d�8�d(a�/�u:55��b��^�ƌ,�1,\5
�/�`>f)������p�^�W���@���s9	����c\!�@�!-[h�}����a���O�m� 07��>�t
yBnŞj�$v��B]8
�cH`',�:Fe�{8e}�鞥��q'1%>yo9iA��}��@�_�1|_Y5Y���H����*ON���E�;��,<�?p��\��QN?��3�l�����?���ޒM�������;!�wy�Wz\�4"e(��>)��gi�������9+^V�"2ҕ_L�F�`�*<C���?��m�{���6�+��V�1,�31x#�gf�q	�{QK�R��������3{��h�0O��E�����A�1`�n����I�$W�������J�	��ݼ���-�s�j{����G�� �4��+>�&��L�rl����B	��uh��U+����
2���˸d�6���x���g��t�׿?�9����`�UH�� xc6	��o������.0m.�������7�<~�w�:��q�Z4i��a�!x�}�֥N��<�"�1{�!�)��ĝ�S�A��"ڼ̥���O��;/�f�W��8����X�SA!Gȇ}9l�H�̹ �U6Ѕ(E=��Gލ~xԴ��^
=�Y���mbB$|J'ࣾ��h$g���^�Ts�-H��}l�A�v�Uܹ#��}R�@%Df��t.�,tU`o�Nh�_�kJ.y�ܺ���km(�K�+�Wb��s�'���N\r�����9�K�����9_��q��\�8�!�u9���������n�b�n�����Vaa|��i�}v�D�D|?��!�9��i̿*�eW���w�$������=�7"`G�o�D
,^F	����2�i�e��3���?���O��>^�q�k���$1NWH�TJ� ��XjV��;��9�%/V�/���l�,��kU�P��(].�jbD�fԙg���J�+:}��������'��e�n}�@9�T��s0�m�����bl�&r�GkG�}�u�c頺jF���ˆR�a����n�D�3.R����<�R����<O���9o�V�.��4 �Z���fP�����Z)���S꧹�N�L�n�ê�{
��<�H��g1P=��|�m�:p*�����'�&���P/�MЩ�-��<nͶ,N����1���GJ2t�i.Z���_i��=@_>��O#�"�&��^���j�c�N����G ���a��y^EJ���!�;� wW�b��bWTc4�b��V���e~�Z��}S�'?�>����nSSY�h�m�"�����r��q������R���6����l����~�uk�wH?�&�OY�M���s+�CI:p���7�_P�<�"j���/�M�di�,�� ���U�rġd�]t��0&C�1��}���CP
p���1aw�Y��PDV�W3�DI��)?�,c7#-
FZ�t��4�A��S�A��+��r�/wj���¡9Ի�t`�{G�6̰Hk*��Ť~t��D�����Kh&�<Oc �K��%s��9��u��Ɨ�N���c����W��s'��9T�d�z�4\����Ў2e��Ĭ�XN��ҁ��� S.sI�Z���^�ϖs%�V�X�>�Q⽕�t�:��G��d��ܿď�S���2�3�o"/&o���#�BJ���7���w��|=��0��sy�
:�+�^�Q����t6U�4�*������8�>�>�5�Y=7�x���瓆�D)^Xjl�.��L�/����A�s�N��׍��ia�`?����P�,��N8�m�LLuQ��;��˚���4������� ?�_�&U�e=ٛ��dxZ<���o�O�|�~'#{�b?��#Wj1\��5��F.�S	�7�����$��� 1��K��~9J9�ȃn$��������S���
���笇�Z�]!U�Ѹ��y�����d{�3�>��'�\��T��T��D��\U:�g��N��^w��:PN��O��!%�P_���4����@@�G&�o�(�5=r�Y뭜@���Aw
^�H�T,��u}�6��̭P�k�C���W�}(�3�c+�7s`81�̒�J_�8�~�iv��/� ��9�E��)� �v*Ť<:���9+�)��$�?���@��(|l$�3����~/�o�mF.5���b����΃��H�+�9X@i�߭_k�|ay�:�w����_��x0��.Rj�{�K��q[(�w��_ti�)"�?�����(�v)qv{��w1�}̂2aP~&��-��.@��� ��Z,�_>��G4obç�@vRs�\�S1
�EW]��>8)�ء}Ш��K����!Im��ث1qɌjnߪ�#��XT�`�bp�W�K����pC~ ��xy`���V���t�_��Ѐ��O'���a��~������oIV��-c��m��~�bũ�	;�Iƍ�265O��U��(!l����_� ���m��Y��m�x�rc�p6��y�j H��;j����V��Z��Yp��^���}���L3d$@1l�)������~�P_�<L���r	"���t��T��]���e��5���ߞ�����������07ʉ��d9�6��P�	r3)k�A"�X9�]�"��B����W���l�:�]���4�|�ٕ	4��Cu1I4F� W���aT�0G�/�s�B��ci���V�����K���?��L���9�'�v_��>���)<�٬i;3q�mʊ;x��?r*�5��R�ֺ�1n�
��c�a��5���Gnwƍ:h_�\��$�?h�pfr>�Wś�T����eBGS�Y�fL-Amr�8��ZV��=�P�4�V�`Z�X��\�_��s
�J�<V�J�21�I�|��Ωe[V֓l��2�}x¹^5�]cq5�-�,c�K�.�+S�=����#���ר�p���*�(O+�wpp�~�7�Ɩ����S����w��)_�M�&k�8`��/J�K�F�rM6?֠?�9gP�����h�&��y�څԑ��@��t�8A��s�k���;���9R����P,����n����R�k9s�7ny��#W�{.�q��Y4��a0ЊA����-��hGWf��i��������:Yn����Y�3b�"�>;���lg�y:����j��]�b�ɿ)�El��T�U�2_s�o������hc��)���4��=�U��M����m\�m�}�܆�HߠdWKS,
L!r&���|pk0��q���B�����e$͏ʖ�6o�2II@ ВC������&�&�+~�Z�p��z��e��g��cu�_���V��l�^������qgup�J@�'`�iL��!<5C�V�W+F(�Cu�;x@�T~��9����)�YCY6j���*<���c��!OL�J��sO�PX��D4S���W�Q��:�`=�����9K���v|N���K0o/���WX׃A��wUz��B`W��Zk�V�Mn�ǎH�S�����kIќ�8%!0]H���8�=�r�Ie�bv\n����O��g��<��l'����+��Tob��ZD�Zǘ�@�B�_m���x�);El�'��,��.zC ��ƴ�@?t��~�t���E��N���rͦd�K�>é]��.¥����T�p7�13S����*6�&1��*Q<�A��>#�)��x�$���a'��e���}d�����ֹSO�閽y�oN�sy6���G��&u y�-��� s%"fN� ���e��D���NL_�����!��cl�È�%�Q$[�B��Oo�io����mf2B�%�kqC^CH�r:�6��3(F��`��n��#B���{&�숀n�
�ŝ+����.�G"g������aY����E+���Y�)�.\������N�P���^��frzϊ��ȑ� Ír��5H|�j������:�p���df������?�8c^�%S��sF���Hf�	};99�����W���ٜB��yH��v�aV8/�G�*,#9dO|�jqJx2���jíq�^5~�k��1��?��J�^��P���3��m�u`�n6��#0��}2OE���_��(��reB�ye�8߆���{b|�nuN�t!%��lm��p������NB���0�禦��L��xv��>.�	H?&�?X��w3c�"���
�q�9g%������
��F�"���C���'��_�c6�^��,��`�e'�K	�Mi��׆�\]G�d�a='� �	ٞ&�9yptgQ�
]�˯��-�ڏM�����E�����
0�Ҁ�0�Y�G�ia0���Gr�^�4NdH��ƴ@#����:m�3�\b���j��;����!����������N����d��E{g��6�J�g= ��[Y��S��մ!��xph��e�=^�jH�d����x>5��=3ipP��0������
IeXENЭ��	�v'i;V���F�s�ޓ�Yv��G:�;���0W��rtlG/ǬI�a���A�Rbd��S2��m*z`De�����^�*^|m���19�5�7ƺN ���N� ��#��V//x�Z���֯�(iN���lqq�k���L�l��S�a�:��0R?K)�ni��3C�ƛ�#P#���P�v��rY��>"s��e�`���@����Ip^#��X$T���n,av��/
� ��k�� xe@���ۛ��.����i��]!	�aY~N������NU����W堺�rn��`B �l�I>��%J�+�n�\6���Т�Q)�K��pA�0e�t֨PKv��_�*��M��ll��m�E>��罘��l��ɧb�@[�,�Rl��s�9�v����3"��B����tӧ`?���8�y��dI��ڒ��$٢p�	n��YI�$M`V�C�1��~�?��i�R&�
O'V���go,͑9����i@�+K�Y����Jo?mYbO�%nزl��)�
���むH��U.�5�ጔ���g��p�0���3��p�,�ɛ����z[%?��+�[�����Q���"ޚ���Q��^��(���n�*p�<
K0�fn��W�N��Ԕ���&��+��\�_
4�� ̄:��~V1Ξ|j׽e�b%,5i�� )���{�Q��X��-%N�U�Ȁ��w�������	�`S�q��il�����=��4X�*�� a�%�fZ�NF�rQ�h���.u��W�̟���^R�x��,����������SP�֦-Ļ�*��>W[��K�X�Y�m�)1H�k�^C=[={�F1+5�v��mh*�Fy	�����~���0#�ל�k�-}t^Z~��1�r#��x�v�ho�߬�' �c�;ͽt� ��j�̾6}^-#4�z����;�T����ښc��8{d�}���q�5��
�߳`�b�I"��t
�]��?�9qe��\A�[n�56j�m;O �Dٮy���f�	]J^$��hb.�O,A�E\Ԏ��mb/�ڕ�7y������[�xݭ���,�s
���`�����r�kҘ�}��/�*��x�*�J/��z�7��c�B��tՄ;���M�"jc /��T��D��I��iN�>W���<y�`m�u�+��a�S
�$?�r�~����N���(�$ш6GZ~I4bN	�s�
�{��}��ޜ�/*���:.�\B����v{���#�3��n6a�׿�qG:8�>O�a}�D,�jERo��G\Cr�xWM
I��pq�^d�M�loQ����IP�4"��i9y�Ϭ�?4?o��:s�Л�ɲ+���k1"��qYW��W�ة�C>����YճfRi�D�v\��n����h�-�E �2�`�_�͟���ݏ�ɲ2��G4��X�JdE7�/�(%�#�O�����T�J���{�f�8�Ֆ\�6I�(G��i4qt�N��_�͘��W9���Fǥ�p���%�G��>�Ҥ�xe!�J�I��@�b��g`�<R�8
D�q�L��r�m��@ukxjR]�Br�	J��G9_��km9ٲ/>s>�~\����-F(Q�����?t!`���G����c�wM9�����_�d.�`���0Z�<���4���
h�^p�ѫQzՓ�� ������lo��5��*8w�(�P{Y��f�V�[���S���K ,�a�Az����*�Q�v���7`�#�H$Ƀ������;�F
&ae�J^��z����|�>�p��F1�Ҝ�h�!�Ln�9��Y���H�!aޘ\F�����p�&z���! r>��@w��r�ު��b��4|��k�Gi�zN��ٺ�~^��*�72W���|�-b� ������A���J���e�
�A�i�#���|谠G�0
.ZV(n�B+Z%{=�"6�k�*y
�!���v'���i[���P���IS����7�5I��6�Jܾ�(�)���W��x�ʯm�M(y�r�:�������Wz�[Ǉ����_�jI�ܥ�����j ��������a_��R?�8)��EF��������kW[_�Q��YE�y�4��ڽ/��-�������<_���yQ1����ef��K���}��>��a��s^�;	IG-y�@2MDv�!�r��#U��~a�m7`?�t/GFq������1����1�2kF��Hf�z"R2�F�+-1I<�ȕ�|�EF�;��郞��=ϥ\�O��	��Q�Y��a`.�K�=��ܫw�%2�͌a��#1��G�2�����8F�'p.����Z��L�w�-�W<#�?���blf���YQe�Z�i��!�B�����##��T�Q�9�z�l��+wf�q�r�w�G�VE^��U6�_R��L<����$��(����g���@
O�vfg**���N�L�!.�o3m��us`s1v���qs)l�Rl�*;K���]�:�ۜe�۵���7k��_۩7ӝb�j�M�2�rV�.G��8'o~�����K�r!� �\?\+����S"X^����?���%����s���5n��Ȑ�l�x���W��8��'��(�����\K��T��X�x�ź�m�N�.��%�OS�F�6���������9�� Y��߲5#~_�����)������`�Ԣ�}亂#����+Xʊ0�g~�|55�7�J�O[p�#%$ږ #��{�2ÈӸ��;���M����mǼ���1Tj2��:c�ЉA,�<�X{*�%���9��R:���|�̡k���o�Xd�n����ԍ�+&LS�����x�B���ib?N���"��5@u��-)�;/�a�lu�����N%M��t����˻�:����DM��(�����G�6Eb��u��C��o��k�nN?��S�@�4L��v52�G�v*�cP�n;�ŉ�Z���_A�C�"���R�������(fc�.H�v�;�Ԉ��/�GţV,�]>q���#��vб���7�����N@�VO�+�%��Z�R=>yM���G��5��3�/N����#��a��o|$�}J�%$�U-��K��9
��4���e���yg��bk��n���w���z�Ta.���݅�&�/S1�[��-�p|a@GQ�+ҠxבN�l���(�zd %Ł��`8�Rb�v# ��}�Ա����[ d�O��M��^z�䉌q<�¹�����l	-��R9����lC�VY�B��P0�Q�	�W�2y�����>�sO�\�7��5��z~�K��'�4�z��J�0���X�H1x���F�1)��LS���а���[���V��u�(�Q$.����V����#�9�J�2�-�D����s謒TRR�hPl@�`?s >��j���~1�4�:/l����|�Д4s���`PԻ5���#a��ȟ:e��욨h����� ��p"��n;�ڧ��[�/�XO�֧��λ<}>�W/�ٮʟy���؏;��Î�³�x-7[�j<�C;��'�8�"����خ�	QDz�����(��W�iO����ӱ�F[[�VӤ��=`���0r��B����q��ZTX+WB�4���iH֝ᝊ�9�B0ƑpX0*����%��*8CH��4i� �u�/xv�S�_��{x���5�r"�4��5�[�äۑ��(8�a�̷x���w_W�[>E��ϫ�/�a�
E)f?�Kr2�\�oLX��J���n%���.)��GX�;i���uػ�\6L��p�������_i\�gPt��!,�L��(Ec�R\NCS-�}L�Z�aWȩ�a�z�n�'���,?QK��ꏊ)����S4�qX�ԧf�I�@�φ�B��{ @~l��xk�(n����X�0��_�z�+Aճs[IER�"��r$���H-��͋,#IF�\�?�~�� }W	�(Q<�Rr?�$c�o�c9��^r�H�Z�z����a�3�q뗐�~�c�d�)��/��t\��������1�d�:�x�F��[{��˨�%W��Zo{�d�ICވ&�	���=p�-�:��uL����u��_B����|�}��6l�C�/c	����fAO�ˉ;6o*m;R/�� ��\T$�UY���s�նZ��a*���l)��"P���yWA�e�,���0�lWʒJ�-��a"(��3�n�e z�R��"t���x�`B?.)�#	��>)�I.R6b�xG�WjȠ������y��F���Ӏ�P���Y�?�q���Tk�$^XMt��D瀝wW�|����GG���	0~Xc_�����A�>�ޞk��}�/���%�/���jA�8�d���{^�Ԕ��h��:�¼��ȼLI����ᬻ�:��_>+Q�Q0�@�������R~�N�: %
WH��<^������E9ӝ@�E�/1�\㿌��cf!�=�M5��g��Bn��82��ʎ=�]#?
��1�SL~pd���ƍ[�f`��Jgb��b{1��ƶ�@诱nN���v��X,�Őy
��-�����厚�o��Z�i�i18��L��IS��B�5�A$�W�~{����[�����K�gh�pF,�ρ!��"E;���:Qپ��I�2v���WrG�A�D�T���B��S