��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~Q������&}��5�稸�sy�1a�n�����Vf
�^�!BLB�?6�1K�@8e��^՜���\�$��[�v9�M18��������ܖ�r?#�r��j�-m,q�:�*�'&�U(>�����͓}�1O�G����6�d4�Ux�X<�lnb[!��.����v��{n���XX!���UW9DGZ�����w	v�'xf|+]�VS�tt���kpa�B��F��Gt?�ep�#1�;���ſ���:$�����h�mYt(+Օ�����m�pT�=�@u#y��Pv�	N�.�鋸���3�>�7����k<��]_�QY�Kr�^�Mn���k�����*�ɥu�]� �^�j�Ed��ZOAyB��jq��4#�G`G��u��j�I�{|(���:�Xx
��Ma�Ѵ�~;�� ��Y�~;f4�����S}��*�^5��8��+�v�qi��%����-y��&0��ن�O�)G��ɎMqF&�o{����.�>�^6�,+m���!;&�Z�(�Au���,.P��C�h��C�b��,&o����o¤�}ܗi�#"�0��f�4���l�� ����sh��+��Mu�
�o�8͉o9w,{Bi@�H#�FE���7����"�iSo��ֺ�.�rB|�"�ޅ��sk��R�B/ =��T_��P\�[y�:�T����3BΓ� ��?MV�`j���@��P��x!����1��4t,��ڲ�B��j�=0���� �31�i�}Q%?&K��x�n*&xAE�@�<�l�#��q ��DC�c��+��������2���<�?N�6�?z��ˎS�|�^�f�kR�d�IJH�-�:]��%��f�ƶ9��6��}q&��Gd<�QF��be�3.?���OE|�vI1}����	Kj��e#���H����$��B�#�7]�#R�}?�X�����}Uyk����ZC	�F��(K�**W�*ܖ�����B�hq7H��ց�Y� ��Ǎ�����N�7��vK�ŝ��f�,� ��k`���t+&m�������|A�r��U	n}�˭��2G��v҉inW���~��2�W�3�y��vrׅ7t��?(U�Օ���`��Đ��d0sS\��������o��QAX����}��6"eO��~ᗉ�1�zR���#?��}�l��d���OQ.3�o���p2P8� �DFͷ��P�'�uSQ�˴)���9�I-����X�4�v~��1�L;�GG+x�{��RP��E� y��q���=��[~�?2�/�CF�ոSǔ�Y ����x!�/[[��LFu�"���ie�����x'��cF�k��M��c'�?�R�5�S�a��A���@�R㡌��lVlx�or� n�M3�b͔��L[�,���bͯ��m_�F��:�>=B\&�tCR�a��� ���B�x�)��z��B'�A�%�� ��k���&H^��=�͡`�������BV1�ȏn<�@0����v��7<餒��O־��,�ob�;dCS�Q}x�Y�Wv}�����8��L�$��/�e%</��ҝk�l7�sV6��F"��KE�̢��!�c_8��ɩQ�=@�`E����*9>��G�z�DS�äf����}�΍����X
�ɮ��1��aNHS9�9�{�h��X��y��wPC!��1I
���i)��u%��_Z"�l�?�6j�E�[���m�ϙ�nO������1�ݬ��gHc�wB���\�������Hc�>}H����u�YO_K�,d��[��	~�6�2�*�dq�jQ|�������2CݭK�+��/���NF����Z</(���Ξ���nS�|P��@/���FQ-�RS���X&��=��{��,�|����$����� �FOh��q� ���#�O�-�M6��f�d&ɲd���������'Z�g]H6���D�im*��5$���C��M�a�}����K�%��M�F���t�pfw�z��DD4Ґ�N���>4����Q����q!��z�TX��g�ZO^Ο��?`�"��.k��vx��'PӎĊ�9</�K����`H�AkP��&�BE0�����v_�P(���ѽP�\��Re��n���_�Ik�f�]�u��_��6�\��̿h�5���3HBC�o^�����?ĳW@k�~���zs��= yq�_񽏐OK� %���	�g�aE�=����f@Y=Y��Ӗn�<��YI����L"��G�ǻ�o�	�j��a�0�q����z�H4�:�5�zҀ�dJ��=��"��{I7�+Qh����
���1R�7�
�����a�h�>���U�P��1�I&rvb����u����Wp�&�"ݔz)�����k2K�����Ȟn��P����]�H/l"�=�+o�O|W{������o_��7b3�:�)�ɍN�h��3j�fY��˼\O�T_���N&�$����`�"�굡4W�6�s5�b� �L��ݞyH :�FX�b���\�ɜ�i�8`�@ٮx�YE������ww\��dzJ��� �<{\�blD�����	�~&z`�s�0�H���_�����ڮ�����~������q����G"���K��	�ѐe�8�_:j�7��

��~�D@Q����ڕޅ�'�ΒĜê��^�a���"|(�}@ J��Q���PAx�%�0ʦ�XE�����W\�{�M�n�������2��5e��)D??5wia*+*?S�!���<�M\��r�>�1���|�k%Vh��h'�Qa
�5E�wObw���22�$G�K���>��fꎲ��@Gl�ǫ�􀎳���0l6��ܟ�f�jT�*�u���y�e��3��`��똝���U��k�HQ�nJhLnT��VCܲr�غO���b/����S`X�]���NO��pUsg�Ǌ�]'ę&Y	EӼx�|L�k�8�Y��O^G�;l�'_��0��$Y��X5�߁�ƒ�T�JB��x�k� Ԥ!%C^����E 1L�|�ɴU��3נ�/�Fx��c�A���w�"��e���Ak��̝AA��Jt�6N8�����K�>>z5��\?��dy],y�?燫��2`*��{5�3<��j\� QPLW�u_����3��]�fK4�R;����1�ĉ}$<��$ I��
:�U���?��O��z~n��$�K ?�&���q��ǘ�� �U�ϣ�Ϗ��I2����'FGM��qC��:���2�k��K��e���\I4�6���f'֑�;V*9%�̄@s�5-�w��?sh�z�d��B@XaC��N�ȁ��b��$�Ώ |�i�
\A�j�ۓ6 �vX���p_47����|�ߥ�a�<*�ZӮ��n"c�7��9xd8��� �>U��&��7R򋾢`��dO�fw���?�ꬣtS-��x������E���k�!��d� /!�������{��¶9��2�pri�,��8L>+�"y96\/{���=Y��eL��q4���Jt�&V�%�wHcљ��&�D�f����� ��}%�;�f&�'�"$]���VY�p�y,��>s>�kr�\����p��ǆ�(�*wo�[)�9|)�L#�"����~��Tw���24D�v�Q���.��c�~fӯ���󾬵Bq�J���OV�)�(��/�� �a(����!��h��i����I����U�}�)d�n�$I��c�s�J�,�hlɰ�;����8�z�����D(K��u�3)x�E�P���K�wx�[����s������?Azqj:PE4<�$x���q�}����I�H*˴��LVu����S�?��+�+K�䟥��ӕ���+�� ��QVP�"�妜�x;$�T.�Z���U��A7�CU��%������U� �Z�9V�-�<��0Q���>\~�.��kR�
(��55~t�j\�w
k���*����V��>G1�ƍ�P|X�{Pc��O���
>���H/��u�w���'e���;����Re�P���Z2�ʸ��l�IsJ.���.%E"k����wW�d���-�el�ɟ�P����-Q����D�AL��
�﫜6�8y��xA�dɆ(`�^��ZN�P���Ī�E�[\E�Hm�[��(����3��e1(�%d���/U�.����.��5��r���o�\���t��k
~a�b�G��<Ε�(�v�J�\Є�X�r"l���^����0��Z&o.d�JV4���O���fJ����ΪU����E� k���`*��!�3FҖ6qD�ݘ�S	o���d���Dh���J��Ϩ�O%Q��ӵap���#�d���ĕ���;���#EkU=0�=h��\�/6��H������x	D�Ќ�,h�;H�WY�D���lc� ���R�X�5$�K�lC���t`Y7���g9 �+�ߦU�-�լS�7�S\�" ��W/��Io���?
���{U3�� Bt~Vfr�D����<�Vd{����00���z�ѓlK�f��71S�'1=�YP�.�H���:��+FSk��f�J�L�j���}��R!q�Ά��8��>Q�9/�߿��F���`����#���`�1=�.%-u��]�������z1��x�b_�X�c��Jc�'�@�f؇+ٻX9}�KL��Swc�nV(4ӓs��j���I��ͦQ�J����*�켷M�e���	��\��s��£�C�!0��z���ն����|�����,�;R����)�0��l�&EW�����?�tGs\W�g�v9HQX~q��0�ݓSr��qQ)� D(ʹ���f���uf���l�!��Wz��q,�G��m��(�1��~�� ���`Xq1��/�)V����\�8p&�ѹ˯ f�w��ϋri�n��ě��uN�d�3L���~�:Jq�2�=#wq n]fj���L'��g(s�R��ɝ��"2͜Ļٴ��/!���94"�Q)�@�"bY�}
�R�B�U�W{�~#�AF�l2I?F����r��ڋ�{�:��!��z�I�I�����xH��XXc0��M���x�p�xZ ��*�� �e���N��������\����+N�M�C�����'/W͚d�a0UזL<��yj�;n\�;��cD�`M@D��n-Ԉwa,Y��r�,?���	� S�+�����`[�ިF��L��"(��T�&����4� ��+,F��\���0~#D���%��󪶃M��h�ӛ�#��us"T��ۇ�Rm��1B�ag��V���#�Z1��=^��Pd~r�X<��#`O�m�p�c�Xb6 �m�j�a�2𡝩X9&�Q�F�j��{	�m��6>'��>N,��.鱡E�J.$c%j,��&�u��8��@yr�}xv�澂�xJ-P��{��z���ӡ����|��Wo7b��bd=fC	�ϙ�P�⦶�oʍ��%`=s��S�K�1�R��5^�����#G��)��D�2�ix���E��$�f����0d҆t$�����������8��ʌբ�;|�Ƌ�u�oqf�P�8�T䪏�H�G����� �K����T�������*�f��=�3�o�P�K�D�{���f}*eW��.TR��>X�
�q"�S6�TJ͒V�,�h���j�l������>	��� w#�Ci�7z���N��>^�ld�Tf.J%Ż��Ԇ�L(,RN�>m�$����j�g�B��l:�0b�����oҩ��=��A]ۄ�\�$�+��ʡ(����8!c��Ϗ��O�'J����達�U����tdI3	�(�+������L6MX�kt�6�#�
�fi�KԿ3M��Pu��D�?���K�J%"q���m�Ԛd/d/���!HY"�}�x2Y�w+:ނ<��C� ��vV{�Nܿ*?j�<��#h7�H�$���Gf$���5�>�X��o���*	 �1��yk:3��ƙ�_﯒��>��Y�r"��޵�(�A�9(��C7�H������BT�fj���S�$mG�6/��M�*�eu�a����a8� ̑v�ݷ���2Fx�h�iñiUx��
���ik4�����MWN+34YG��SS9?QJ�����CܟcL�:�!�$*�Ƅ�Lo��Τ<����a&�X����q�yVc�4q��"x|����԰A�:�[2O��o��?;{^�$Z@�=�>(m�|�`�O�R��ZN缣4�{u�7���p��ov� T1��b��	3ØSyբ�o��h�UH�˻��<Ox�K�(�u�)>� lxXu�h3\`ez��ן���!7傹h\���^a�|�4���s��{ˍ�OE������2 Uc$�cT�����8�G"ŕW2(h!Gg���A-��a�flKwr��Nk�8�{�t�����]R��Xd�PQ-���?#�ܢb�O��B�$�����A��|�]��h���O��=���9�q]����`��V3��K���_�wU+�x������/�DQ$��x����5���������av3�� ߼^��s���@*�7��(�4ݕ���]�Z����t�.)�
x�5��9# &�R*L�����n�Sо�>JWu^��ѰHN�RGt?g�5g������KP�ۿ7˘��B%ZXV����V%��F�.�;�nS�k(D����R�D�nQ�1�3����P�D" ��$��������|���N>W�E���D�Q�WC���n��b�5�t����m1��g%�5ߩ̇ZA}O$9vk�Ψ3���<�v8	�O���qÞ��orٚұ��	�~u���m����.x��=R�G(1U����c�-n����H#U�v�rh &��T=�ȳ� ��r�,y!FEׂ�%�s攻$ɎW0�<�J�-9�$�xץQ�v��e��zM�̩Fا�#U��s�𡓢ɘ�s�͐d�h ���*�-P,�/�x2(�"v�w�f�S�ϊBc��!�]��3���ǽ�G����QJi=l�?�d���'�"�����6Y��M�!߳�1e���q�$2V�J�1-c��YhGb�b�e'C���g��y��˱���)x���d�~Q���U��".,̠"��Z1�L�Y0��|$[!>i�L��!XX�i��==��l]_]�D3�l�-���V����9�b���1��~��wG�Kk꽰�l��-��� �@rg��Y�\%m��;G=��`(T�r�r�{~��@Ha�Hw�E�^>�b������]� �;�cb���;�WT=���j�W{���WV�����S
*U���D�����o�O�)&��A�B�j�u���9�͍�>��_.T�Fwş~�d &�=�0�xh� $q�`�G�)����O��łV������f0�Ss��F619ȡ���)P���)�{Yxt۴9N��[�դ��7r���7Bŝ�PRN�G�h��C�QC��~o´W
	
�i�
Ӱ�g��TAf�Ld�-�o�ޭ��,[�)ե;���1�k�_�|���as���R�8#��;���h���s�|��9�N�?���}��cث��]��Q�$x]7c/����:I'�38H���o�[iވ��#�G �q<[���r(b_$ʜ��O�m_�?�]
/ �.In�Ry���j�!)����Y(�+�u*��n_a��|4+���?�c)5������x.�Hu�J|��PX���]�G�����'�&�N����|}����W��K��e�=���24����{�5�K���.t�@��8�#��L��D���7�Kz9�ᗥ�,��u损E�M��y��ؗ� ��G�8�����s?#�SO����'�֊߂����x�=HʕЂ����p�!¥/X�?�>�x��Lī�O0䪘2a�_��Z�?
���/���a�g/|��99'�;�$Mu����2;��Y��p8][$��E�-LMw��c
�y �	;"	�#r���x�whrr�5�'�������Z#0�yf��sݠ<Όg�-i\�jN1�ƈ>�@!H�Z���9S�Y�O07��W��k	�wtW�3Z,km~��؏�$�ɺ�U�MM�;�Gd` ��ׁ.��jA��SM4/�?�'(.V��YA��<�><�h���k�ؼ���HC,2�s�1f�[��# q��7�'���D+��[���Y:طh��4���21�-̞������`7sɲ�H-≁���;"�������I&w/�?�y��˽c��E�%+���a4�lK�^^�v��_G|ߡ*���OX���`q����2�~��`&
ّ�����n�]������9�1]t�خ��v�1��u"��}��z/%ǅ��QX������0��r�J�;��C�����f��wڙ����	��-�:���ok� �Mrjz���M��D��?������>%e6B����#v��Q(ri�p^����1������%�n�e7��e5�_�����'4��X��n�+�H�KX�mqc]�_��[��(�'��.�k�LDⓁ�������C[{�}�wJ%��@Z̝b��N��x�/Vhu���/&xe4���{~g%�fҖ��������\��C=��q�R�?�O�Ȣ�0�~#*8h ���QD����~�uf}��,fS=��^����Oܖ<�\�T}<����}����
�P��,\����xc��!w��6ߎ�ߜ�~�Z2K7�/\͎�Ӹl�?����iǳ���=D�-uЧX���m\+�m̴���N�9�b��c�w/�k�)���v⺏��6��Y���t��'�"<m�DWa�D,�<X�h�5�c����rO\���:}�2t��,���� f�|�߃.�s|���aK�o������h����R�ĭu�x���[`���!����,���t��N�v�&S�.R<Ģ��a��LA��*>�ðb�.��r��5��Z���Hk��$?�O��X�h����LP���*>�1������̭w�ia�.�=�3�e��I�ݕS����Z���}_o�?�ԏ3��J10�Q�^HM��>�Q��B0<�Ǐ�?�5^G��R���k�V eS.�_LЏ>�s=Ն-
=�f2���ڝ�Bw��t��0��<�����p��������e�\7�4���`�8�ur�%�E�
K�a�7���� �B\L8y��R=�9*���Pךp΂���YN�Dx��-���ɂ�[b��:��A '1��pd�>�$F����t0�4�'_l0��ѕ�^5�5���k�h�t�s�8�<ڎ,��H��.�1���6;~��Q��w��r��c�/ގ�����F������ٶӹ�"ڹr.�?�x��;���]僑H4AT_��g��X�~�����NQ(��;kek�L���>ĺ�gq
9S��H?�	�\��:j�+�9,�k;��cX;9۴G��Bbby1���wy��n6?�����RV^�h"���X�ϋ޶J7cn�߆��CTJ�Hl䂄>YQ8��*�RK$W�9x	��V|�q�t������ ����vE?{�x<��6�Gz���w9��V�d1�&���' ��⏛�J�7|��}FZ�﨣������y�tP`�X-qa �h���lE�X2ێ�����0����*e=`usbUP��*�1�Ś�:���.¥$�2���u�Յ���cC:?�%"<Ս��b����Dq���,V��M�/*��9�7��/>>��Ý,^Z�H3��2��a"Ei=�0��l(F�D�DuWDZ�Qs�s��M#+$��N�FÒ'�8/�g�ɠD�E-��%' \��"�k}���HX˚~!w���� �[�ƥ!_y�[��[80��/�CU�r4��X������7���D�zB/�,��5�T��p�����K=�H�U��+��.��c�1f3�+�4��({�`7��~]�c�'��kbY��4	LsT<��_��1�a�2OTK�k�\�1.�_����F@3�\�?��{��Eg̉�K�wL��*��c1���x�L�m ��W:<Ҕ����8�5���{W
m�r@��Rj˚"u;1��B���Ȋ9�Vv\���}ۿ��-V�}����c�>7iD6�6�/�H������)���y,����#$�fKZy���O�&&)�7�9��@M��۬�L4��k�*=���&�i�L��ۨu|J�^z+�X�ƑL}"O1�:v�ľ������^;:ms��#LI�M"9۸�u�e�q�o��$�7]W4Y�/�46V����M1�x�5��j*g�J`�%hĝ�9��%-��m�hl�u�U���B��m��8�F'���4�.�ς*/a�"щ#	��s2zZ�"5TKD�a��T�[� z[N{�<�PbR
7���ֽ��qeiܿǚoתU�i��A��(�""�J����R���X
���M�X��*�k_�V�e�� ̔s�8_�(����"�����D�ט�t9ɤ�nS�$I�CF���۹�S ���5�i'W��`ЛM�,H[�q�)���JW}vpKO���-��C�/�Y�1P�����#�*���޼q )�6Q[ة��s<2Z�*t`���}Q�����'�P���ڢ���("h��$ c�Z������<m�:&����'|�����eU�MyS�Ve���#.@���.P�R��G*l��W�C�EN����XZڒ��Uq�iV)C,Q$�L��F�\�� ��B��m�}Jl�ƙh� �w�����n�3.�!�Q	3���8^����22e��07w$�v�?�SK�2���e�J����A�U�	�l! w^�ŭ��!~�C�x�7��9�=�Ya�,̡A_��#><�	@r�k�U"h��;�Y;��I��MԖ�g��6DǍ[��x�?~�ݖ���R��Ƒ{,�e�N�$H� 4�������~��iӁ��=��� ���ǖ؁���T�&{��D�]�g�����{���vQ<Ud�U϶~+�N�#T[���|Y�vś��F�#���,<¬|*K:���K�zj��T;�r�$�q?0�H B,���/�,��M��n��}P��T�rI�[���ؕ3�'�O�������-!�s8)��,朢�?m�/�Z9���Bc��$A���������G!ЙJT({�h�Ul�T�]U�����h��gc�M��X�v�^��y�u�I�s|_w�s�ZY�Fl�;j� yN뫳���K����x冶�?5��,��-1�+���<bN(� �M�����
V�R��W���Q�srjѧ�����n4CM�G
jm.VI:�*�e�b��ʺ�y��%�?���4ө ���?ȣ�t�uY[�V��	W������ٔɒ�`Z$2����r��0_u���!����fjO�Z�����?��M!�J�Ր&].������9%��1@\����|���K��f�o!>vxq�u��F&��)2�"~3�JS��V��崑����b�h�w�-j�=_��=lŋ��MU{��;8���LzA o��˞���oKu��$�i�&�g���"�JI®j½3�cwۓ>N{H�%��ᴩ-�#Hqnbj ��3@�����9�Q�+�١p��Fw[��8c����4ٺ?�%����5�Ay�K��n�pr޵��3�o�1w��n�-�3$ʁ�J��W��0�@w	JՈ�U2�=��i?!���{W�����|���l��v�j��웄��(���hd�Y
�br!<�t�N We]��|��g�dR�FaR�̠�6'a���3[����}��&���V�����I��9�� � !��ƚ�D�逯���DG5n0�k�MT6�ϵ�V��2n�m�f
�	���ga��K2�X�g�T�f�1�񦏭&�5BEP<��ߍ�]�&����Az❒��#���FK�OE�����;�߸c;���U��D6��v{*�������G�p�O8sl����+���2�:C�W�C�z����|��,�����q5Td�g�V�Nik����\Id��u��~�X ���� m�2E�9	
ڿ��X�������g1a�C��=��-��(]�f���'>c��|�t۫b�#�CtW#��^���KI��,tRGk��V"fy4��4���2D�dZ� ��S-%&Jaͭ.���*�+'�����^ު��7�w�`�I�x��Nw�A�L��ns4�&cvo��[�g�$�/_�!�F�[�} �S�N��x�&+����0�H��p��S��@�%[�&>�����ǳ�2ֳ��	ȶ���K
����uD�A��^���.�vKf����q!/��+Jƙ�ڙ��_�q�<O8�����)4��>��QaT�^��*+VEמ�`޹ԓw�wt�$�P�ȹ�h{nmx^U�;L����:����6Z@��Ә�d�F���fi������D*��g���Hɗ��Y�~9ƈ~R���ir���@��H�|~:�>I�+w��Dc{�����F�c�sz����3�8����g��ݼ����;t��'�0iC�`�@��y�j/4%.P۷W���n�����ҽ�n�s���n�}��dw朦��������.���2���?�f��`e��n����<�˃\F�)͞\0<�2��S���\ڪ���<7
@�~m��� Z6�_weT�~�{-��������ۡ`l��S��{�楙�j!��E�W���ӎr�]Ld۴�^F�b���Ȼ#���v�56�xq{D!I�Of�#m6��"��ԗ�A\�<�z?WlpGS��>hA̐"��;f���.}��8j�����yW�Y��rH���ucP45Ů�/X'�;����h[0�Mj����x7��ԧ����$��3� �oM6� o�O!��,D,����?�=�V���@v$�-b3��Pʛ�a�^��!}�UB
��_7�ur5K�t/;X7�OE���23u{�;���S'Q2pr���6��:i�،�Y=�{׃Y�t���ʔ���g��_�~B7�uL����ϙ�pU��22��IT�Հ���)��F	�V���W�Mi�*���.��[�@�?E�Ah��O@6c*��2��6�>H��m�A�.(��$L���u�S;sIy�;ܨ��?'� ��[�Q�fRZ�C���40��.�u���v���VBԊ�x�ˀ�=�AVƆ�6�h�NGN]<@ȇ+2�lc���V�������<��TI�8hX�Z�mN��O��0b��}�e���)����QKI]s�p%�?b�����u�zL�G�݃A.l�uݐ�Ѳ��(T(W(q��:+�l��t�r�-o&e�=��_> nTZ+�ջ���\N�IlΜ,�=����/$Î��^�����m��Jf�6|Jqh}�wV���~���/q���4���z�TC<4�ض�0n�^�N�˖C#jC;��*��T�5���]^��0�j]X�zp�ݫ(p�EΔ���.b̜��g_H�Ӡ��قr?�׿Ui.���� ���v��΀�Bx=�Z����,���.
���?m��h���u����<ٮ�e$���&�9Z fۣ�y4��Z�F��B����j0�$�J�/Xt���O>F0m�>ڝ�Nk�y�	� �\�G�,��ߨ]t���*l�D�>�Z�G�Fv��}s/�b�nH���rM��oeqA�>�y�&D�|K��C�怊���`�O��#��KB����v�ӵ!:���ǥ�q<:�������c�����א��Re�%���Eߣ;�&��T4�A`�č��[�%Է=�iy���ڼ����L��[�������;X��-�D9x�|��qM��:U�+g�m�Ѣ)���%��� ����z��'�t!�%8�V\�]̄CV4[-�ނ��-���ʟ��3�_(���Hi�Th�b~&J;4����B0�/,ۛjtjjM�7/;oXo��y�X��K�ф���+<�Q��/�z��d5���^J
N��Jƕt��Cs���F����~=a�����b�+�N��:�L���:�XG�X�A�.SO(���4c\iR�>�<g���R�$��rI:�M�#�'��%#s#�������>��ƿ/
�Rz���27��{p�T?�Y9�=�|�Ui�b3�e%����۔Pt���Krp(=�#�ޫѫJ0ox�i��h��=Ҭmf��~S��=����X `��whD�G��q���2*�\S���>�B; �?K>A*NEjI�&0�F{+��!��Ai�\@V�@�ɴ��}#�s0K��[����^���>l'��7W�բ58;W��c=4�{l�K{����m=5�g�1�5��i��$���gķ��U5�5�W23�S^�TN��|]���E9U�(��$�u>K�S��յNe7x�O+�MJ;V5r�[���a��< sV��`>�W��oY�1�x-���J?ɘ_UN4Ub�� ��EТ"~�m��UK؀S�	��?��I��|���ȬW�4�h�����3�i*�7�f�8��me�Ğ;V��*��ǡ�������,
�~֌�6�p��O1iM0�W��Zr��7N����6�.�Ƶ��d&�b:+׊��wPЃU�h%���C��؜�j|�z������V�Z$��9�l����c�m����$�Y �!��2	�aԅ��##/��69̌I+��v[�J�(�������2a��PG��>���J��j�QB���g�s��e��r/��X�|(S��� � ��ɬ�8�x��S���;M��~d�l��O�@]+���|�bɱ�Z� �����-��������Z�8����h>򫞾?M��]�Ė�zj��I��V|ç�5�7�O��fS���6����%�FI�8\o%�Q�S�2FWy���V��+����7Z�>��Q&��ݺ+	��|t�vp�c�p��}��	#CI���	;����|�X{7���<aL�q]��{(o"^;ߌ����F�"\�r`��7�i��2�$gI�]o=�bXXY; �8���Lh���1�=ah溟����L7�1��'�����}�2�-V�m/�Ͻc��C3��y{[sxf<J%H��QR��{���"��#(���V�:�T
���c�, ~>�h2�b^q '�?2lʞF�v�D��(&?�{�\�����lwo�ޗ���r�w~�:�Q_�2
�X��q��-@��!Z����ּ����	=�C )O]|%EkT��PH_�=��+��v��-/�G-1�{:B&z��Qv}q�l�w�	�{v����ٜ{ԏ?���3�ӭ�[���j�1Ce=6�GF0g�x�V`�{@�nw��]��+���� �u�S���t�ʨ*�i�A4�>��l %S*v�Siݮ�n��;�q2�����E���_8���sW�nD�'RhL��yqÃe�3����Wke�LрC��-8٭=@����D�$,��P,UN��$"n���0J��,%*}�ؠ��,��+��M���[rA(F$_�,���_�@�E`N��ט��+D�I�~�G���v~����X�ҡ	���F���"��pB�$��mn,�� Vk�}2�>�E�������+�NOS�!ӯ��b��V��E����>߈r]S3�*�x�y�\evYxl�S� �j����|v�K��2��x����Sixm���y)��ҹ7���u����|E���O����S��eg`Z�������̂�r�#Y���'�p�6���-z���.�����1uZ��Y�5���Ԉ��"B<Þ�?��!��4�������4�/c�춴+*Y��Y��7^�:�	�V�{�*y{�%���C[T��d&>�]�wN_��.Yh�(`�t:Q	bi&;�����nid&���G�Ϝݱ=ɸ֟E#_�F-���w���ġ7�����
ђv"ԯcHr�$�q��_!};�Hg�׆z,l_��5��$Ɇ��p��������z���B�8�]$�R�Ƞ������_�+�cl�-�	E"Hn�Ժ�J��=�9� B&��,4Ī� ����0�T��2~����)Qd��b��&�C07b�A�U�M߽S0K�Y����f4`�j���PicO��]" Q�a��S2��2-�w1���<:�p�
�G�r��P,�ӷ��2�72fܸ �(R�=�|ݍ�V��]1���A0@�n3����`u�Z����D�G	�Z�@�������@!�2����
�W��ߒEC'�{�Ky�θ�)X�lM�Ao$	��6s;�I���CA횅�E�1H,�t�A[X1,��J����b@�:l�|DNal3�K׶<��#-ɇ�d�n���g	���5V��š�B�U�-��UIq`B��D���z�,��f�ʅ	l,3�IaV����Q�����pu!��@��Ƶ�yD>RIԶU�A�g��aZ][�;k'��l��u��C���_�6njI\�r;&
�J��PKZ'�b{�3QA�I�2V0ɬ�d�i�R1��Sd)[���i��54��$��V2d��i��i/'�4���~1��f˧B��/ͣw$�H�p��LN�ʕgt�׷���)e��N�o ^C`��Ma� �H�S:�Ԉ,�����	�;n���i�[pJ��_E<˦#\:�*ev���xO�	Hם���ա|�pd��G���h�1�.Aq�4C[�� �@�aճ�q&��11î�D_�FϱK1c����QX���Iî���f/�5Szd�Pm^+����n׺g4��f@Wn��x������F)��S�鼴8׼f:L��Ǯ*>��$k�H%������7;���BX68Bp1��q
+��]��?���lTcAr�s�l�m K\0��Oe���.1�+P��#�����|�5���33�S�~*���*KS!�o��T-
�	�mX�F�U��Fأ6�&L�������e/���;����.:��]���m�\���j=��<|qk[�9��d	jh��Rs�=�F>Ƞ���nֿ�tFpj�#3y��4,�7C>�v/|qh��s��Z��PJr]����j��M]����~d$�Dc~�̂�!�*LKi�u��O�\Vx����4�\,.,��vkI7�;�'������'*Z��1��o�̤�wR=�u0��[j˗>Җ���P^�����m]$�~r����@���2,�,�P~��ԩ�i1�C��p����{Ё��峔)$
.�r�x0�T��|׊vԔ"�Ub�®q)�fD'I�Н��l�{R����X��8:�Iw�T�
��i8���[�8�m9@x��6�q�䮮�5}	a��С��r��yS��<����1b�=_H-�N���z�"OR��󭼮;�*0� ׯ��M"�j2b��Ȫ�`[.RI[@����r����;JoT��lbG�A�'��A)8�Ť�D�����H��sZ���քX�1��J(��i�G7,5şɷ�h�>0ֱ���M�Ŧ��c�4"�����pqw�Re�-�s�d�̐�ԋ���$��V[�5~�BҠ���8L��]+<�R���/�Jl-��<ɦ�g�ݫm�QaSS�8I�p?�U*�f5���ï��̩�I+�Q�dcTz��'�P���T����[�ȞI�$f�xM���S�K���K�A�[�apP�����x�UO2;�47�WB׵�F�YS��'����G���'㤝�C-Pڐע���0C5�*����,�����Ԝ���.F�fKp:��G��|�����"�"N����CPt/!N���Ļ���p���;�5���.R�����P��"����Uާ)�ט_"�� �xwKVT��Zs<(V�˷�b Fq�Ֆ�w����.��������Q*Q�摀>��^�+�?��A862��E�4A�=����|��I���<U���)29���@��-D)JG%8�R�=0$(�q�p���$���g=R{i��SiE0fSm��Z���e���/�Z�FEWa��|#Ӆ��8�Օm��p�MC�D~��E��dk"�rӹ�u��g Oӆ���!2@.O�R'M[�;�/��g�/q]��A�
�9k����mNE:��u�NvM��<�����a�>�eY����`NpL����u�C[9
���>���M/mm�k�[@h_g�EV����"�6��*M��%��7.�co*.��˳�5oBxA�W\�XӡPE�Ӧ[�Jw����_�8Y��+Cڋ���nTɕ�U*�L��^@�<}Űr�q���p�v�"^r;'������z�J��	J]l]��4�
�dב��6:�ַL+�1J�Re���(���!׈>��2�����23��j#��ܞ9	�x��]5�}��q�b�� ����l�_O�}(�2&pR$b� >,��o���%W!��2�ʛ��<�O!o��8��8���dO�u�_�`np��M�0�����y� uÄ�t�`�nb����&���M���H�#�Ҡb���1�:�	B����NHMk��� �-����dڙL�MI��a]bm���WlX#b�x�M��j2�ƈ���(ǝ��%��^N����/^l%Y;�/��&-�(>�~uM��gf�kWa�������s�!R�l���C���#ӥ�����՚�E�