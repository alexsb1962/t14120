��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aЫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�g���)��V<Dr��F�@���ª�ƨ���������;�4Β�����ǈ��\Nl��;��}����MF3�+u�9z�E��y�!i�]��Ie�E�w�����A0�<'�x܃����ĳ_%rfע�mk�Z�s�~�ǀ2#a&��{���pO�H9%�z'9�\��ewm\g2�+p��zBK�w�gcu�A�;x#�B�G<�CA�L�#ܤ��nHA���!r-�T����g}Xc�m��7�%��pg�N�S�o��9w^���
� Q�f��r�z��pc�FX�u)6����ά0�Y���g~L�i�����c��l;J{�'�����hFWI@�w���1mC��ע�T��;��2���\*�������.)����=�_��5�R1av-\�'�0�e��_f4�H��lV&���kC-��z�'����M��(�I��z��3O�46����X���Ne�]����0}h
^k���>ٮүm=:G�h'r��	'S��#���5JRJ�lhFK����������o�GU�>�hj+Wy$i�/�l��d-�X���_��˫���}>�j��Rn�]7��G�q��u�֭ot���֎{����g}22���Y>�a�,C��ި4���$q�V.�GDK)��6��`��ԣD���8�t����`۟w���ͣ:��pW�ZG��I�5�3�����^�q�fX�"\�f'����s���	��"u�0C.�����!�>G2��7U�Sމ�Ie�_<(m�9��,s��J�x�!B����Jz���)���hC�����k�ZΚ-
��-�a��Kх�uxy|�M�����NG�wm�74Y뺣6��L�$њ� �Tp��ɓ�^ީ�R������%���7���:��t�#�[�*�#�<�0�U��׮ŕR�=sVl�p�ɻ��VM��bmvcZ*�-j T$���u��I��r~���$����?uy�'2V5?t�'M�~�26�7�˚F��ж��E�9�w�:�m��q�*��E(�D�N�īKc_�����Lsg4���,��D@�)�c݄g1������	E�~��7�1�o�]���,?5Z%��XY���|ۿJ�/d\�~ʅEz�#���	뷹�Mݏc9K%P�t�\"�S�`Q�
�>B�sZ<�ڛ��*-�i+\;y4�Q��8�gW��Ǔ���:�s��"�t�����Vz�WZ��Χ�!���V���J�B��8��[�d_9��jP��.�\jNޗ/�Q�vO.��/������y�_��ﾗ������\�(����3L�:U�q���ĕ&Q/�������Fg
�X}U+M���E����Z�{�=��x�k׭ֱ�I��3��.z�~o��[/�)�����`��ǔ֢?���D��� ���Iqg@���Y��Tb"|�De�����1�Q��&�m��h`���pZ'Es'�p����q=�}�	�>ßl��E�0��s��8$��y�+߿E.V�َj)��q��`��fp�H�e�7�0X�KY��0�ʒ���ǚ��Ӛ��l38�D��y\tŝ�ա��K�"8K�"dhd�>��	�s. K�0|:�%�\'(�e���Fո���5r����;Ek�|�p�`����`�u��p+p1� 2�&��8�_�@9����}W�5��$5�A���袞�R���0��'^������ؠ7փ�BAK`lS�Kʜ�.�-r�����Q����$�JT�˭I�����X��ۀ.@g��Lc�KD@����p$�������RGo�B�V/���������>�HX8y���6��q"�u;��5�
������	���H��dYi�Ϳޠg����#xJz�Q�@�'v��K�9�=����%�}��������֮�3���;�ʜ32��U���0xL7�Z��^;��������z�7]�)$G�ٵ�����fZ�HH�r�����k@KL<��,��_�ćY�/Yܲ@�`��� �\�8�����fA���R����;�К�l�bD�fđ�y&V��=Ab���Eq4�f8[����Ǻ�8�ח���  �Q������U��V��_`�EE ȕC�D4m��:dX v���Q*�}J��;�=qd���k��F��Ⱦ.-4F<�@O�w>�WԴy8��YkiO�6Q��Ǝ'��g="��.��;����>O�J\Zm%c�qd���}q�"6c����n�N�W��E�ؿr�@��B��H7��u�z�b$��SO���w�˄�]@���9��i!��������d����� �w�RsIu6�&u�Bkѷ�_�ӓR�Bl��8*��-˵�$�˲�~쮔�
�_��2�(����N��?d~���?>B�9�L�r�=���k�Q�Ie-E�G��r܈.�C5��뛟�
�h�ӥ�$�?Kie��΅xG�����_��,��~ X������C��Q�}3�0[n*�6�J�YI�������o��7��.^������H	��a�Jأ�2��Q��⩲���Y#Y�L�̜O�hP|�~ ���E�*,�2�%�ɏɬ8��h��UX��jU2�:��~�ݩ��ΠMZ��n�v$���ҧ����؜At )H� �����<�c/g��	�?3�j��ae��c/8�(�{tJ��.��T#ʤW����	���PX,`?Ua�"�Ա�����4�A����aH���M�#�����<5��a�0��8d�TS������
{2�g5s��DD�eWp@t����!>r��^^�ubR�4BaK�ސ���]�ˬ���ſ^dݸ�\�
�t6�%�(���r�}�Na�Y=᪗9)2!���C5�%ș4��~�}!�mu��W��)��:����#���o]�g��$� ?�^�:�]]��?	D�%J��2(H��ؼ�f�UԋhX���"-]�b�Z�g"�v`�����b�� %���?�?�/%���Z�ĵ4r���b�A��iv��s�y]6�7���]ђ��!Os��-b�lr����Uq��RF♪,�=>Q�b�?��w<���0���օJE�z������
���hdEYs��:��Ҽ"/v�軡�}M*�5t|q|ڛZ/P�becڱqv�*�˹��^�~g��0_n�"��{���6P��P�k���|��:�d
be[�B;ǥe�G�x�3~�4��۾	rQt��.��Ĕ#���8Y(�b�ܮ�n�5��$���Q��k���9(�<y7.���0��z�&B����/C��q�1)b����}u��"�"�Sǳ��3֍�t�$��������T7�j���Q�ߣ�.�ld�Q�(%�d��c��%�T�E2�|�e��p*�gz��S.�b�?�_9xwk�bY	9�w������ �܂��І�DU,��&l���%�k�G7�uE^%QjY���	T��-�G�{ی��&�W�@�۶�<h��o����Eӵ�F{�WlP�r��G�0��Q&����""�w|���E<;P�0���G��2�m���4,
r!-IYZ�g_ͪ��ck9&9����!�<`�Q9%&��`A\����K/�(�,����*��o.`��:��xI�4��Xe�<�⩴�7͡��i�@?=*�Q�nٻ{��!}o�]&�Ƶ��E��ôt�	�ȳ=�<t'�(�W݁�֛7��b�+T��ϵ�X
�<�I��[���^�uU ��\�d'���=�E��}��X�������<�`J�Z�iǲ�l��!إ<��cI�8�Sw�t���-��a�h��#"����! n�R �	���pX�/�s9u�!d�&�O��ֽ������cͻ7�FyJ6 3S��pm�C0�
�����	Gǰr�5,؜�/X;;��v�>��߈$��U�5�^ʵ��H�vSX}�������޶d�C&n����kڤ�Z�Y�}p������f�5x���ڌL���V��4絴}�q0����޼TsǏ3G���}���v�A(��N�m7�%��O���]�73d�Ȥ�"�Рi����l�<a�7�3��Z��K��M�_0�GY��;�����w��Y:~�{�钬B�mO,!'5����Up������w��H��3��ד�@�K*R���a�rH}1>��\�vS�^���Xw�Fd-�#��}��>��q h8��Y�Yp���>�ҋ^�O��a�� t^�-Ƕ�|<�%��T��y1PŜ�J��|��$�7Z��U
w�">8�(ND�1���)B���[��[�.�:�tL�B����	��d�n�,Q��i���*l6殅���@ƅ�������_D�G2a�W2���HT���gg�E��"��Dq��q,�GK̏�����1���_�!Ƒ*�����t��`1>�g�3Ӳi�U�L�╈o�\��]˙I�wM�HcV�C0�l�S/\�R�R���g�6��`�1a��z[�=�.7�:��Ӣ!:�l�@3�#�p��������\}���gnqKBkߓ%OI���b��?f�������Dp|�%��3k�uN�$���0����!7��(�k�[�V��ާ{V���72��'}�<�1~�X;�LՐw�ZO�Րp�-�R����&!��n[�;5�|��B	KG�*�H}u�c� ,xڙqK��Z�bL|�`JфZ��)�)<̗��|���&%��~I�p��_*�"s_�|�`7P�/4�����\*�A��X)Az��'zɌn�R�"M^�U[d�L��-���@�aͧ+�lG3�d"�G��4{�\�J�:d�����x([�ak�N1�6������ٓ�ÃD�[�,�ܨZ`N��&�Ȯ�N�eul#�B��<�KO�T��	8vI��`��>1`!	�4����%|����s�����n+CLH���TQ��;�.�ED��y~���!��y�9���5��&-���/WKa��D��#�,E�X�Z��h��^J�Ɛňx�@)�p�=���/�*U��*m~�FF���-��L��&��d���$�p%'xbi�t<��x�/�	���s�����^�z9�D����q��d��wJf�Ssv�w�Z�7��]�� 	�%����o�<2��&9���-?w�#[`cov�X%}�s���tNe����5�ήUv5��8m�+(�\��_W�����۰6�~��R-�؂\F-� ²p���R�H���S'����4{-�
��\�U� ���	%B��F��=?���+��H�6�4�����V�V�3R�3<s�#�Ha���}io+݂c�Xc�2 �~�h-�w$�#A������U\���7�u>�	�Ec�΋���,�ֻu/��5�VF*&T]Z�p�W����:�Ŧ}��z�hQχp뇛lJ����Plko</���:RC�s|]$Q���R)�����U�'������HNcuُr��KAjE�`�2��HO[��^��=���8��8I�=@"#���R�����֗'$�Zb��Ƌ��R{?�HdS;�*�a��j�P=n���؀<F�wH&Ѳ�	S��Vߙ�5��]"�2ĳ�fc|!��JEA%A<c�����b�z���R$��c@�V�(}u76��,���4��"ƴ����VVH0W1'��$@��a�H�0ox��۠*(m��[t�'K�,@y��=�P�4u�r���FB��]�Z��3o��vA�	^�a���?B��v�Ǆe��A�d�o�P�nbj�r
o�3����8#Dد��� 5P�X��D�/����ci"��:pK]��-V�
���c^�4G�A�d, }�	����/�y�3Y$���d��X����O҅�#*�;ШU�#0S��.�i���pμ��`l���l�,�E�
���Ȭ�����98q�P�V"%[�O��Ϫ�'W!b�ދh>����A�5j� uwB D��4���|�I@L(�Km�c��Ԗ(a�.�i���k?"�^$q�G!.0����0��Dݷڑ�LJ/�5`��Ф�SP_1ܶ��r�N�Z)��{O�XQZ^�W��1���������߮p#������;7�W��/ޕ�N;[���������� N;k}9�Z�(F�˴�-�T���ڸ:i����Q�!����&�4���[�y����xd	hY��h�׵��n[?���{��2ֶ�2㜾7!�_VUޭ�Rh*"o4�H*�x�@l���Q9�L1�z�Y��o6��`x�����w�v⑑��A?z���}�=�v���m�5��;|��<P���}�q��Wz�D#��C̵����ܙ1Q!�<�8�W���7��Vs�s��vH���{�LvJ�$���=�0ov�xt\�N���9�����~�� �E�R�J�E�tr�K:�)��"��i��H-<�WG��|3S���Qo^P�rCzM�N��T>���S"�*�&�ٶ?麸��"^ڳ�5�7ظ��$�~�^�zW�Z��S�k�e��6(N�!�9I�8N���j��Ҏ����KjJVJ���삩�Ƅ��c�īJ6hb��`�C�%��O�R!e�UA3�d�W4�f2��X3�3�M �S���	+F�����~��,@�����o>8�<�9I�q���Ќ\�g����>~>IU^:N��(�\=LO�$%$�7�lPH.O\�1�� ��OOo�P�����c߽xY7t������{�å3��)�4��J�/p���?>��m}�P帰v9�	�9m��W��|kY���&TQ���̕��e�~I��`���K�1�a�MEn\�Ԇ�����"Q4������y�*:,��=�6a��p|.x�=���`Ѱ��^W�g��}�M����	�q���&�m�؟J8��N�f�Ũ��x@�f��-v��L�;��E�Z�;�������'���&���Scå����8E���QϖEO�8Р�l��a�~:��[S��!�x�={Xǥ^��[L���.��ݻj_o=�����IX�7�� ���C�L�i7��:��`�����-#��v�:-:lDj�5P5��v�S��P��&	�ᣄ9jo�"rb �T�3�(�.d ����<�(�l/:��������6Z�(�;�M�����b㔴��~�d��Z�,|8e�0h�����8�Wu�'�u��%���Df`�@�P,�X�!@��<��߶Z���a�פ� ��6�b�� j��}ǌ���tE�Ox����,0�<��ǕK�OTbC�}�[pUw����׍I5x�\�1]�����y &6����Bm��=-�p��U:���}�?q,x��x��kF�%_w�rXZ	~��C��F݃�f����Ȑ[�'�7�[�6�y@��y��
��e� xR˹���XZ���? �ӱJD��ĥ��R_o�J}�����ʧV��`� �D��26FV������g��6�b;�K�`�v�����u4�Ѭ���m��Y�&��m=)�@�1��=������	0����K̎[3�K㣜,B��,
��������z�k����^^`�5#����eS����;�l��пq���Ӫ�_���C[e�?X�:��!ҵ�8t=��ƥ�a!%qm�u��7��U�Q`/�m���!* �G��ҵ�!�cB�^�瑨p�:��xS8!\��æ�<�w���Y��Ý�U ��2eӀ�z�éY&�1�Fz��P�GK�-�^��2�!peª��Z�ԜA�Wd�X#]��K����D���]N�*���䤷k�H�*|�Db�l�ÑlU�CW�X�̵^�g�Т���|;ѰE�S��̹@�-���ŋ`Ռ�\���F�q��~t�P_��t�LPf�a�;GI"��
���ƾ�QAU�H.��������F��(�@4^��y+��F<�D�����y��8��w����8ga\V{�)2��]�&��bB���)��	݆���Hq��.FJ�)!�cֲ��*���&�Z�R���>�NYf�[Z	ݬ�8品X��v��p:�J�8϶%,��]���hd:X��aS��٧h�^-��4!h!�9حn�K����Wq�7�G�YѸ\�;j/}i���
�o㎨Rt,��Pk��]8�U�$"h���$�	j_��k����BØ<@��A��\��³�p���tHt(QZM��A�u<B��{��ꅠ_)w�'E�IV��ق/k�E(R0���K7�3W�"�$�_�͞VOC+��z���W��W�f���꓍�7�D�o1��!��1R�+HY��K��'��6��߆6x�Q��,��)�_�	]%�Z���f�9djC�N��)�@�TY<���H�+Y��.�Cn/kP
��?񮞂�ਅID�:��]�j�۵����I�i�(�{g�q&�6%��[�Б�� �@|)~���vYg�WZ�#S����5Z!���S�ȅWɩM���*p���+�=��EM���e����1x�*��٧�Z#2�;�Q� �����EYU�����8er�s_��2`����E����',���|�&+���>5I$S�8=h��r�YʠTN�q���%H�|�J�k�^�!�uU;	�ёaPJ!+%�ǥ\�t+� u�e_V��V��4���B�r
d�l���Т�{���ئ���םn��Ԃ��̞�C��iJZ�Lƴ�h��P��4qm13�$�@}`��g��i�	�J�RJ�w[�+ ����X�v�����Du@s�8
Q<��yn�#��� �de$��)��W��+ǟ�P�*����VC����wU�;	�d`��׈�7�hy�x5(��5f�w�N�~9l�܏���{�1��1������b@��@q����L��K���8c��n��6J��D��J@��s�à�	>���XoY�Z������p��hY[ޥ�*/{2[`^M!�P��т��(�e>�OQP�t���2+b7t �i���7�S����	���X
H��~a�'��T�i��S�����E��mv*7J�ʛ(�����n�4�!5�M����n�\j�ׅ5#�)�#��#���\J�o����
|u��ad�E�:Z�7����@����qU�y=q�&4 �`����������7Ca����<��'���<	�����`f��aͣ�)�T�37��b�^\Y�_㨓���6����߲}	sq?,urp�Wl���Ҧt~�aѧc�ЩvDÛ=;
Nh����O�M�NT���8ZC�,$PR6��v��,k���A��d��0n��M)g��qfv�
�ݴN����sC-��٘S9�ZgE�@�S[��>xD�k��io�ф��
�;h|S}�#k��BZf�y�z��x��#tq�ܻ�~�\g�ăyH�'r�̯)��.�}��"�_�P��5B	۸�ζ5�lNcW9R���fG���¹D���A���1�@-��eG7��T��k��ܯ�z�	�ݞ�͈������w��Sund`R�hlv�#�3ʟ �Y
��&����_Ǚ�$�#U�jI�[H�6KM����:-�%z�6���*�*�S�������R|l������ƫ���+\\�.%�C��XĮw��N�t�!q�,8�	�K�v�6�Q}��m��8�}Lkt�Dp����Z����M����`0j$���_am�:��%�A�	�
��v&Q���MB,(�v>&���~O�)�]��2��@�U��CTL�����e��Z��d���|���?|W�ǡ�=��r��/~�1J���'_n��	�t�@�s���q�PǙ�'`Q2 �:��\�GӍ�A�kS19�72�P�AM�Z�=��0�%FϿ����C�z�൶Ǧ� ߋ�jc詼���G!��	�E)d� c�����J��
hB��!b���r
�G��<������&rgX(���p<uX��`�F��:�kk��th���ha�o���Ӯ�:	����Aӣ�! �$�ʸ�ދ� �3P��L����5�[��&��#��l��Φ���$)��l��M�T8���E0X�j�(�����ט�����u�k���&�]�=��r�q�k��Db7I��NX���jiK��ܮ��8��))��T��Uyd���utP�'�o�R��,Wų�A3픻/y�|ޝ�j��+\Eu�e�����2�ʞ�g-/X�"����.Iz��6�o��V��{�,<�vc��u��02�����T���~Ə�ᑭ�{���{`����1T�*���i^��<�I/3B�)�d���}홋_��3��������3#)�c2�����"!��:r�3��������O3��Ю"�ڽ/���stVphm��^��c�����/| �|j��E`]1�G1)=\�B.?�ִJ��)86� ��%/2���M8	��V��)����m��x�(����&��JT��hL=K_BIVa{��Y��}��2~}���'��ph+ig�Sԥz�'��gX�R�����b��_ks���D�`� ���&'}�^�hԧ!ѾX�!Ih���V+@�D\�V�ĒW$�#�y��Q�N1�{��.����&n�Ȣ)f+f��T�F�Q�D�n��G:�2%�-��
��MW�f��f������_��_�À�o�����(�-�b� 4�&
 �;I��'���W/,�ye��WC桁���ߦ.;��Gޓ������A����Zit�	��$,!9&�"�$%���8�R������*��&E��:�7'G�'���k-�jKѴ�7�㎀�0��ps����6g:�[h��8^2��ZS� �Ƴ~�$�R/!a9����p��[0<�-����׊�#�7��+�c[�e]��-�(I���	�d��y��u_bz�)�C9hδqU�uH�PƢ@e@|~����ޣ����YU�G�`�6�<ܐ�*���q亙v:k�f�)V��LL�$?o�}sÎU ž�>N�4sho�~�P0?X���o�Zp_�-��Ğ�#z*?)��6�⁵�%pi^�����*>K�5jddK�U<C�uI�	�n�;�P#�M��q%�ր^B��XgtB��X���|�+~��Z2v�^����?�kyE��Z
�5R��S�>;�"0��9��5k2����"�y9