��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������;U7��б]��uL����x�z���^��:�q=�n�[",v���@���Qh�c��t޻���0S����b*�&��@R���Af�/��Z��:@w�fe�5�p�[��V�3U=�.�i1iJ�E�����Z�U;��~�%L4cK�d�����bneɥ��sˉ�i�1Zzͱ��N`��F�?'+`��O�9[���$8�Tz�1\j�JWaN6�E	��tj8~EC��s�z�L�H\����!������߬��9�w�E�q�86 X=���/(������f�
<HaV���6�����m�mχ�:�H��"f���+,Ü��־:~�6MJW���0Dg+�-فL@�E�'���!�=���Wu1��bG�?�2���ՐЦ�ʲ۝=���k���&���J�J6��z��h%���b��Q��Xf_u=P1��cJ^�����C�ɋ����85p�!=	Ƽ���:�B!���-��KFN��~��aW�@� *���I$�1���I�M�?��/�3i�,�	Ԡ���\�_�M,G�46Z��j�R�1��3��\]��x��3}�l5D�gZ�0� ǁ���$��G1�kS��7�#h�Ba���4����7O#6~�_e�,1�[ CCy
��V��lv�~��5����sN�x[�ʻM�W�I��㘽��x�ֳ"Y��&6¡	,h1C�x�CD�Sҿ>�D]�P�ىLm/�)s0�c���@���rY�Ύp�S�qN��G�mZ˸�oԕ�5���ϒ�W�*4�
�g
|�<���;{��)$�I�2;�6+<
�c�}&��' �)e���U�*��iqQfH*�������߾�&�d<u��(i�id�7WZH��vo'oR��<���P4��rn����_�t��� �	f>��(��MX#Zx�'��� [p1x8��[h�l{
�zV!�ϑ�!I��L��	�扔u�չA?����a�+������i���)�#���<��r�����Nf܀�ȕ}١P�GW��..Ř5�:l:^�V?��]�/w0Q�
���X�h��3W��t�SA���tY襄G���'�:B��7����颀��=�ؓ�!D[$~�����S��a@@%_}-�׻�6���#�]-���_��9�A"n��l�)ݕ����#Gd&=1�����^QL:�x���˾�(*���7����<6ŵ�����ֶ8gٸ1�(�`�˕��K��%�͸3 �ܟ�?h>}��?�vU"R�>��PF�	��}5B��99�^d|&��?�U��ۜ�;H;߄���^�K�B0Ԩ��1#�(�a�P/�����n�E�$��kդJ�0����z`�s`}��=���&���V����R����^2��FX�+��T�m"��Z%��~��
�EVp"��D->H�<#���Җ�:�l�:п5��x��'a�-,gH�+�z������`+����E���A"s�<ׇZn:�4���S��FH�a@E�T����8�����K�7��T /���f�od��hvYW�ൂ�:�@Y�b�}�+@�uh询C�H�n�W^��K<�"���ld�����qA`�]1�j�D�e���R�B����q|ه(&������O7��~�J��M��M]֜�b�Ͽ������3�k�vC4�L��S��z b��5 r����I|k�lf���L;��y���}<�Sq���bj�ߨ@�k�����m<�����
��YیM�� !O��:X��}˃�~�X�qYd�O�J�b
X���`/�Ԙ�ϼz`L\+���3��:����I}DM��ǲ�é΄.n������5���h^sI�T�5����:�6N������[��>D�x�*�f�HI�k�U�����$�&7�H���2r2*޴����j)]�2ӃQ�t��f�{P�,	��P��o�h�q ��H"�B+<��0����o�s�ŴKڵ�0����ٚ���~����d��-e/���
������|����L���*?��)��j����#�5���,bBW�~�}w<�o���_�k#�f��Ȥ
�C�.��~Z.�"E��*��!
�-\���5$kN&�g��J;�:�ѧ�����h���d���P�*~�J���|$�Y-f	�����/�K��x���c���NBu�|��T�@A]3����u<�9*�������|P��o��8��Y��nz�)��"�i"$j� ��G*�d%���Q"�NPX.xAA&��"y��>�SGa9���1���{T��j��	Q7G���?���a��N�
.Q�!�����ݷӯ&,%�j����7�z�� ;z���WppS��dO��~noK{Ar�U1�ӥ��p0ɕ.Ի|Ιҵ���/��a��OD�NK�Y�O�ƿM"��Z�W8	��0	}cZ�+ò�
��-(JY��:��Jxe��`�}P� ۃ�����K1i=��0�$Z�5�V�ܱ=�-�HfT���ҡ�ˣ���i��K�6X+n)9#2)˞�P�.\4���GP�β?b�&�M������������A^b�2v��x�8<������[3�	B��6��a�P��X����f�0�C=3�m�[��Eh֝r���B�T�9�b�uvN̛ٛ�AM�@�@�I���?j�#Y5ݯR@݃\�,���}��53)	� d>ڲ2�M˫�uj�հ �k.��䎛��U3!���U��nt�ن��w0E��|9�_;Ղ��Ӡ'�C1����y�c��`exc¤��?ŧ�R��V&����?��g4��gLvrL�o�{�M��+��]�L>3R`�-MnV�/�G����D��!���ֺH4�f�na����e�]���K�H���CP��i�r��Y��3� �Iz[�]�;��p7��O���S���QO���3H�c�c&A1,���(s^Z�/OH�_��ާc�0�E�#{y�3ʊh5�u���w�ҳ�(Y�F��D�#�"/�rwvԜ���ZԶ��������+�C�#��j���~�O�7b����l6�Ԝp�{~*6��M��E�;�֦�n�?W_�v�le��(m�m{�k�7��I�O?h����a"�`���>ݡk��S��r&�������f)I#�":�S ,�X���4�,;�q����k�B�{P�i��@<��{��.����y��^��
4�?�ç�X�3��Ru�n花܇��Z�����?h�6��0���=؂�z����z{��E"��L�T��`�>���dX�#DQ�����
�А�f�J�Ȩ��m7�/D�����[�S�˝Lj3�c��%� %n[pra�#>�oG������@��[h%V�U����ތ���XJt��=$O�r
����f��Z���4�pm���D�����"%�VZK:�M�k�|���V��@�_��ۢ����YW�:�&�߯���	��Y=Ю�~خ�,}pa��� .���Y�cB��n�S�*sF�Q�J@�Z���Z�v�=#�xj��P�Ƈ�7UO�x���{��6A�MQ���b9��/���q�|a���<s�Oy��~�T���.��v��[��ƴ����Xu��?m�t
�9)�(���֚��G^Qh7�6S�շqmRC����LJ%x�Z2��E�a�2������ iš�U}��C+��h@�h.�c��ҳj���V���u��.���$r���~��e\��ҕ���)i�b�f0��I��M&��ʬ��"�&o�2VI���x�hpx��Z�6��.�;O��U1�*(0��sjYD��.��sK��˃Q�]Z������BL�IGf.
<���y6<�S��jv���y��[�H[x������V��iV�0k~��T�3�o�t� $]`>���(��=�.�qxB��pQ-��ǒz����[ʂUĘ�ıW�NA�L	�'�E�������L��0,�*/��{b(�P�/��_nඒ�oʂ2�`�1m4�q��#��=tM���]W��^�%��e�-�88j���\FK��llp�(J�l߯���6�|�{l��2�݀$��^�B�y�-@0q�V{�M�_��F�����-n�h�E_wF�<��턨K��`���L�;d�[L��!,t�4v���ϥ�8W@^�LC^���V9��J�"�w!��%�:b���Q����.5@�
q���� �"�/v�^���b�_OM+z�ڷ	JZ��Ѳ6��x(�ʋn`H�������r\h�������>��Ћϝ091�+�!&::���	����Y��[慝I��v�!����M�⋹Ѭ�I��}�R$v���Su���1�/ʺ��DR����Acm��ӏ�v�i�RE�'QT�O�����?A�@���5��1z��Bp�*�A�|�gz�mC���4�&�u]ŀ-�\"5v��
&�z��̎���B?��(���ߦy`e���Wf�C.�9�Y���zy ��X˨�z^�Njҧ���8l3��xiN�jʂ���?�, �^?_a#��]���[R�S��0uR"���GI �d�W���T��-�0�ܽB�ꘜV�[�"�Δ�yH�b9t���Z*��=�iԬ�FN�m���Ӏ�C�㌋n�` LVh/3�����B��T��hY�`�ǜ��z5���݋MJ�
��*=��MJ�R%�#����jE(�)Do3-�I�7�P���#��q#5<�*sL���^'r�ے#f��q�	���8 ��E��M)�_�5��E <�\��-���s.0=2��uGj�G�b�'�pn6LWm�0�4�3�9әz��@-t}ʅ|jIWe�Χ;���b͛y����gb+	��l<��"�D����<�b	���H������Le�ӌ�
%uο�G%����=�T�.ũW|Mg&������H�a+��lN�H�}�������V��.��B�Ŭ�nKhJ��k�srR-�1�³M��<�+N��i�#]��v~;�=��&~�d��g�����\�u�i�.�*��6�A�2����$�6��Ѻ`饡����
�+�Jp�+ G�F����ฮiy(>��+}��]���
h☉,h%�jf��2�?�c�kImI��#C\�-��O�6�t�З���߄���Ev?��/%'	L�į�ѡf\+Q�ܵ���>:��,��TMb�7}�����2-i�Só����a�X�Ԩ��(��\o4��*�#���ƛ�~K��$�z�b.��]{�x���OY�72D���Y5��J���-DΪ//���p%�4�<#����vqd���s�M�tgl(�b��h��l�ޕ-�rV��C8aY��Cv��~IF�=��h�+�۱�8d�7�l$?���JΏ�7�����8f)Qy7ѡ��A�\s�>�!%�X�E��xS�>�'@}+�f�Y�:˚@]�L-�H�o��\�6JK:,db�)�ٟw�5�_F��W�
���iI�bg�qGO�;��Ms��E�� ��(���*�,ׇ��Y6���N_���qE�����i��g�2����g`�ْ�{'<�+���l�-�4���*LNl�m��e'X,��n0�
��g������u��q[�߸>�����V�|������?��lK��<� bJ�4��6^w!����aȂ��XX /���|�Kࠖ��ZafY���������(ҁґ��^%v��詪�co;#<�����{C": ��#�BN�/݈��!�=�/;��ݔ��).�t���[���$TaN��B3jS�<kN�L8�
��M ������?�"\��	{���Μ�n|��S""�-4�:�X�`v�S( �Kl�x��.��ݹ�/�t��4&�@�6W����͑ ��u0T�E��R�^8�H�&�$��('�2[9Lڳ#��Ag������
>m��`(p3p�=�_��S`EL�����I�g��M�Hr�|E`򳰽$��Ll�d{|��Y�[��a�d�I �PԆ��Q��1F+�j[����b1u�W�\%qa>�0W4��<(���K����h.wR.���`xq�G�m�~aç���SL~55`���	ӤF������9|�=��)
��l�w��_O�Hʈ�����3T�K�;��_�F�|o�2��c�G�o��NOƶ$�Я�0|q�a���#�:s�b#G�R��MpƳ�o����/!LHW1���D�}`ZJEMQ��s�:l��*6�Ѻ�皠#Ρ(�lo�_�R6ڞ ���6���%%���4C�"�k�B���t≛����䔱���m�(�a`!��!ko��r8V�ff^��$!�����Co��i�p�/�G��Ԏ�d�2�w7O�;�A[����JF5��M
МK�ěݷ�h&�K!�xl���`�8�p�&�9�Zy^����v�$���Ϭd����	�W�i�D�x��P���E�Y��ѩs�N^i�-�
A`�wP#�(��Z�;T�z���ѧ�p־�n'k���QרI���=�XȮc��i>y`����=p� �u��J^	 �H�:��UV�D�7���<`��G��;�N*�m�6&)ӥ��U0��z�W��h�]�[1~�o�<�0*��8��5(K�x�%t�����|fS/���~�
#�D�mG�0
*B�Eң�޳l/>�9i+>9���%����*�K�	�R�	@�^)P����Y��LD�]��}�[Q�^=�7������Е��zMn��b��:�s���֏VkJ�/خ����z^�҇Vعs�.���}���r\�ųc+�u}���]��uL!�z�f�pBko@7]���:ev(4Q���US��v� ���BF�^?�T\�l����Ir�2u�V^b�>� ���
B��Pk��'��+��(`ύ7���:�1[PB7.l"����-��D�0RGO4V��q��nn�}�V;B;���J��?�"�]Dt.��]4&���%�C�?a� f��^*3jmXv�{�j�KJ^���I�G���Kd�}�����ň��A6�'�pѨแ�9���S�Q�ޝ8yT��C��е�Y�<GK�㖿K?p����������#^D��%K�;�Y|��W�����D�V�p�:����p�B�"�ApP,�Ƭh��i5j��{EU���~�������2z�BB�zN����~=��M�Q��0H�N~���F��tz+���=��k�?�-����Os���G�+�ҎT�9⥠�c��cFPl�/���WQ�[�Y�XTz�.FQ��H� �{L��H�h��ZK�ĺ��HY.ă��n3���'s��VEw����#�Ȧ�<����T$ڨ�9rD�f������\�7d�r@yno��$ +����u��z��s�D�(��=�l�9��7��B����b��"�t�S�"����1!���7�M�f%|��n�3����ծ>��dm����k[{ !k
�4B=RyD � �Xs*��E6ˊ2⁜s���,���&"�qތ
·�%�q��Y��a�93���ނrM��Cݖ2�<o�*�W���ERvRf�rT��EL8�;�^s�f��X��oD��˻���i[�(s�Z9d1\����wN����h�7q=z����gL��8Fme��<���r $s�}������^#I��}����a�9)4?��(��:�G��"��}��JU���y�Bd���qcX��߲B�ERx�_����[�2�D�舍���̦4�堕�$����7-��K�9�f+�l���5������eZx��5Z�(&�}�m|��$h�P*��p��k_�[a����Tq9j]���	[��)�9T�lؾt'�q�K�f��@7 �)�"G������Ln�$t{U�����{ͺ*��0�}>�	�s��̭�E(�a��������%��uWVb�#�(�$��G�lA�t㙃)5;���c �߱Rj�o׍�fus'�L�^&k#�iVxR��,�Lqֺ�D��Qt�Lb��@�Oj;+`_� ;�H6�0r�
ŗ@��C���R��>�M�@�Iϧ�zG~�ط*���1'F{/;���p�E9��>�h�zt+ՕVV��*\�g����O2h@x+���hWu�t��tJ����r�W\.`�4T]qm��+��5~�����N%U׵"�o��H�dCin/q��{�:ue�l���������yL���L!�6���A�6�:Jjm���P�'�Σ��k:��es� wx�o#�Q�fyY��Nꕗ��#o_�$M
��$ОE<��.�#�����jkË{B�5�8�8��P8��ml���?~3�Y��,:moo]�",^Y=���b��[�}DY��:+ǚ�}6Ns!(/ω����E3��rέ!"�=g�GA��0뚪0��~�׻!�oC���se�N:�����pTJ��((ɪ���Ґ�7LS �ԡ��5ar��o���̋�=dy$��:�>�K�T�y��P�d�@k���9�������[�!{f	�c!ʖ�!�%@�G(�<�V���Y��^�iQcah���d4BxH�0�z��'����t�������W�N5�/�"0N�'�t0��� �@���>�6��]��b�h��O�#Y���xY^��S3j���v�o9��coX�.J� v������XF~P5�]����lt�8�-�M^��;���RY��/!*z�z�!?��m��q$�zITk�U��X�-��7��� �{pmM����pu�!̀�@��$��Ue�R.A	ީ�^�zN�Iϼ ����9v�X�7�Ǎ<��Wȓ{�=�4�F����t���\�da2� ?���8� w�����\4Ϋ�t&��9��V_t淕���ʉ������=���VT���Vf<V'~�L�=f��G�U�qy����b�59�Q3LEF<�u�v�wh0�h����;�<Np�8r��4so�c��g�2�;;k�.���k\W�SP��IHZ/U�Y�6���ʺ�B�K�D]Dd5Y2����9�c.����M�;e��:)��T��*ܗ,L�m'�Y=�'���M�9|�!Hcxaj:xU:m'�x✒�}sc}lZ��婟�c�!WoC;lybs��$QH]@�Y���n�3|WAb�lf�Fs�zc�pK(S���]��ލ�u�"���CI)��L�lB@�E���G^v��umw���S���X���c�Kr :N(����q�d�J t�ã�������4P0�,�r�s��V���-����Q�KJ{�%㺅����7u'q#O�RB���n��K������������XEDM��8t^�U�:8����|=ݕn�#Qi��uB�C.�u&�0So�{��)>g)���'Tn�f�]Yͨ���`+�GN#�rYݪз6�o~����}�^ә�����O������"2"��� n���Cp�U���A�����_f)"z�q��V��9jĸd*
%�4��NF!�Ni�lnK�c���R�H�Se')_we`����/��K�l<�&k���\�Q}Rt��<d�6١��h(�)�W��5Z�/�Th���잧.�r&�y�P��Z�p�hu?�r�0��`,�kմ�4��w:�HKQ�k��嵇d�S��Ɠ]��+��h�먶�-��v��P��B &����y��q;|PǱ���=�h���{���uUm��op]ܫF����}H�~y����e�
�W�X��X+x[���S�GM�[9 ���?xfܢ�������Q�ڿ����<��v����I��3xz�f� s~�#�Y��a�ehhɢT�a����v�	��!���8��=�w�H嬘/����4l��m�_�5�l[�^x��Z�h;�������kn '�%ā�����MY#��n�BS�Ğ��S���.����%~߶���(��!��Hm�J�m#��6Q� ]�������8s�W�	m8C�g@��t�m�ts�c/s�W�؏ig���X!��O]Rg�W��3�m����Ֆ��1G2���_���ݬX�'�:���t��S�KѢ�D�7���N6V�Z�D�t[SrԔ�@[�LY	���"'��%������ܑp�]�ItV8��0v5j�*����p�)�Bs<���T=.Wύ�i��E���\�I��Q��_`�M����,��>Ȼ�M�u���+\������/��)�8�)�A�L�i)i�����(��j \,O�ѓq�0�Zr�c�MD��P�E��h�^�7�.�W�h<%��q��;eDʐ��&%9�C������α��zas�E#�]�nn��g ΢����j�v#�ћǓ�'8��&�Q�t�l0�hx��`-=Ϭ��VD@��/*O	A���u�-���o�*�\N'? obR�;@�N���R���\��{���XC&>�l`9b7�ߏ������/�d��x* ����|� d�NXQ����H�4�:$����>7@�^g���ǦQ�ŝ>V��8���ǡI[��w=�Tf~�=�J�d�-�U3*ۖnA>��qRc	9�m���\ˡ��w� c���R�9i������W�n֯$�E������WA؊��U��;s��&��24b�@�/�=��E�����4�`�ѫ��
��9�6�	������������O����P���֖�0?ʂQ �u!`<�`�����[�5�uz��$hxL6��Ǯ���b�U�'�{J��ZZo7�(�_JEY'N��Z���%�m�Ѐ���c�˭��r�jFX	�k6H�\����␙N��3z"A��M�=�K�-�-Y�ZM!�|DDe�y�̄�PGK�7�:HF�\j��=Rf%~�[�0?~�$3]�c��tx2�Cz��v�ռB�!Od�MG~:������W�{����fȬd)9�Q
:[K,�ުu�戴?^���Y)V��5��j���C��>�u[�J>�'u� 4y�����y.2�p0�m�h)��|Sk��qQJm���"�*�{o�8Ng<'��0���E�5����P��/�j��X�Vi�w~)k�l/�A��9u���A�UA�� �ft���QM�{���,�v��f��|K�f���|��P	��R%�#O��X�V~@��̺�-4 ~A�mĔ1�	�g���΀�
4X�H��А& qΣ���F�p�RVeߵ�6_ʖ����^Mn�a�BT��4Q�M�S�4��7hm<���ɟ2��^M�e��*��I�n�����srd��*kT[H�����ѭ�|_D�Y�l��	���涨��#7e��n�JӮ����.�ˌA;�������Y�k��/w��F*DU��)��[�^ҽzc���qड़+M��nj���b;���?_�"�ur�9�˂}sܠF�%���O�aL���.�XZD~�N"��ӹ(F���wU�B�Co�
����~��XN����eW׆xx0_PӼ|xU�Wn I�#ԩֻ��h`�~�������__�"��7I.�p$��Ͱ���_�8�3��-+3��7çeA}�*�=h:�LC���EB�Y1�j�K�M���^L��ND�s��,���J� ��[�B���B��x�{���,L�9�ݿኗ6�*L[N*�S�#�X�a�XnS)��ӓ�|?y¡���$ڒJ�U�#2h�_��\M��)HOoBg��C#�����,�au�#�^/�"Vˌ,*����ܥJI�3@�T_ά�A��|�SϨe��2pu 9w�L�I���SQ&PO�M��3��I�Y�f$[��1��`�bV��Ț��l&��Qr�m��-J����`0�n�J�@�2�f&�[my�i�[���|���B���U=!p��4X�����3;���1EP᎗���Vb�%�����w�E4 �Wa�����N{�E�b��f}�NgO�r'tM�����w��ֆ|/�mbs,d9T�t�8��8�Rw�g�;���c�	[	%�eّ'Z��1w8����R�{� ^.�m�����^K��,M�����6Ѧ�gQ6��L'��K�d����y	��9˒��t�۞�:���>����-U��+��i��|��t��"�I�d���� R/T�gDJ�y	[�_���c���e��uy����,½
�i�8�w��b�$q|G����; w�DF�{b�mgH�C��K�Au<�2T���� ���d��ؕ��l����m,f�@G�7&{z��,W�(fBQ+��]�4_2�/*����.Q��Dni�I1�����Ѹ�r��bc�����O`U$}����U ƴ�M愐oRN?�<�;��}߱�)�Mq�5��i&��?�!����o�������W�7k�6�ϕ~��HS�GqG���C��w'R�M�˸v��3�DS!�7Yca�E���Bw���uT�f4@]�
a�Y�佧���jEp}w��5�Q�� +]���a��Bf��Ҽ��3]�� 1b�#(�S"�##�L��/���TXl��N�	�7���B�&�p�m٥�4`���� k��C�G�W��z����7Ti���-Q8W�*e9�h̩6�J��4�<�?Na{����A��7�bqǥ�(��ת��&3_�,�ߣ�FJ��{^��#�)���z	���t�\&Nq�Ʋ��0����t�ܶ�˖
�ĲQmw����ӫ^��И]���1feS���A���1�Bz�B�������j���٤u,ӳ�����������џ��a�bX��,�j�xH�F��I�L��&6�<�O���qV.N41@���&�ljH��ͭ�E�e�R�«�c�O �ꂢe�߿��#�d�t������%Q򓲟��๖O��x�n�/n�hC�q����K���=GP����]:ǰN��_W��f��ṙ3㍖�x-U"致,��5�������� oi4��1���fOߺBL������?�h����y���"TP��l���X�XL�U ��W�����V@��A�E�c��:��=��L�_`��"�t��B��W�L[}��j�O��(�i�����Z�I7c�yi�����3�,|z�S���.�{�׹��ѝ��Ev��d���=����I�Xz'p�����F_��t�$�d�S�����i����T��}�ԛ�%x<~���}��������x}��o�3�Iǎ6�O�`�>���Jro��1�0�8�������R�D����`�]�6��ɎSŪ�(���Q�%�7�>+��&,�((��MS;HQ3%������Zh�a��x��Г[�AK� ��zS�FK�4����ѯ�u�*�StDޖ�!G=
7�|b�5�-M�h&������YFLh������~�¿P�7����2��vӍ�|i��t9�G4F�o�1�`���|n;�Xy�Dy]7�pD�.u�)�&%�8���s�Bb�3�T/�  أ�\�ϻ����7r�[���Sm�
FzU�ѣ�~�g�	ʔ�*I�9��l���ڶi�n�땚+�9˳�=%��~CeL	�s��﯊�"�
+,f�E��|A�Rl�tTZi�BK��9"
��[�'��[)X�(�V�ݳirE��Y�q����RY���ѝ4l�I���8�%��V|%.�i��5�8+��;��==��A`�i4~�S��
����O�v��)�����.������y�@�ʁ�3܎GD]S�F^&�!is��|�ܦ�.�P���,m�BCF�bo�:���2�ux��U��*�j��Մ҅�eJD��'��7���1�g�ڋ�gj�-�:)��M�NY�؈Bݛ=�}��kw��0uWW!�R�k���2���g��	�bf��L2�����$�q���=,@�~��?���>B�b�o*u�Aս�[?�
�	��E�O�Ӂ��QHV��ǳ�&�6�dOCs��n��sr�ȭG����Z��_W�t1���Aَ��v�����r"�~i�W[�����V	�~�X��C,a�(��-��'&�f~�E[���6qj�z�*���p���������Q��D����&���Y�$�}b�F��W� 5��l\~�)�|���(����餟X��B	
ك.P];On�'ۉ�᭰�A���3��ݽ�g��No�'��ѓ^�9NXH,�;�hf�܆�����{�/�D����#�s^uY�4��W����H4�^�Q h��Y1w"����"d,�)dV��;����4_��lJB���Ѧ���u^�SO�H�����\���=.U����u*bը�ڪ���
���ۜ����V>��[�����Wf��u:2/!>zN���-7�҅�a�ؘQX���Ď�S�o'+���,�nA����+瀾B�Ư����o}}U]� ��J:J���e!��Y #�"�I�MH�6�z�D�n�j ���y!�����9i���|PX���s�<k��jZ�p�d�Ƶ��T(v�/�~�4�N�����4������g�Φ���}N|��]o�06����$�r''�ףN1c^�4� xl��"��� {	��^�{���bX�w6�䦶^÷��aU�{<��ڧ8�8q�<�uV��왇�� 5I{8�C�ݏ/p�M�����W�~�9G���j{V7z9_N��7�5>�K5*�c��C��YҖj