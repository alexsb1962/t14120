��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	������&�RS�����c�I�����`�OiM��ި��-���	�6-�l�n8*�l>A�����+`�CاZbC7��ł?h��6�ņ=*�C"���)m/yk�GM$�V�]�Z��qs1Y7�s.5��D�< ���(��OkO�# �3A�wL��L��M�I�Tҏe�=j���Vֹ��h�־��\n��6�5�왦.8 ��:�H�m��#��E�SE��H�#}��7�*0�2� �����Hj׻T��l"=�=��Q�d��ɨx���mn�����U(�` ���̎�N+��o���yrS2\�i�u����+Q.nU�\i'��oV����NDG��|�To`��~hL�%���hzm��D���E���Vbw^� �G~k�7�}+Jc+q~�W�rJ���;kN�F��=7^b�Wr�)�>��}-��oB���u2MAΦc/O���0���1`�ߟ#��F�>W���o~�_W:GlZ�b^L�.�gv��;���
_�wƲ���JA�o/��ǈ��b"-�/@��f%�t�������s�ֆ�	� Gƺ�0��H�lD�S�p������G� 1��:"����~�92h�����AH�m%x@��b�Ղ�6��Tͧ�~΁@xʿ�3�uz�E�Q��,�ݜf���;r�{z��+5���$�5��^m�/����H´�ꢿE	�����M�6���T?�\`��+?w��v���#M�W@����PVٮ�殣G����l�U��o��G?��N�|w�SŽ�U�}�AɊ�x� B3Vn����0��<�DEi��b��I�.� y�c��KM>9^+���3Q��F.�Gw2���j.�(y�u��J�q�E6�@@NU��p�kH�Q_��ۓ�Iu���㹯��:6鐗.�:����s�>�JCz!UB��$�S&wY��?�&�C�	�na��1����
�Ћ�Dl6���QH�l�q�?Y���P�o״�I�i����E���.��Ҹ�l<�������l�B��^܄E"��1!��.��.����1P��OY�����,�,�՟>ZR�5�����To1�v��I�X@|m�s�V����Xx��?��`㼒M���6k�@d�	�Q$.�}1�ۮj�	����$*P���͜��`�����nNA���E��T�K8�؂}�
-��43#��"kC9��4`Y�"�d�n?��F���k���>���.6]U�iL��}��8�3T�LGN��_.��Ag�d�'�BHS0*��tL.�5��^�*>�JC9�)�k������'R�Bk0��!�Fg5�H����g�aT#���	f{C�U���� ��#@�������ѫ9�v9�H{_��T�r[��׬{��J��)!�5�G�F�i��� .8�$L���"�dMH��1��Z$�[vZȶ�6H� ��S�z���S��·t�r&��,4���2�j�q��8lC`\���5�I�Ȳ��b��M#�@Z%r�a�u��;�����h��j	����d0h={>�JM�1�d6k8��b6%)�/����6��e@� �u�bŰ_KЉ�V3�ǋ!¯Ӆ�����Hm�/ҰQo?�VȦ�o/�Z�ː����lk� F�Zĸ:��9��e7pҀ
��9� "ǣ}���X�Y����O��F���%�D�|V_����v +J��,&x��7��h����>����x�R*��0M�(�%+��O�t���im����`���DDRSa^{�<����Pl�V�^�2	�0��z�4zo�|��S�.�7Ga,��V5Tm��ق���2%�f�ō���Z����]~�t�∻���*8���e�Z�-��p������E ú͝����3�נ6�h]�&,�vG
a`�"|���3�^L0�UU2�&P�7�\�q2�I��1c���B�1�b�]A���z�m�hzx8xт�vy���m�9�n�T7����� 2n�r��O�Z�Ɣ�x��?D�C �֊�8�����>�Ð
`5����zu�u����v�uv�I�s��"m7�ܩ�T�٣�7�u��7��3��s���iB����Z�p{^D�,�N2\ bM��]��(��;l*V����]n���C��/�|Np�!I&L�A��QAm��r�5��bF��o�S"�@	n9j�p��eZs��7�7-��h����6&�thN��6!�s��tòWk�Ά�S�!ni��j���&��1�r�T��'>�� �Y�fQ�x��
u�w��#��gr��͏�7| K�W���)�׽w��l#��p	$8�y�rbĢY�t2ӛ��`����$^9�#�� #�N��/o�zX=>]�5HOL��3˴�%�?���p$ ��b/�:��@��X��YcL�a3�=ZMjg�$>��)���<7���Ob��M�K���&xz���O�"%k"�o���8 ߛ-�8�����aG��>�E�No޵������2_]��^��Ui	 N��J�v}�;`:��ʟ�]�XY!7lY�n8eQŊ���v�YYڀ�F��k$�:p�򧚣�;��T����K�a�6Q��F2�;�:ɼ��ϒo�Y�RhĨ3?6��u�!�W�/���n�g��?�ZI�O4����=��A��@���FI���Y� �3j�
*�g6d@Q,(� a�۝��і���,!|==�h �n����9�&�څ#�&Xa�<�e��4�t�a���$"�h7�$�zϵ�u&�A����#l>u�5���QhL�8.�c��p��z���'���Y>��k;>���-��&4�U:? �R5�Y��$�Wx�ݫ^!�7��玫��O�1�42 ibJ���FHq]����?�o��kCqKK�kX��"?:�7��v/7�ՔR�@������a"��7��܃p��1��N!�l@��A�⭡�����f��ۧ(�h��yS�Y��P�#�ܨ.�Q�{N'�t�����T�/^S�%S]���)�2��ᐵ�$�Xy~ù�˻Hm��Q�~L?���(ߺ��(_�
�s�^����R�}^�R	^�����"�׉�o�nk��I0kCI�U�)��K%���<��> B�]�Dm;�'�����Ks\�*�Y�6�N�nVHa�~���x�����e����^��d�F�T�##%�}ҦN���n����"�R;]x%oR�%Z��h������Q^��/���b��HbK�I�
l�{'� [V�D"tG_~�R�G������Z��&��.i�X~n+u�'�z��ٹ4F�i�A���踸����� d�#~�t��OS5܈��D�	5������Z�GQhZS+��M�B���dk�nl��"L9p7�G�!��D.C�02�1t�7�i�6vzi�bZi���
�����ͦ�>����o��n�[*�u·�ϻM��P�����po<;��{K0y~,{>���,}�,��h��B#5F~�N�Q�6f9��IpA�r g7�eB����/'Edk�4����x��t��mrv�R*��g|�gܣ⮘w�¾��h�^��q���IΆ]���w�nks*����W#��3����������z��;~����C��3k��B�Lʺ�pz�+l��&!ci�ɏlE��Oe�$|�5
�=�q�ffؠ�9�oE1F�̰�n�mʗD5�1��gQ)Ӌ[gs�y'W�N6�M�d~|@Vuaa4�E�y�lPE��.Kdk2fo�a�4�4����t ������6�Ahz�`�0���,P�����=ĸ�`�������Y����'glb����{=�E�S1� #5�L=�5�5UW��(4��d�W�po�-+�)�S^�#M��I�`n�'��H�%���[>|H���K��G.=��˖8]�Sfc�i����m�f�%�H�SA@�ҳa���$G��Ţ.���� OC��a[ܝc�\�f%��������|xd1˼�G2ȿ��~�35ǖ��N�a[�E�H#����,%��	a�>����DL�{�h�[�>JT����K9j�+i���S�1X�?q���Sd���Q�J*��m�\h��*e�4��-�6ɮsF6Ձ��{��mb�'.~�N���@����S_��-�Ik��6>�6���J���{D���"�j4hp8I���Ss�!HQݨ�j�$\��}�Gmq�w���h\]�Nn��t��K��
|��7P��ʱ�R��5MJL#�k���#�4f��/�V-�g_=�	/|�s4�+��s��a�4uX���{�{#��3rl�]��,֕�o���do��ơޜ�t��~L�:��,W�:"�$VU��ʚ98��y����]"sy���T&]N�e%mTx�s�]����Ҽ
fI���5.a���	4 I���ʡr a��b�4����F���lIԼJ�w'�3�>�]��N���lZ���d�`��ͱ�7�V�q6��K ���b1�VH�C��(���&E�y�^|���]]�[sM�d���*?��aR� hW���О;�u8p���G6!O�$x�q�ͬ�*sՁx`��Р4�����G,��_��f,���E��.8�cv!�tץ�)��v��
FCiG�4��GL2��M��VX�a*S�N,����u�t��@�����fW� q��'�����H/�����(?��bֈ�1���϶9Oo
�rv���~�1^J��������7O$�g�.R|Q��ZBxy�a�t��v��U�]�7N�[s�[�xC3<Kĸ{�2��-8@��YPf��hŝ`���}��v�N�^���9��	�ͭE4G�}Nw�,Z}^<0%մ��$>ߖ�s�rP>����-���g�� �wH��j��}~wx��^��F,���E�
��ȓZF��ؔ5��'���4l�*aXժз��wY�R������(=^�VmM�}�ٶ��,��@� �SK$�>��5>�o�ز�~@��,Ǌ����������x�bI�J��"�%�ovȦ����ΑF��ݠ��ҢŬ��
�;�JXt��/�jҭ�u+�8���w7�h"�4�azb�`�^P$l���~���dvlo�r���J�x(���x?��?	 �9�~�/t6ה�D����!�3�k)
,��m�&���:�(�
�c!(�+��;n��:���A�X���Ib'u-�F�	:Iv�n2��I���^[��R�i��c2��NCpIՔ=��U~��VP����ּ1�3L����3���i8��a��#K0�ʷW#��p�d�ϽH�2��'"���׸�r��:��)Ϋ����a7q���(��#&�[t֟#�����u�/ ڝ�q���+��9����5F
!O�m��¹�m�	�e�lc�V4�Q�-bZO��zw��������ڋ5E�k�Nz���a`i���o1�����ף�h��GT	�t���ǲ����X�t��QИ5�eq�)���Ivƞ�Ѐ*�����_Q���`�����y��_(��j���S��7YSf�P�S?S��_Y��#����9Ó��Kb]�ڸ��]�pu�D� �0��6]m�-g���2��X�խ�|�42��k�$����?��E@͸t�����p�&�����Ӏ3����yn�8�m]t:��*iB����t2�?�Yd2��!��G��,�TT˂�Dr��`Gȃ�z�5���~�2�>��G��B��4J@���fPN�f~��;��9!�F�Z ������u�2�3�%җKh�:u0�i8b��R�L� ��Pȭ�ҽ�~�_#�NpФRk0�)J_Q���F�� ��&��'����n�j�p�z�аL0PT[�N?�,9����8�����
�I�N�/FB���9��p����4�]M2_��8�C��L�8�?PӡHπ�<p�qHl3�/$&��4�"=�����/$7�3���G�/˫�a�<w��^Z9��Ox~ �C,h[��)
6��Y��!7�]�0�".{)�������"�E�3)�Jc;��Iٛ��������ez3�VBИrD�7�%��nQ��?�BEK��a�t�
0���׏U���龂��anoD~�e�N��)z,��F�z'�H�.�6��%�ɜ��ډ��C�f.������d�"�����,��^*�.��a?�w��\��U[��Jc��dÌ��[!�[����"<�c���:��;�X���Q�?�ZT�z��N�(}��S�g0HRkщ��� d�5��^��re�����?uP!��Q��QM���-v]����V�{�"۶x�H<�[v��[�6�:�'$�]N�n�;'~��~�4��0��!�Q��G7on`,�7Y eD�����,Ļ!���Tf�˒I'�4����v!vN�z�^�zPa����]���e��"d��Ǭ ���N>'0��S櫎<Y�M��R���3����Mu�k';�P4����>U�=hF����Y��aB*oo'�?%xqP�d%��	G_��&�<�Y��4*))��p���
������i���U{آ����	�?X_���$n�v2�����,5OY�s��e|����vB�Ι�����!5�Q��>O"mB��\�N���p�h�'���)v�@�5�n��@���φ�r܆)�c��9I�"��E�SF��A��7j-���.�s��{t@ސ^u%�//7��`5���(��EMY��cy��G��,aq�I�_92�����Rp���I	8�by9�׍���W��â�~hY�0���D��t)n�W�?w�CG_s9���1�̻S8�K��.
�5(�c2���l˄#l ���nJ��|9�w�Q�p����n9I��A�9�'c��gz���-W�#Z>|����Hf���.vMu��wT����?���OB%�8"q�G��&���C�X#����u�i]�9�8��
$_�<Y����,b������v���л��{	;�)��������[��_���55ti 7�G��ӫ�>�b�'�c20��0�w��]���:\.d[#��4�i�Z�����4Μ��rT�Ȋ)ʞ9������Vc�Tg�v 	����j*9�� }j厛���%T!��+&�� �/��V{b��m�����jc~���7���s��16�C�S�q
���� 1�%�\qe�F�S��D*��%�4��0p�Y��8d�7�%��`�w�g%6��$B��q��PL�t|��+�{|@�3;}\�� �~O�k�O
�E?�O)I3o�>w(��:�OX�%f�$�q���8���=���������9王4���t�C�e�ST�ܚ��1k��*��JI��-��K�wm@�2����yq&�B�����n��0��\����9�Y�d��>`x��x���Q�4�-����)M�O��)}�D��Fo )�KC�6����v�/p�|˖����
�}"f �0��Na��M�e�+�C�ۓ��SCOB�T�|���j饩<���\_N�AǧF3�I,5i�@�Y��	jL� 6S���6��A;
xVdI_���u��=�C���GK4@q�F��.+�q�7$-���q��g�m�u#2c#�C;"���r��(L1Q���m����-��柁Txu������3�YQ���Y^����?
>� c�#�ѿ`r�藙]��Z�mv #�$�-����5�W;�/5�e�(�|dYh��S������D�j���J�E� ����_�+��Mql�X�_-Wy���#N��)�@�Y�"Ѯ�4Ҭ|��5VvV�8���(K,���S��SKw�&^옏7��Q_8�C�7�vd\����-�?��mF��(D��bG+�ő�^������脖�*�s񏩹�6���I���I\M;�6���1{'9�6Vz]X6��)����q����[�ApKa�����'�"PR�9�./g��c��4.Ce�ȇ׎S။��Uc1���Qk���m�KO��{�I@�a��-Scg�&��]������o��Eh��2 ���R���u۫��AxFM��y�3Ul�|��NP�Nk��hK���Վ�U�b8;6�����C�����'I{;�{ �Vx���m�ߜ`�ٸ9�$'�R���З#>r�`�F�qe! `�wϴ� w�eة��)���T���?���2 ����� i;�pM��u�Ct�j�m��hEnI^~�&%��z�$�l�.f���հ�o�P���l䇮kΓ�����]�nR�Ŏ$�3�"4�P�'���]�/Osz�9\��0�[�� �"�=.��nPi����������vМ�ڭ5�G��(	s�8�����֊ b�{
y��	��c������I�$�<[t9���ޭ)q]�O��˷ad���$'��{��UM���y, -Vẵ�������$��O��Z�Z�U�F��EѦ�
+��	��ʿ�f8?���2�[lqO�����?�_��l��2$$I��˽�+�m�M;�za�Jd�c�w���O�)"پ�듥ñ����"Oɍ����&�;-^����?3�
3��0A+�?U�1�IY#��G\,PQ~j�fi.mP����]����C��Z�o���SҲ!�hS�6t�9E�c%cD��ߩ<
#\`������4T��b{C)W�IW��ʡ�-��,f��U]¾�{�(5޼Er��BI 5R6#���Dg��ԙ��fu�u��~j-9yx�QkՇ���ν�� V��ʮc�0��ݢE��A��E�?a���k+�t�:gH��y����/�d����Xnorf,
�K��>�mR^4��~ΰnnGJ�}I�}(�����35	�}��HE�'B��3�]x�JҜ�p,c3�+�B�Y������R������oAq��MݹPD뤹T�"O��.YA5yT�Î�"~��Y�ͣ��ϖ�_)K�xG}�3~rs2���˔��$������C$#b�C��(��^�ѩ/2T�@t�X��F�����=2�Ǳlx7��,���̖�w-�6}�;��������
�ݐfzq��|��f&����'��A���w�~ƅ��j�xr�J�ɮY��lYMgk��� ϗ(�Q��WF��sF��`�0,ʠQm�)�㖄Izk@o�_���]r�s$g,缶4@Y`d�,�A� �B��F"/��)դ�ݻk��l�_�� #$L�`o����渪�i�Zqr��HU9x�@B4����6(�ώ����:<١������t3ܪ�CO�.���VkH#�>;�F)F�
�܁2��-����e����|��b���	�8�v�L1�̐o.�I񹕅�^�K��]R_a�����S�yE>w"7�m�Q�1|�AN%9�3�ejV��|k����~���os(Ew)nκ�,d�H��$	���|�!);L���e���Qn7<g{�:���HGJ�Y���6/e����@gJ�S�����n)ʚ�]���p�Ï�������T���E4v�g@*��rUr�WB,1��k�2�_���ǏQ��m/��1�d�b�f���WF�͑"Z�r�ֻ V䈲p��,8�l����p:Ps�nt��J���-�Ig����󟎨9璁��ʫ�U���j7e6��ƹg٪���y�7�ʊp[E�Ǥ԰;�S���� �#�t��h�ꈫ�d��%~�����?�����mr��u�y4H��^0�'�����|���\,��ZF2�6_(Cw�}]k��Q�j��j|{s(OWz��RY�pP���C���������J�"�w�3$�+��l7��.�}���%>-VY�O�R�\B�iٝҨ H��%���	��Cׄ�Q��k-��f�pfDu��A�p^+����; u��a�f���w3>�������E��~K�LQ��m�GN�������}Jx�
hM�IL�{$+9�t����{$W�:V���΁��HW�Yi�ř�K����e�f�-?ɯ�G�`�JA�O��P��E��9����l�$��[0H� 0����e��Ȩʌƣ"��bB�,Fpo�;7����ܽ\����73WΧ�34 a3lQ��Ҽ�u��~Z_�Ϙ��`Y��մG<��U��	��'pE~��4K���v��}J�q�%��S�vq-�Գ�m�)�	�􄥂��\:���O������9|$����̫���/Nx����+�/8���I4Vb�k<1��O)�����jx��2w���샵�F�/t���)<Bm��˷]�
S㙙�,!Z}#h�"�G����|��)�k�ǿ��%F�lD�>�_���B\=a%S\pr�_��%5G������0�q2IuD`�
���g>u�IX�S*fN �o�1e]��f���bYgY�K�;�<k&V�1M��c>u��Knt�$�VЅ�w�iג_�������O�_��<�ˡ[����$e�c�@�	/�]�O:�[����^��!�0��_�q��,��
��o>sI���an��Ѽ5�͠���6�ze�cL�f_;�H�_�\�8��^da�x����XC�!$�I��w'?�I�1}k�gu{A'����;��q��:�v�@uL�^:F.���P��vX4r���"A5�m{�PdC#����BO�d�:^��NU���6	��s�7��]U���L������ J,`\Wa�)\�b���i3��9�&��_�i�	N^��HGi��`�i�qjֱ���|��]��1z-B���m��@zc�U��LH ��;�8���5��ʮpȱO���EЀ�
��휀P�+�ֈ�9�`�L�(� ��4��ٰ��ؔ/���w�6�����۾Tzh��-��[���ݷ[Dm��J}�W<eՎ�mV��aU�Fx4"iȰҖn�&7�ފ�Y�ܯz����/ޟ�n���ۓo3��daP�������5��}�Z�ܿ�p������Sǂ�%a��(|F7��V�L�:�g��K|
�һmwlO'q
&E���N�%n�\n k�������@xv�I���I�fVU�O��&���6�M ���l�_��a������Cd���}L�u'N�*�C4�Te���m���h\������#@?��u��Os�c^h�8��5�D/����R�D;O�4���/���{��gӔb��Z�A,�Pl~�n(SF�`���Wj�������� Q�*���d01-�7����U���W���j�AL��ӛKE��,R��.Б4֟o�8,��ШHI_�e'�Q���cTgmu{�S>h`|E���+t\��ڕ��C�8Ø�/�;�P���/@7hH����뢂�� ���fS!�}Qz=cI�ZoĲ��Q�bR`!A'M�ܹ�O�1Y[R�͹^�,�M����\;�V)����,� V26���h�|���q^a<ɯT�=��"�^�fT9�9Ȯn������$1`�uMP�<����iD����?�
�V�a�2�չ9T1&F
��Nl����S���]��JҺJ��/�툵�����/w����ZByH�:��		�K�|�Y�?���#�c��IK�*��N��Wb�\���3��IH�t>�5�b�W���:I=���ݺ���	 ��r6%�;�2���46��&��oNC_�"˽�{�j�>.p�͢(Ĩc�G�^Ww����1�*�$���f�[�-w>=����)\��*��7�&e8�[��U��O��N�*��v�I����*���C�*�gD�Ľ-�c�ŷ����pJ���Q��/)W�|�ϼ�>Oc��)�eۿ�5�B�iȝ1�|�H�*aWx
(�`*��b���ESO�@Y�w_A���d��G��t�8I�P��i)�E����"�SX$�� ���	�;A\q� ��ck�+VƋk�f�>��ޑ�N1Z��,F��X�Q�י���]]�2��o����z�ͫ�������c�-!�.Ɔ3F��E$Sb�?�Dc3�ۄ�]�6N��B�r6�]1vGh*ą��d�U�*������i@0�s� �0c��4��Í8+光&�Y�.S>m�\�{��� h���>���c4�Sx�ն�Rn�O��'�Ѓ�9�ٚtV4�m����Q�V�����4Y Ї�u�&v�0ue��?#�7p���c�=�_��bS,��H6�� y���o �7�.%m�3�3��7h#s�9Ck�5�,V^>�p�_H��kt�K)++�fֲ婦MKq��?S3LA_�5�����ǳX�2�5���D�Y" �	Y+Ֆp�y"u�ǹ[f�@rMKpkǿ�̾�����U�8u�k�O�ɝ2o:6Х��r���g=tSv{�7��*���B_��[�!��i��u&�����Z��Jhُ#T�����.p��[�ᚍ$G�l�h����7ր]a��5yI�@�̭1D�N���� y�O^�����tǛ�;n��!@���[���K6!x3>�ƶ#�Db8J��2��;^E]��0�G�rx �Ѿ^�=�'�B�`J�\�_�����r�2���DX�Fo_��@��)��0���⎖��R�L^Fw	z!vm�����ș�Hx�OQ#C�<"��s$�.����=^C�Ow* h��x�~��%)v��f��󵘄�\��]N�;uC�y
�2n�x�Q�jg3�dE3ԭ�b��P"�"6}IX��wg��r�c�|>N�~ߵ��+[@k@��'�bv�0�;��}l#
O�,O�GZ�+���d1���Ძl��㵶 ũ�[2�-1]�p�*e$���մ�[/�����~�&�K�0�Cݾ�u*���-${�����E2S�xB�թgg4�W3UE��fBJM�c����	h�H"q]
7vJ��?"��_u��)q�Z�iP��<`��͟�3�N<2�[?-S-�I����{9�u�L�pd�g����ǘ���Z��KǢ$}ՙa�џ��DD�ߋ�`��4Jp�T����V���N�������O_�N���'��I���d�7���eɧ�?~	>wS�z&k��\Sbu���G3�H�{s�D��D��Je�͢�D�:�4������ը�5�k������/I�/�W���!'vH�f҉=�sw��݈�I�h�x�T�Cvm�g ����Ap�Z�\����1� ��Ofė]�(��
�S0{b&*gG!��ګ��7�~�G��cH�
�����R��.�m��n�R���Iwjw���׎B�Ru�`�b�)c�aP�E�W�$�-���;V?�<�	F���-�U��A��8��d���&i�)P���7n�?[�#�k�$;_�`�o�$���`7�qIW1�A��t}�����Q���
����#���{F����b)_�n�e,��d���U��j(���n�`4�.�u:�����>/`��3��[� �lϧ$,MQ�s<���
���A��ͯ2GH/`ۄG��r��������J�ڊǰ�YA��Q��CUS����by���'�>�+`zɈ�dO��G�jj�B���oW���H.۝e+��Y3ʜӷg�B�=������ǆ#bNB�x>��Sݮ�4��CE��,�m�	ё?o�*�E@���_2�b����e�Jj��#��o��MNL��u0��ÓR�}�.��^���"m�C@��}�;� �fo���a	����>�z�N2lW��<�>a�PqGx�K-A,��}6����n:Y�m��xv��(i�Z]D�y��*Zlv.z�X.�M2ܞ��k\Xb��j00��Vc*`�s��S�B-y/��̠��.�O v(�͡p��i����0^nU�Xa��W�nL��p!j+f���m}Տ��v<�b��0�16JZ��j�H�c����\��� 6��Q"g�� K�j�ݡ�*x�:K�~�PY�W䍿}ʺ�q���cʺ)�&�iS�s5l�p����:��߁��^u��d���s�L���L�_�+hzW� ��%���n�ȣ螠X���ܐ\�V�J��U�եX3�խ�!��<����X-F����������	�N����<�S�^Ӌ`��~t'�*J�髮\��\��z�I�!Y�ׄ�����*/�����8�НeH�ʸ��<�n#�i�z�0��?����JQ-�^�ū8��0�1��)16Ű5��Wg����:7�*7����#~L/�Lܖ�!���� ؾ���,!JA�q#2�Y&V%��k�����X�3�H���W���8>GZ�!u]�G���g��P:�b�BV�0T�8]J	�IZj�z���_�U]����y��z�H�,����|�t����i�lt�,�Б����g���D�=��}%/ѭ����n�V�t��g����я������6?��m��Si��7*x�|�y�,p�A_TJN�;-�bL���
VV�^��S���8���x�/�
c�^ENh�9���j�ϳ���BC8 ���I�Θ����R�{��&X�2�]t
�Gb~�����@a�U���K���������jִC��#��q���ղު�أ�|#�xU�f��ս���:�7��� b2�X}ń�SZ�5d�~�����Ͽ
}4�|��ٿ!n1��̘��P.>�%��KJ/����]6�S�~��_�2[��X��8����W,��o���Xü�7(�o��[+[򿽅�}�6tXe���6L �k�w|ց>����?d������{d��FNZ���k���T����@/\�|��	���)"v�̤i����KGj�9�nF��m�a�i��Q`�+t�Oj$y� �kYl��`yH���X��U-�����bz��E�y�
ш�Y�bì��o<-50t�N���Y��R�O�WOi���[l��(�ؑ���ck�7����m)&2�_�mӲL��G�D<e�C]#k"6����\^j���9������+���Ava.	&�Zx4i������.?�Z���\��#qB���Ɣ����J��
S6Bk;H�"�Ќ���nV���|>���M���u��3�w�&�c *#��cGe� C�{�7ø�� "7l�P�IEPB���V:?��M���<t�gGI�9\e���ht��A��Rg���+�7�T�њF7��a���������R�9l�S|Ѽ����z+n�[�?{x{D{�Zѧ��\���J���j�y��z}�m6�л||��5/�J$� A[�gz���6��W:�B,��R[�T��y�D��Uh��
�i��u�������{�[�ͺ9ڋ�".4{y�I��j�|�)�v4ev�c#�8�*W�+�e1�xD��2�(�F��%&��
�lӫ���h�S��B�ժS/��%��k�%i��WBݩS�F�_�D�N�;�������[��:��lz�i�pd$O$��C�|�c"�ᅣK��%���qz"��6�Uok4������������N�ç�����Z��qL��d��lH��x�/^�"}q� ��~�Z�@�Z�S6���54��
�6����N��lI�_�h�����:��8�J�:�Pt6Z{wFsW�X�5`��"!q{��A�K9dl���'�L03�8�v$��	���l�J	־��h�O^Ϋ�bY��}�O3������R��WS(bs ��~��������,�"+��3��f��V7j�M���ZI\�.*R���ey=�W���d�^��5h]}^K����_� �7�ݗD�p����t��^�>�b�rK�S������w>D���e�����*���k�Vǣ�L ���eB�K�nC��@�o�n�f����������z�Wf�I�'����f�'���f�wv/�}���#:k��S�Ģ����0�I�h�d,ȳ2��|N�<�_`���&�;�
��6��l5dr���iot:�N)���?1Cʸǖ�z�\g���@�E����d��
����M=�$MR�\�A瞒⯔�]O[��7�݆�����=}_kA!j!�z�O0̉o˿�sL��T�( .z�6��+,5�z�b<�j ,�N¨G~J�Ս� 2�\&V�u�m�*�G������}�&�+'�{v��>o���t�Co���Ac?hl����L���O-_�9����7��Q��a������,<9Ff����{���B� sq/D7�V�,�R��^��yę��d��������6X��G�t�u?P�8[��	������������w�� b;��ᚡ�2N��tY�������-���vܤ't�U���}�IV["o��Z�H�F�����)�_X���o�i"ҡ��:.���m�⟜vd8�$�e�8|/@8�%�^��6t���Y!b��\�Ƒ#,��$ɲ��Ɂ��U&�Ķ��Nś�谇����?5�YL��-�a��E���HǏ-�+Y	v򂫮��G�ۃy��aXb�b9�w�蜥�@ǈPZam���˰`�+����������s�~k罀��߳..k�Z�/��\�pgH0{� ԏ<�!h����FG���;���������M��%�őf�̴��b�J���b��?\���l3���r���X����&(�<ɚê��n�$	���PCq�z�E���r'~W�y�ZĶJ\�%O-Z��M�2R�n����G��P�9���G&_�O��K�
�`*����"y1�ٸ*^\��hڋ����\��˺���tKC�6D�̕#���n���q%"\t�`�|Q���9�_ٽ�����8�R_�<3���7VH��YT�D^������]��DJY���=k,Pc�L�OD%�
������f��nr��N��ԑ	5���t���\��/��b�0�+���6��X]�p��qD����
w��́�u%�U:#��%2��8<;�O]
6����*�m���}�wU�Hj4|����cP���4��a��VG1�a����~A��{-����q#w0�<�V�όS�����fժ��~��Ɏ�s���)���lPv��7ڄ�Z�Vǋ�:ކʜ����z�eU�e�҂T	�l>RQ��g�t�7Kb_ �aEGW���}���z}�I��#v��C3֩I���2>�g� ��l���s�!xF,�²�G�-	����D)P#S�� �>����~Kn qzI�eč+���b{�:�G���/��h`{ė��n<f��0 ģ�V���-TQ�_؈�&�$��(l@��A��x�f�`�5��W���]R�����R���#��h����4����{"Z����eF�\I�N�|�i�/��:��� ���jM���dS��2D���Y8���(�+W��/���mT*�0���~��K�C徴�:�a��ܒ ��]���~/�ֲ��ޞ��}�\�3��6Bbm�4ѭ��Fڈ!Flo�2��ݧ����%�R�T�C��=�S���-�(�����&���� Z�j��$}1������֩~F!���*��p�=~H8$�^\uL�@�����2o $�_��ƥov�aΑ��r�f��FS���	,�#:Rz��ʏ��'��@N��!��&�$����c�>b��ɩ��2��f>�x��ɪvdn��PP����O��1�u��U��֪g���Z>�X�� ���Z?%@1ꧦ�E���,t���Mu�z/����)-��)+1m6�F��W���[�;�[D�v<��f��!Eε ;�~ܾ!��1�L�$��\z��{*�e6�\�|�Z��9��雕��%[�A�f�a�tF��i����v��yx*e�UҜ2�D�S����-�Q9��x�	���3!�|T8�*b���C�V�;���*(6r��a�a|���FJ=��M:���t��?�xW\���x?�<�]�M��̠����#$$���.V�N�� �6�����ܺ�b�,����u�å������3�N���d�G].�q���6����nH4�ڳ� \�=$ʍ�q�\Eqk��y�c��0cQjK@�2ӯ)qуGgOx���SlH.4�:��ذw;�W��T[%Lkԣn����/ְ��NS:x�h����C�n^Ht~c~�$w��4�sh_�yYp7�nS�W�h��-] %��^�߫R�Q��v���B����V��Yyǵ�m�F��w�O�p#Oݨn2O�B��iBϨ�2��3u$ZW�ås3���e2IL��!������л]JJ���nG8K~8]\Y��x��Lb@5}�����莅9rIL�S*�.�:���P�K�ɹ����8��)wx1>�`���uL�K!��m���	wm�3=]Ԝd��𜒼��N���B�Xz8�s��zT�>8�߱k�'3���}��xA����1U<F�s��
o[+�&F�}�Ɯb�j����ȣ���E�Bŋ�l򱎖$����p���:��+����j��	[�����0F/0����q.4Do�Y��2�l��RF

.�R��J,u)�	d�?*D�
5���e�G���]?K	�MaU�^ڤ�~5lx��D=�y��w����t���P�|��]��>��^�S��($���rL_���G R	��A� b2��C��0�viPEn��	�=Ke��H�с3e�_Y=�ҧ�o�[�BP6| ۵9��[� dQ�n�w.dAԧ˘,yW�����N'�l��5-T��b�,	@y����>��m���])	��������eh��˗����gK��].�8�-��He�I I�׈=Sɉ֋Dn��L;�����{�4<}([�C�QG)w�}�'����3��ԁ�L��Y&��@�V#����a;W����+^(¼�M��mSf�};݊	�Py�;3��P6��q��!����Ĉ��:4ُ��D$����O�ŨvŢa�@O>�t~%��(��:G]�4|w`�����"�" )���nFc�/$�f��6rw�D�x�א���!�?^5ZZaI�2�N���R~%�p�ɨ��8��+X_�;��_׶msf6ɥ3�NJ��͑K�f�I��B+����J�����NH��B'L������f6���c��a�_!�E�Ma��+��Z��m���r�I��U���
�^��s&\ű�������T�M�$�Fˣ���L�j\ճ޸��S�}��er�X̈����'�Y1^���½V��H&|D�_1�?@���<Pdg� �� � d���ډ��K18<�dx
���^��jΦ�0X��$���*v�=�Vu�L9���*1t��EP��:�1@�">�{k�u�9w�*sJ�6��¼�0���a�&��)Z0���)3���O����T͑��[���eŕ�]�LaN�hw9�nG���L�`�I9�?�hk��S���m�Q{��t��dm�ˊ�i>\�y<�S�ֳ�7�ϝ��x��g|jM�4�q-H&�O_22�R�1+���<��@��L2P׏JF����n���O��^���W�)P�%u�LBE�9��������j���4Ę�i�� �Qw�DWɵ���P��A7{��{/밇uN������G�mi�\}�p�]�~��b9�RD�B��':�9e��1W��|�e��.��
k�-v�{�e��|Pi
j��(SOc�5�{�T����#h��ml�?�a-���������s/�� B��Ed �!"H��Gl��}���bF胓H�Kr�Diu��
�	��<��b\-�,�4
>	 ^����R˷����e(R�	#��-?gߪ	=��]S����r�!m-��%�5/��)ۅds��R�eZXݝ���ۈ��;{�	���R �D�Zڑ{6�\$�*b�E+�l����T�e�{Xvu[��u|�R6�s�x�Y�L����9�0���{�
mg��(T�G�$u*<c�?Mx�FW2f�j��bK�P[�n	5#-N�t���`���0�؊�j�;^��ZR�$�g���Kc���0&gBp)��V�2kQ���"�9h=���
���$S�&N����[��t@�����I�.�i��H�)d��!���n����GK?�!`K�[P-��PoH�"ƴ͕�ΨZ�#>y���}�G7�d.��9���4�����?���I���J�˯'�nTRw���Gx���H�x^d�s�]'���!Q=����E�֥�b���/�Nd
4�Q�{����U(�x:7Q��>��R)ѽ�S]�~�}TrT�Qx��f<�����W4L��n5�wo��m���������3`;i��e�0rBq�/G����kN%\Y≾�ʸ8)�Yj��3rR�p~
�}�a9,���Pǵ����a�|�N��]g~�<��vcBɎ�ђS���58X�xoFe�yA��{�
��*���-p�+fٽ�e�I�J͔ȴ� ���˞UMA_��7���W������|��=#J���l�?n@n�9����Q4V�Q�ea �u�/�Z�f���"1���༮�հBG��Y	��5z�ǰ<h���s+O���f)�@񮂳Q�~�u�`=*��T���TQ+ⵡ`Ҫ���ǎvK'F˜Cr��u��� 쀆�c�V��3���c@�����^���>�W�2��b�G]�#�d�P`B� ��������Z�x��L�j"�-�n =�`�q�"Q�h�Y
��~҅��D6�#�f~��Tb!%7��"U/Tb�m��xQ�v93�O�:���a��ݶ�t��6xw�c��
�5O/!@�Ġ�����uT+B�p1l���库%����6k*4�(2��Nu6����k�D���-B�נbN�9�/�~�!����[��z�|J��v«G�f�b�	R�A𪞳k@L�^_���@�Z>��Zo�HʺH�c5��7tg90���`X��+�_�%TFq$m�w<Cmg�i�`*��tîn_��>���e�d�KW����:Nm�-���*�p�!�������֗��}��nï�X�jPڃ}�z����9��7͂s�E@��ߊ�)=I�Bi33��GD�U�lυ�z���e����x\
���n�V���,A1S3���1uxfHl��n��|�~$�����l�3�zF�$o�`y��]�wz_?��&]>Q�(��L�����.��U����n�3�WcG�rɽ&��4wx���W�>����&D��� M�@B�0�'=�Qۚ�tJdZ-87����I0M"�$9��	���X�����Y�� a-b�3�N�U�$y�u��q5��ƧcY��Dǜ]�3e�2�Ŏ���\p�F)y�ޮ�$HK����'�R&6�:l���W4զb P<�����l}�>�Jz�ƿ���=D��eA���f��?F�Ni
mR�����L�B���vKx��F�%��s��X�I���~7�7(��7G�?�.��
D>�)�NnRms�QY	�T���gʷ�~a�W�\��Jf���(Ͷ��+�<��=3 �C6 n�#�q"|�]�^�֐u�ʵ�yRS�Qʳ2����Fc[9!lRV>��h��gȘ���T[� m�uM�������5�c�RQ�:.�}@8��
Y0i��N69�d]9���v�i��;)�ݐ2��C����� ��"��"��8JK�&�!5�T�7]�P<ɥF��
��@��p�f�4hɠ�F^Qh �UZ	$��D�qrf
x� �s�5�*{�����{Ҷ`�O��'3�~m�r�������7�� �z��Z���@w$@J�[w�)B�L��5������x��ѽV�~��@��I��_o����Xw�7��Gc�-�s�Ca�3�"�x4�}<�"H��$_��ڨP�:��#	zЄ"��/�z��E�f�pt��R!�Y��Bx_:ZW�[7�9DЎ5JKA�8��U�����B��U���`L��l�lrkr�:��G��T+�k�j6���D+���Ό7�+�N�n_E[��.ˡ=
���JX]�� w�)�Q9�C�O?ƍ�jU��Za��L�P4e��sW<0Uݶ�5]M�n��N�঻Ԃ'��&�+}UR�	��%�|�CV��姵ԊR��ȕ��۽�2{h�=�~���TY�����j�d#8;���?�l%s��S�7vذn��$�R������N�ؾ���0"Cs�c�c�_$7k5��2ˊ�J�q�S#��;x�?�v�]�D�W����� N��qb���>�jo��+Ru�3v� .��1�#@c�\?���#j[��6Q�~��c��k�@@�&E����'S�ݔ��L�1]�[?��O܈m�����;�鵫2��������7x��p�v��J�����u�0�P{i�  h��4X��U鮜��L�gg�<__d "<���<�<��X;^P�g�^<�v��<���߲OHJ=(��;�Nɦb���+p��A��k ���)뗖��4T*>�Ķ�����//�cdG�P:G�c�~^*�����XhK>��"^����k��$�G�
�\�Q<毃k��ֶ�D����7�̀�@����˺�z���$���ɽ�i'��]�s�)8���-Y���� FG��m���śCP��|,�)��'tB'h�����	��q�*�JJI0|��m�����g�����x��N9�J��l~`��:�[������j0���إ'�Ԋ5����-,��aX�f�@O�ֹs�.����Dz�å�b�2|�0A�<��E�&�9�t[�"$=n���+�!��5�z�k���y�;+��Ў|��mS$��G5�����MR�nu�F�6V��#�ýs$��Z)���3-`�D�)E�W<�
#I�U�rOel��:�Q�%f*��ӇW�0�{�0x���� ����W#��|+;�tpXd%MI���F1pY~>����ʞ?��;�667s|������\��%iI�0Dڊ?Da��3l�D���R ����XL�߯�J��N�5�	��@uVy .�z��O�+���*�jM�_`D�$� ݑ��H|򶬏M�����a�1c"����W���e�dBp�����'�H���s�;A:|�m**�M,�Y4�:�y���+��@I_D�_�}@̓�u�{�<��e�?��Kf��������dM��؃��IӬ5�$�Ph���EW�j8��E���|��N5�>-��(�읢v��EL"* q��:oB&�]��>(��π)�Oj=>Ƒ�A�A�p^���h}��2qfCp'����4�P�t��jC����qP��2�(8�<$޹Ÿ�8��,vyv���8Z6oy�C�i¨B�c9��c�0E!�r�ŷ���_}�#�-�E�)���_l�&k�vgG^���9��aQ?,�Ӷ���8�|�,����	�����*��݌���)u
"��s�K���٤�ڃ]K���i$��B>$�ꂋp��fD�LL��rTOo) ZG(�@��_����T�Z�%f^����-&<�%�Kd��>rHLj~��a����Ƽ�LQ�
:k�}q�������%���8q��H��᐀L$tl��Y�(x�����S��3�l[�@΂�啐��ԑn��� �w��x��=�J%�]�c���a�C��r\;���Zy%z��*���h^g��p��o A)p�f*�	}�J��If�u,����U����jY���"W����$4�'��Mr}��6;��"�W/:�&.a����5)�������7݌�rv��AM�ƌ���N��"06�vi����灒����yȥ������'!�j�T�q�7#��1����*Tsf��m��������3�ӊ-���,`|��v~��P#�0k#���;v�x�l�-u��ڙ��4�����$�HФA���9�5���mwO�������������1d�]�z�On��w/��,Q޺�Z�Fx��������Aa�t�m�}����\Ӭ��ny��FAˬ}�J�����B�r?܎�l��_��fa�Ϟ�����Ƥ���-aN��7��z̷ƦF�SD�A�?4�BU���P�����oF��\�v���:��x�B6�B�9-����c�R�%|�@l�f6��4BƼ(�Z��{=A�o(_ceE�O5���8���P�;���*����ġ��	*8�/��)��k7��]j7���%�'�\(V0�7�"o_���-M��;���3������!��s:JNv�*��k%��禖�^/�������B��^I�f�m�s�M���<�(F\���K�r�Q5jkW7D��ݡ-�� {�Q'���x�V-{R�0<V3q}g�H+�3C�~p�vH�����Kz1z���!�����}8y $�Ȭ�}����a�/��Hq#w��n�#�h�F{2��gY�(��D�J�;<�ᔭ��:�5}�F�gs]����]F�LJ)�"H��{��I�۟~0�l*mp�R�1��i'�φ3�#�����2K�����ڟ0jE�߹�j%��e�����{.K��M���i3�D���ŗ�£$A��U�	��($hIB������B�]~�$	3����Km.pX�{2I秉����N�9�!�k}w�����S��E�C�2�ôp�Ŧ���vռ��g����3�%���jR�H��@$��.��D��9��T��E��q!�x4�/@�v�H���-�5,���'im������>�$�轝��QVA�U�t0�;���ia=�����ΪtE�Q���";$�M� ��a�G�������Fޥ�f��ˎ��(ţ^��}�#�������J�U��d?�|�g����N����Zc��ÂW*�L�Z�m�x(R�wp���.��+C.Ҏ�%q�:�� ��V��Z�L�т`�ºP��M���&p ��D܁bU�ǁ�(�ʩ��i�����Pߌ�ˮ�?�u�	�W�b� ��#^*l<���/�����<�*H�!
B� �Fe�(~+�w\��Zc��hS�rf��c�����"b���StN�d�l+�����j� v�Z/�t���2�$�E�W8Zh�߷#ZB�H����'���"G��'c�@��1ا�k޷��ɴi"}|�.���۾ 7��0�7�g/@���$� ��B���a(���Aw��8�/8��w2��G�h*/�UǧN��}����v0?�ңֶ;�.�����9l��ȳ����"X�.{������A{�XjfO���W�S���\�AQ�n�T�>��R�ޏkw�u��iY�uq_��:�#r�����'~�h���X ��2�y$י��L�{��$�(z�/
\z��k�յ�@�����7��H��i}I�K~Ҏ�&\w�-�B�7Y�2���2��)������]x�O�]�l~P�	������������I�^����Qv�KM�<b^�'�W����������-݀�s�=C�D�{������|�ԈE���i(�z��>�xWd�}׈�k	�o6(�(���T�f�LW��]V��Q��E�|&��/3~V�^�X�ΰE�@��e>��z�l�����d1	p��+R���?^y$��X`�,�ƞs���R��v}���zVqM�.-Z�Ӡ |�1PFz�udH_+_̔��z~�)�x+��jR������Бl��'7EeC�����r�h�U3�l���	ґf#=��I��a�T��&�����ɖ���ќ����	���Klh�δ�K���$N��70��^7�{��	b`Jƞ%\r�8U�1�93)���cx�� ��>d�A��^�t���s2��x��
�L����l���y�~��H��� t)Ƚ���?���7�M�-y������f^�Ц��[o����ucL{���^(D��6IB�F=�!u�˵i�~베�U�_��Jl~F$9��� 麌�^�q�P^Í�?�K���`���.C4��v�z�[[����ꃸO �R���?f�_u��G=t|y#�B_��73���p����O �\l������{��O|�q,wב�/���c��o�|SS�j�a���jo}��R$[%�h0T�[0�,/yg>����~�˂�ݴ��0��l�%�R�U=$d��Ne���g���4�'&!�O��5�p&t��c>�u��h��C����	g��Q�q]��a���/ȃ�d�ʡF��7�?f����-������>H��v/�h�@Ăw�|M�N��B�*���Q��c���*�W��rX�΀n����OP�2�������ѐ?��Z<��1�,:e7W��MD#����kRB�v��X� U��v&z܃����ͣ�'L�������0�.;��0�uSMb�̪�/��*FXF�"�<Tz��n
�{�O�BQ�c�Ll���O��XC[p{�A���t�ra���:����>�Y�[9��֡��<j<���F���mIr�Y��#��{�<Q.'��~_<��l���A���
	�,h^ͪV#ʃȰ���L�$Y�z��	�)�c�&��%�q>�2CY��J.�>�Ơ��e�_�U���m��TA�HNR����s��������S^D���c]�����ݨ��a�d|�aq��+�3;��|}a����o,�]��{��M��d��Z�~�j�ĳu`�-p�j1*b?���:Q��%��k*�܎"R�5Ʈ�@:L�ӂ:� �vN�ןs�7�5e<��L�FQ�;�l_������CqK��:+zr���{�e���)��ƽ#�]x����}��aȬAM����P��!`�mok���G"j���	j�~b.�\������T&�Nv��o��{����`���2�d���2g:� ���CI|�A5l����}���x:�E��v�F��)���|'b�M��n9ܓ�V֊;QX�(`#]R�o_W:S�O����W�sV��'t�7OpV�^w ����
oR?jd��2�=�L)o��\f�X���	i�e�0酈�N(��;����N'��!�� ,�6��L_�.U��^�����1�cw@VP� X�PdP�IJ�Ӎnug��[)�����LN�hI���0W����p����[t���i����t!���X�Z��?�{��\qka�FZ���w)̒��_*�z^�u��{_����%��VFR��]!�~+�JeB��:2:;��b���Aj�E{����9f�Wn'~��S��yxi���5Jp�_�����D�gb�<F����tS���ΏQ-jXYiN��������		�Δ������Dw]�OC�s<{�����K��P_L(~<nHM�~:����P�	���*��.���j��M�|��7�d���cO�pu��8��u���OR�:,�ߙ��/�V����9n/%dr���%^qa�rI%Yw�tg+h�M� lR)�!���KS����F�ȸ�Z�ܲ����	`�B�1�{ψ���_RjmS\�"U��NM�����w��Oڣ
������BN��-�,�&iVP��@k>�.�,@Z����d�����r>W�Ͷ�>�%�������D!�����Y5^Ÿ3n"��N�`�W3���w��HΛd��w��~?��	��)[�B��	��]�~���'4�Dcf`�!֬	 �����E��_&���U�u]�ǳ�c��}|�+��:���ʈw~���==?6ҙ��סg��@'��hƗ&��"�+�FdO�#UUw�e��`��w��%�h�rx%��Z�<�c�9�S$==,q~�/���l�Մ~{��2�� ���iEɧ����Pcا�;8[���TW7Zu����_ EA�<*��Y��+�.I+/��|��/+xl��6�k63�TQ/〺���"ޝM$:XunkX|x�YG/2��N�p���8�y����b�~�i��z���M����;�Y$Rċ����}��I�`�⩿�8#��"P*�D���QՑ��H"�J�7m���t���{)�ª�ZmI�iK���<B3m����
<�J�[A�6���#$��^];I�@���K�f9r�����EL�W~b�}��]6?d�S<�_ ����"q��2��a+��i �Y�`�؟���<�[u�|"( "9"BOhJ�m�a�*�U􍌟��7��T�Z�YP��-�^ؠ��U�u�@T[r�E� °ˋ�+_���:�����K��G��b)�b:V
?1���-v"��T��n��(f[`����vfYҧ|�����×��W1�.(���ࠆW�O�@�18��s��`�Uc�a�h�K�HΕ���Ȅ?�>Dc�0A)����!���y �����"KM����_��u��\��wjj�����J�,A��?���u�6��<��1"A�$�F�vG�.'zPeڻ���ȍ9R�4nҍ��Q��HhP�]���s}�R��5���"��;5�����08Zw$s��BfQ*0�ׇT��b0�zF�����%)�kS��UIki�Y�E9�0X̝�(�mG(�����fM[�5n�%P�&�J��m��wA,/4���������=�(���s���2�b8p*��?�L���4�#N��N�J�{�Зo�2e���k�ԡ��&z�l鉫9M�_�Bf�=��e�i\O i�a_�sz[��pvDGd�{4�	�EG�9�9K�|T�?=�*�	=��kDj�ŷ��L���+Լ�����z��l@�_8���P�XF$�d�e.���\�2����#�T ��i�	�_'��F0�����X�Jn,�*��l��v��7�p?L������`y�'�Q��u�C#��K�@��lL'k��\R���Kw<���/�����\rNW��nm��G����J�+D�ZLo��K���[<l�X㡱 �"���E�@x3a���5#A�7�(�_yĔ�=�[����5�J�%U�v�� E���#�1~h�a|Ҟh�kc:%���wrQ�~��:+;9
kJ��[�� WS��p�>���]�������~���|~���͆�?9�A���Z�{h�V����`�N��A�x&��j>�F��^A�� d����r`#�Ǉ{��h�D�O�c�[��a�o[+10p�y跗�r�w�rd���-�b�����Uö�G�&%�0��n��Q�pm�\�X_SB�)*fQ�{>'�?������\����'D,X��nt�d#�\5�h��Ř�%��t���j#�� �&UoDh�����=h��NR�G��A$�T�Ćւ�,�Sӫ1n��m&�y��KC�����i�M+QE�Ѹ�ħ������F[H��+��+�\�\0{����TR�n<�߀���s��~�8p���pÕ��غs}�-"�π�y@I��:�G�⽥He��Z��_i3Vx�z �֓F��u�������3y��-w�����\��	oJY�Uh0���1\E����T���'���\�E��ە6�QW�J��@e-���uA�28��x����8C���T\�5�e�hv\\�T(�A�1W@�Y����>M����)��e7A!�d�('�
T1�9���3����z!��)�Gח�K�w�<�~�nڧ^�����E�*W���I��t�cթ2�"@(M��e�?�K�M������9�����S��<��e<��\�b٪��;�8[�cQ	�v�ȯ}ve�C�H}5�5hkG���3NM�'�ఝ�����C��X�n����˺�\�+���^�5��_��1�pۺP��6}���)�9��� �)����aFr�a_��nW�����a4�;ZЯd��ߊGQ��Ć�LwI��b]��k�L[���	���S�1:��zl�Xc�� �N�bp�/9���͗a=Ӱ�'^YMk�.��>h�
��}D� QMZOHx�4���}��/���G����fg�ĥN��N�a�P��GJEM�ۅ���CE���}07j/e<ujP*�|!a��K���酥]tf��7~�U�I!޶s����G�0��A�(�r�d?��	�9"��ر�G���$�#��t� C�s+���U�n_����+j���N�aU>/2��(�N�\3����:�1��]����<��8-�9#�}��G�ۖ�*����|=�'#����*�Y�2�gU|�H���D�D�b�P��>����#���r���_j��e/��IY�ZN},ԝ<�HC@@��P �$	��Ï��Z	�+Ɩ��?yzj��"�sG��԰�i�$(�]ע{R0����g���z�mE�����X�'�5��gd�Ubp�'
��C�$���qM��M^��(�:V�+�:�A�8e��5j�c3�;eC,B�5詉�~sr-s�U�2Ftq��r�"C�N$\��әG����Q�	/ͻ°v������w���#����Q��BT�%��)/;`������X����P�c��߆�B�S�	�ح7��;��1�9 �É?�`�4��,��Ϳb�����8S������i�m�s8�����><�B���k�Q�k�߾&�0Z���D�J��#	:q��Տoe <H�I��X��#ь���x�F������_2�($G]<]�h�r$�\O�	���w�ĨT������� �=�YL��#G�n���w��	:��4ႃbym�߂W�C�Y0y_�*h-������ޛ�q[,���s�M�.1�L/N���H����yl�xeTWe��v�Ɇ"醫=R�:u[���o_S������/qv��~R ��|l$��+K%��:ώ��$x����c�r��:p�����l��c��q�z����U-[�)g���eȔz�bXv���[�yV��A����@�\4�3����j_��o.�N�XIۇ���it�X�^���F�Gb
�̈4�_�c�W9'��g[K���ٜ,�*	�^,�7�����T ���VH,�e�ҩ4�B��|�v�ځ�C��W�
��6f	Q-n��͇v��Q�B��غ�}��9���Zwz������M���Θ~j �V�n��"� 1Wʛ �1��3Z�@pg|���3���Z�t���;�ʰ�Z�4,#ׇu5����Ke���-���E�گV�Ͼ�E%���O%��MZ�w�TN�.rϐ֧��Uڭ��iе��L=n[,ݞ�J�w���὇�#��Qꛮm�h~�SQ�|���d?�T�<��y�YB:0�絓��C�7`f��/)�"��;*l�]R���eH���T����O�/�A5w�r��9]ϳ۶	鵩g��2� |��@�=c���oY�9S��+ޢ��g�2)���؄��u�^�����š�9�'LT�t�����K��;[�w���ri4���ц5R�#���bڬ(�1��w&u�ч�9� ��8��-���5�f
� 3�	c3��ׯ�h���X�G�ަ���%v �O�<��	� u��}�a�/�+����A�#B�|���;�ϋ	�%X��� l�Q��|�V!a���X�?���
A���,�j	�)����ҠR���Y��V����go���\�:Y}�����A�O�N�蘆ԯ��iw�C)���l�	�vP��^�o䎗�lm�\S_1mf#T}�y+:~r!vtLFA�A
t�����c�#�����0����A����%��
]��;�E��!�8�~�jW����J1"z�X��N
��|f,Ji�0a������'9\�ֳ+�-4B��k���n�n��*��KW������<�������bB_Iᾛ���'���l�F��j(�E�9��Tcmo�f|���2���su�TZ�/�e����7%�K�4��sx��"|X��5N�����y.��섨�5�`օ]) s3����M6�C"�C��0�e7D-�R1x���W�@��T�X7��W(��C�����.6���q���&BQ�"O~ ;R��˃Ou4R���B"Au񤙭5���O��M�����@Dy�V�հxF����,\���;��̄S�5�9Vq������J`�!�5�>�m�2.��I:����U���\Ǳ���D^		�����_�e�Z#,�����_���i}��a��~̯�$�4̹��^��Pa��Cz���/2�5|��j��w�]��]���p�I'*�u&b�vr�R�؉d�5�Sy������B�s�>C`�T5=߅���F��-�H�H���+J�$��V= �+�MX!2	���V%Kg�^R\/q{f��K�Ͼ﫩�����H!�J��4�D�_���_��2�g��#.zՎKૹ#q�kn�H)Ȉ�#JXڣw�Ǵ!\T�sS�o}��7�5��������Yn�u�M��સ?�B�P�ID\@�����3D����e������Ʈ�S��
�s3W�^�G��_��J|h�{w�9�B�1CM�6���a	@i5vʝ�oi���|Ë�h��g��Ņ�%7�l��PY�G��&qV����N�(��cQQhHRa���͚�8�N
�Xy���BW�؎-$Y����1)<�/r\>+eKpC�}7�z[;�  ���k�(���C�*qr%Z���Ri�ŭ@@B���S�N�<ܮ�:xN�l&�����` -�ƛ�
#Q�K�յ�Rh���A�i��⌯���o��P�e'̢ůΉN��x�ڞ=C��K�� ���O���͟(�m�h��.�8��-����K��-��n�!�HTdl9�)����h�r�Gcd�j�yvR���|��zj������nw�>��XIiX�B�j�A9s�8
pp$,��QE^�>2t�\���OR{)[+�]�?�~�PۇD��S��8������4ʾ��ģۆIg�@{�B2��D��4T&罍4|#m.r�t�i������O
�0�+*�rgD��I����Zm�{��_+U�-�:".�����Ȅ���-I��M�BO?�Oh-�Th�d��K���!��|��@u��`��7�"]�A�7�'�iP�)S��KJ�K�CEl#.����֥w{�R���+���]�?�5�9_{� �{��rN.Il�<��^KM���k=�*��A���/���mV����H�bPA�9�&-|��<Ʋ}�n'�;ƌ	y���(nh�8|XobRVYL��W�bG�����[��A�/i)d���l'�UF�'J�Pۏ����g�b�rU2f�@��#��2	�e��};�3X��`��(c'�	������d�����N`�{"���Yhn��!���w��ϫ;�u0�&b���A��p��E�Ϭ��Ɋ+�1�\�V5O�B���f�t�ؚ� �F7u�7�A�tK���4�%�d�q�(UDp��f�{����̕�� "}#ՃF|mo�M�<�$g�G}�l�k��:KA��/DƧ��*s�VP�$�����T�r�n0�C�~+��D�_a>��%��N������<4r=|L,zyaSG����6vO� ts�������׋�s�¤y������^>L��	���d�ldMP�jblQ?�Lވ�_hDb?�������O�5˒���҅���E�ΏaA[r�����h�����v������;5p6gV���r���d��L��NX&-���V5�)�7o��������1�S^@�trP�0��O/8en���pU��M>B��Ќ9���[;��w���@�H��>İΜ���+w�5I�^#<XY\7���~�_%��W��ڢ��P��l8�rV'��3�T�W�u�ns�����g��V��w$�"�F�9��1�8���u��For`��v���M�֟F����{�b؃��}��-ĝ�AZB`���7Jd\Nn����ņ�F��4�ۮ�+��ƺ�6��s�h?��}tu9J�=7�Rk2U��0h=)�]q�ś�K����g�'���bJ�#eߒ� x>�t�/����e�8_D�����u�5Jn�Y�&2�|�a?��:� ���<�Z@j�%����Qp�cvX"	�"���)���L>���(���w�E����-�
���R�I��TȊ�)
�Y�"�C�'�׶;U�CP��'��9{�>S.���N�u�I,�^���g����ɘ������f��i���W����K��Ŋ}��8�7�]M��_b�ٽV��0S�3�Kg�6���c���6�{���������p
SrV�|��X�7���<N:������(����ߥ�Z'Cc���F�>���Y�Y��;�jU�� �J�3��-r��߯q������"M��%�!���޴�S��U�&����f��Ѯ �~z�����\������Ӫ�ط��@�'L*R6*�mA�m%��Mt���!cp0��_�����f������ݖ��)�
��5^��D'�	�����I*28�^�y�.<�]�֥�&ё[y�����̉t��HAT�%�h�+�z%򺩇�����X�\@�5<:CvM��zq#2X���������Co��R��Q�������-c0�u<gF���2��("���\�%v�Ύ���l4ȕ�f����b&y042ba��_���^���X[���ł�}��y���@Gۑ�14�;� �x�ZG��
���l�T�v4@��q���sUH�����"O��becIQ��}�N��y<q�'�-�O�y����BTI��"��Ӽ���~�2F�����o�TgN��'��5��?�7�J�A�S�&\,��Q��7
p('�ST�sm�ci�?M�$�{I�u(�M6V�����y�\}b�Զ.�@��5�(��l�֧�����Dn+#�^>[���Gk:�T5&��]�	k#���ͯ�?�r�sc�Ҙn��MJ,>�F��c$�K���r"����E9��4Ⱥ0�Y�3M�c��.NM1E���;����Zo_o��1��, '��B�!���25ZڟeKN7ȵ§kf��r�%zTX��{�Oa��p����7�S��qG�;��7M��| �Gr���.�vF;3Z D<j*�r���Ʌ���G7�>)�5:�I����F�1�����Ic@��}I  ^u��O�K!��,Wr��Ӯ��X�`��-�	�@a.�,c�O�~'P!��LҤ���<�d��������bLDґ�z����u�D}LLE��&9�I��я�֍�бQ�?D�����卜w5E.��4��|�M�B#H�.E�1n��E3�fj�vZz���Q\!~A�Ђ���~Hj�Z`�;MBw����h"w��cQ��s��9\��֕-S����� ��B�NXZ'��\?݉�^����M�^��#~KYkl4�}2��DW��u[�� ��3q��J�l¸G��쵫r��� J֣`��ea���������x�S!��T��|~8�a��\?w��	��39����g���ybA��l�s!N8���V�:*9���&n̆�mwH&8�ݲG��K����z)��wa�pHk�o�(�xD�}�l�5p��?ei�!�g���!��ޢ����8�[:|C	��}�iί�]��U;��^��ZC�4��Y��o��k0Yp0��@N�L�;	����Tއ��!��4���L����L��܌��9��$Lǿ�c��|�
�7tD����!�[8{�.>�j�se˒�vG������<8\HwW֏�	����@����^-�Xc��m����JA���2qh����d���Z������F�a�r���4G[���J��ۤ2$@	'~R!}f�5�s��7h�k�!8tY���R�i6�|�.�Q��"s�R�|���t�:U���{JD,z_8�n5W*0��J��
�'�;��-(�ߍ�/ �����ɾ��:'�M�����o��Ε|�I��Pw"�\���>VW�B��Ȳ���K�B ���&d�Q����c֊�~�xX/H:����>��-�{���e_��>0ڨس�X��| ��GB�ඵ�Q����v@�Y��}����x���TӽZҟ�*��l(͠+"#L��j�i���zR��U]m��d�q�8�P"�T��
�ϸ��/h��_���ΰ�
E�ׄ(pkk��a�a����@I)�����)�yѩ#@E�ƨ���'�Y�T�����d��`ń�A�l�
��:������ؓS���t��R&��yJ��Are\k�uf�`%��#AH�Q) ���4Г-�V%��5�0��4�e:���G��e�T/ohD�����~6*�i��/�g{z�9Ja*_M�=fճ���`r]�}lz�i��*�D��).1�=��<���ҙ�}��V�gS,��~Wo/�i�%�tFp`n"F��'"�.��kvS	�8�j�g1�!8��
k�>���'��j���y��033Tn�`k>���
����i/�ck߸o�D��I�\�	�Zn�{�'����"����mi�=/}������J����w����nOб�BzE���^�. �ñ\��f�w��{��Gұ��;Fq�o����8�}MKY3�1P	r�����r�x��H��? ��Ύ�d������O�#4��ž�l>m1�%F� �R<3�ZVl����Ǧ=X�櫱M6iph����0ܡ��m'��^X��]�ʪ���q�73�$K�Y;���'�9�?��O�B���׵'��'��j�s�HVA(��Ot���To��B�����;�9���S6�U}�sQ�qf?4`��wӞ0F���	�y}�S!+��5��ڔ���;s;$%�;���'YK���8I����a
�(�<c�O7��%�k�p�H0�����L�K� ����$�ZϞ;��G� "�.a�r�.�"��<Ty	E2���>v}x�ɉ0�V�b? @a���y��
�ŏ����0<�r�,P � v� e��`��\��+�$�Ω��S�2*k+��ͦx�ǃp���ؿvI��R`�"�36����yE�Q�>��1�q���a
��tx�9���|#"U�+B�Q�p�r/�R͂@Ê~����<<������8#�9����u��}5�u�t6��"]��;�{Z�Q���;s'�e��^�*�n����0d0$Ԝ��'��Qn��jx��=��ic�=M��ʩo���X����(�=��p��@v-��TN�j:����%A3(�|����JuW
 �͕a��K�ܝ�_��0�?��o���Y��&%�K����Ⱦ��F��OkJY2�|��
�~�������`Ϟ�J�U�����S����a���)��xu׋�v��
]�a���c�+cYo�wATxǵ������w���Wo��WxFU�5|��{���c�G�^�(�mkݜ�	a��i	^Ij�} A�<3KC��g�!h8���g�!��.��C:�Jp�#�	�z�E��%[S�k0j�u���j��КAM�y���'��A H�?[5H���W��\0��=�m��찚�ӝ���'F6���/�fOzKQ�9���l�Es����Za���$҆Ѝ�K������xOV*���3f�L���;���	���/�@#�[xp>�J��0;�N��ҥ<�Lg�oԉ2�M���"[��G�����]���i���*ƟMF��80�*��쓑��n�ߑ�� i��-�(J#��IWU�%vͧ|W�A�T]5��g$%&[����$�np�o?�}�������]�{"s����_뤔��y�
�������v^�4D�����/��f�ln���K�t�鴯]o���r'>���?���b�������Z1[0��=�;d���9�i�Ơ3�SH�M&wϐJs4IQ�m�R[�[�MC��q3�᧝���p� ��Um��vjX@ڹ�c��l8,��E��������$�P�a ����_���V�M��Y��!Z��g��`9� LAQa&'�