��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~��_&kQs�\�K�v-�Y��!�M�Ɓ�����y�I;|`��e��懌Tv�fD������>a�v2�oEo���\����*(�ί��S)T�B�p,cϸn��c��2�b��>ޣ�HQv�j3�0�w��M��7�U��yzC+�Oic�&a�֏���hy��ϣ0��o��"*�t'�|>ڏ`&�v�EW.���5Vbg]�P/��M��a�����>C�Z	_�o�[�zV�P��#Z�]�IuL��M����t`'��.h�_��~��CC`1=ǎ���G�K����5}
ՠC�2�����,�<��W�ƒ�"٪+W8�ql��t!	���z�[0ؖ���I�T=�s��x51��$�{&F�~�@\'�CѶo$p��:P��\E���V��.x?:b���b$.ďV�}ѿ��}rr�ȏB}��/$+�1�g�V�(++T����@^`g����4�}u���4D{nE�sO �AdCP��\h�F�h;T���쩎)�.H�#���:�-r!���Un1p��E�Ӫ=�>9�W�$d���E�hb��h�W/�+!&T���0k�Y��X!/���Xg�&�h���l�>��� ��Gg��\;�����^�2�o3��7���J���J���F=������C����+��n���	����?NO�g�)#W:L|��-x]�{6(�ٲy�������"��YH�{�"�Ri�4 b��u�|�հ%��"�j� � �����l�)$��t�i4�ܸZ��J~��!5�qZ]�"���5J�vE>`l'�n
v���������$
VB_	Ƶ"J;���k;\�.�B��%��Be�.�Z�Cڃ��4��&>��Z�?�2�Z�"�A�W�s{ƒQ��\G�]��_� ��1M0 �n_~v2�=2Hr���� ���%���%�S�����q0S&'���6~�_��~'W��DJJ�dĪScԭ:X��@7T}#����(Q�^�G�obu1l�l�ӕe*I� *;ȴ7�9f=V�П߯���Ɵ�I�\�F2e6Ւ�Kr����c�&��KM������Vứ%��ڶR���& �o��V���-��e��1��Y�lZ�B��;%h�sOp2w�`8.�O�������רv�5mL��#��(�hw�M����x��咟�Fof�K��nΈ��63��K!dU��|���pzO���'�>]He] y6�WE�b5H�� �n�sԜ�0�p�Y.7`m)gݱh6F�%m�k�!�T�����S;{L�v�)�9� OC��ÌC���]�X�wd�7GB�bC����{�H	��K`�������Ɔ�?���G��J�%�:�i".�&p7cd�ȹ�G������#��#�2�c�W��Z܈ 6v[y1櫨��dL�plv�&�%�+Oҋ�|�)��29��i.����,({�=L���d����
(�Д��D��n�G0�/5��ɹ�%d1�/�R�8r�#�}�I_М����|�D�r)SU0���N�
Gƺ�Z��9<@��zà�`��$#C�)����+�*�E=^ ��҆���/щ�!;�x���N�!��C[��M��;��s@�.V�;��NM8�Y����Gl<=}%ގ7��w{m���_�~�?�X�< ah����|�����@w�Gˮf_�{ۇyJ�JI �@�wZw�<���d��h�f�~&�˱)�P�Y'�y%[f�F��4E(A���_�P��=��5,XEx7���[��Μ~V�������:߂޷�/E�Y�IyĜ0�}�90��uV�7�䲍���������
��;�"��Y��wRt�T 	'���!ȺH�dmu����N�'-���G�j�A��>�I���\{P��f9�g�<�R#���-�`Y���=�%��Ma��a��,%XA�i��^7�pG�&���v>�V�Y�$�]�Uec9��bs��{5��$tR
�恸������ְ��ĳ�!�%�4�ai��z�Q��Z��N`_��(;g5ǚ~�����ѩ���2�!^+ñ%ם�Ӏ(��E$��ۆA�'.#�rf~L�Z�H�2s����Ry;�#�F}b��J��;;�HM���L����2�23q�7�ٳ��u��0��g��4��"n<9���Ρ��k-$st�u�>2��a��.߅�UxɊc�O��_,�IO���;.��OV��������Iq�˥��	%����1����3�F�zZ�:eT�G9�_|_7dL
Qo�����3��;U�m�?�,�/;2��>�S!��iI)r�N�V7��${a��oY���T�"�?�,%��Y�����sy
�i��M"��,K���oA�7�ɮd�*m�󓲆���P\�[���8��&RD!�͢xh, ���Z����hN�M��lYJH�SѶ��99#M�����mF���"W�]�n�(��0Gl} �#�1�uVfH3sح������Y�~���`��g��̆�ڭ���k��e<���D)�0�DI
�|a�	V��_�`��:�d�J}�z�[*r�6ٰ���B:=��s:${Hdؒ���ꗰ�Տ�t|�e�h��{v!�wu�8���*h���~��Fi��遇�/�f�+�u�'�s�V�^a[��1Yj�=>ϧ�xF��yIn�X��ꂪ�!f��c
�p���~t�v�N���6��Џ�p��"$3����x��=`?Ĝ��=5���8<l��p�)	Q��Ҿ-���rU�z.���,��Th�Z�~�M<���C���Z���9�>"_��Q�Pd�_���!QQ#<{~�ϹYN,�4 u6��?�hx���5�YHQB��A�H�~I��6Wj�WX��5)x6���ƔAI�%%]�j�˽X�ҹ5��E�B���er9�3-k�P;q�e�1��I�����O�t�6KJdy����N8)A�v�5/�!٧�8·;,��Z!�Ǡ�Iz��;PIr�Qϩ_e���*�n�˼hj'=�*�L��(������l>˜)�=A�)����M�{~�p�i�S�j�鵠�\�S悓S��SN"PR@��.��U�)��ș%��h � _�-��]ɒ�S�1$�r�mTR��zM����JyB�[L��s�x����B������(*��K��C�c����G��wI�|4d��|r�lw����i���A�b}n�q�KӶ�䉊�u+~yU�n�����p������� @��_�I	 &�n>�;�pZ[A�yH����F�I<���.I��g�2���;!�,����2]�^��:G�����'Z��������̷��w*�l�ļO����&^!�9�<�3X�Q���!�c�X�����6ˡG\�~ì�A��h�*��M{�{���K��e�l��x+�
����Vn� �j9���ŹEt�oH�^ק2�a����)ǎ�\�ɢ^;�� ؃���~��Bu��^rZ��j����f>��Ex��\B�s��w�rÈ�&���#���/�)(�Ȑ��w�N�T�*��n0%'/�w::�E�׶��2�t}_��>�o��2y@���2/����z�h��������H>l?��q>ɳT�{UJ��0hh̹6%�_-~]ğF�+u*�aZK�W���k���Ky븠v
�`lu~g�W
��j�ET�*��ow��_sT�Y̺ V���GL �)��ь��=7.�>F�}%3#*��Zi��V�Z�@əMk��c�K���{�UI�3�Z�e���������2�K������x�a1��X�����R �����I���_j`����U���R5��d8��b�i���*��Yɉ���1"*]a��G9@JUSqs�K]��;��"��f��	�����Idt��j����9)�r�K
zB����#�N�F��{�\�׶?p2ȬPs�l}k��c�IA��4*~*��t��Q_9�?�
���K�́���I�¬��n�	�Z×`�B��-�P(p�?ك���c�F	��]�Ҍ!��d�����K�պ���Q��'G�+	��)�^/5��5���j#B�j#'�����}K"�C��R���e���)"� Y�Qq�Pw¤mV�v%��ğa�j�w������4(��Eª��T���A��~��I.Ss�i/���x:����|�|�1�V���	�O���~=�����3) �вz	�߳�0��*T��ͭ�[`���j�g��F�p��{a�dXVD��N��>��Zw�de9��A��W?�Bl*�ċTS�j���H�
�ۥJ��|���T��9���֔�g2����}N鯒m��b!4�h��Nf�k���Е䰢�$��t��B:w�_=N�S�x  W����/O�Z�q+�U 0wJ�`!����jZ�\�@���b����>}"Ēܮ�X~�R�2�?��;S�}�� ~����G ����E���6^)ی����iB,����R����Hw1�E��TN���5���+Uqix�������R$0�T!�c��U�[x�+�ap$�xw�:��Q���75`}�!A���/��6�{�~�I���r��خDν_�^�Q�ʼ�d|���t�
N68#�$�8z�_@,׬/xW�Q��XP�J ���*b�M�)�^UÖk��7���>�@"f�~�Ԑ������7HN	(zY�z���������D���F��Ł�����!����z)����_=���F�����:V+	a�9'�SG5*��������Zn*0ƃ�� j�
 =�Kj>|�`��m(= wb�K���6w�
��^��C��
'�M���W��ca	��M
����
͔��mܫ>f������ɚhw���rh��-ӣ�¦W3��S���Gzcɲ�����j�#*$����a���)B���N(�)��uO�L��}�G��g�+�T����Mǐ��4��	��^�w&��� �"͂b� �r�%$� �L��DA��#�Jo��x�+{_�J{���=*Eq�B=���u�b��+�0�������BA������=�VhI��ʤ薽�zO�4��c��%��MIЧD�y��k����J\�
�VE(R���96���]w��K*�e]�CI�M(@�����>� ���T�ɮt�r��`�<��L��O�E�.ݔ �����V���^J5�+�%�����ح��+H'fT)�{�ew#W���46��}�[DaM��Vi]�,.G�_�ђF��µOa=�
�)?fV���$T��ې�%20�+<�N�3\�X���Ϥ�5�k��jD�h��9����1T5�Un(�"̦�{K���,��'0��փDj0&���JҞ��AA�ĳ�����J�d4�"c1q�%�����AB��]v��я�����WKlr��w��9���[�5�������{OWe�s'�9`�Ǌ$C��T�^j]�/����S=���g|Bqi�ٝ�+���-���`,���*��6�^C��[���G�W����хA�I
k�W��;`_���T�J��;ȗs�.�,:��u����~��Q�����f<_ux��~�~s���p��:��(����ߜ�X��b\*O�ں	F^U�P��H��t��9��v謤 vi[G(��R/I��Jk]`�o@��1�i3L��OͿ3qI�����ǚ*?�VHTj���8w3���	�z��)凃p�z���%.ƽ�5�,�؋ۣq�
H���2�Ƴ�qK�^���붸5���e��:>#�O�2[`^> ���U�G.�;��C{SX|[���֯�uE����J+�bz.엥e�flq;���YK賓f�w1�
�u׉M�r�eyF��T��"j���v�o�[��/�ٍ�'�x���!�j�H]�4-���*>F/����⦈Z��Ü75U�R��7�G�=�k��[�Y+#L�ŧ�cu�d�ҷ���n��1-僴���,s�p^��zlIw5���>ˬ�[��鯱C!n���m�M�f��:�#���S}܉��6��T�R.*kue�;�x�<pH�OP�6OW;�����]#�F���P�G�Ai^:��T�)�'*�7Lu���8U�"Ism�����h�M�Ƽ��%��[cY�~&ǳ�V���E,�y��'� J�[C��#�%�������T@����6tCrc���H0�b��!͹gm����2o^1��mF�=I'��9;FH��U�:`Fo���p��
V>�H��ᆽ�Dto��]W���?C|���Qp�z�F�.�P�/��ţ�3��+|��yj��3�a�R}�������H���Ƙ5_���`�
S�-Q���Ψ/��+���~��`���c+����n����\�K�%��'���ϒvG\C*
���"��*� ݑ��zD�?�(��X5�����!�jl��0/��W�!r�����.W�&yPM�7}67Ghq7�+ULO̔��;7!Z�p(h崎�]�9'���t>�;�IZ�t7��s��:�b���t|,ل� g=���9둆����^3���é��/�j�J��9��qϚ��3�.�c/���UP8��2��gE=L�窱�B��̩Y]�  R�+����	��h:���犯9�8u*Z�
�������[��3��i�.RUQ�>?/LM�0�g�5p�kZ����s���,ۀ��7}3)*�a��|!@�Aw�ڦ�%쇻 !^�$qs���t�	�-ӊN>�l��-��$���s��
?�0+�-T�-4>��OrK1�/�Hh55�@]x|�#>C���O;��^�|�)��Kz�J}��E ��A���K��^M�l��8���mJ��7G`}|Zd�Z�2����| ���뤲�u��%b�O@k������ �.�=����� ����:��-N��{�B~H�b�c�ؽ.�l�'�;8(�{��A�yj�`
��B7�;�+,��]uv5a�~�����3$	���/4߳(a�J|��DI`� �^(�>�� ހ��I����Sz�s>;B?'K�k����/�9���Vp�K0����o�������4M�k���2:��A�f1EA�S��C�T�յ.����C_����t��gt�6$�u*� �g�<�.="ڵ�^��_&L�㻯�[�ꑶ�;���G4�ߤ�MG�Y�<�3Q~���~�I��͏�z�[��B���lg�ɮ?����k�Ȭ�