��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟx�ɅT2n�x��p����Xh	H���9�Ҿ�z�1�� dT�h6��[I�����B�?Oq�_2�9Ӑ@�p���G:26�[�6T%,&'�#JeR�+񸊎2�Դ��E�Jc�������5N�{�����Jz����+�:��G˦�<�_�	�'��k�Ov-��5l��|~+��,�Z��r(?�! WD_����J���K���םcE4��%2���qb�B^���p�G�A�tX��~���tIݹXT��Ps=^�����a{;h�h�u��@9����*1�\^u���x�#�X0gR�Y@Pt%E֠&��-�?�*�ݎn鑷�-��E*F%�}��V��?ZҀ
�C	:_}�ZY`+U���۞;��F�U/� l 㹄�<ĕ�1#o�Т���{�H8r��,�W���5��V�[N��S�T�2s;�R1��'�v3�����0�o���֑�8�ea��O��ֳx��@��8���ت����H��_�xD0�{�\:b/�!�LX�R�<F�$u����3O;?a����w剹��y��\�3{=4o�>ԛ�F�M�� �I����Z�u����f �.�6T�z?4P�B��ߩ[�W�\$��W��� BdG�g���گ*y}�X�>E!��QY�iGI��v�*Еʉ�F�pK���9�vЮ�=���	�g���(p��E�����jf�M��=KD[QhˍJ�E�w����Rnf���~��w�aG��s!�|�E�������v��*3��1Z��'D�$sN�v{�4���;��Q��ŏͻ����wiH	�he��)�4:��J������O��I�h(�;%�BF�)MD(��B��of� ����d�yVJ��'�LQ��W-�N�ˏ�+�e �����?�?m�#�P��7G�3��P�}��I�� �'�Vod�C����D��7t�,Y�`��kٰ��RDc��-�s����1:e��"��C���b3;��gB�S[�	Zh��Rn��!�'L�Kp��H�`M�y*2f�fduZ�=��}֊�_t`�Vg�SL�.6�5V����M�ؖ�����n-y\O�I������b0�<�r��'$W�˩)Zs-2�dN�k�PT߫f�F��i=���#����C$s�vZe3w4d�1e�i�d��Ç�`@����G���N_��g�<����Ą�t�e�W*O��<�P�d@�^4�6���i�_zO�Sr/)�E8@��wH#���y}����O���Y'�B6�O-V	ǻT��S=���X�V�@�?�Cjr�Ԟ�[�w�@��dS��a�0a\|�gGs��	�	�EB�;�9�r��\pŮE��XZHY|2�'Kw땇��>�]�#�|��}�����(�4$ȏ���S���D�3a��ut*,���3�Lx���|=������e�A�5�iI;����0�	��]�pCA�TP�G�A�x
��yg� AqY �u�b�c����b�e#}#������J���$�XW��Bud�B�8]�胗ř'|�B/�.� �0�D��{�a�MV����.�/��������΂ڮ/5�t��+�h���dzH��I֊a�
�=a�8b�T��+2���0,z��X�lZu;p�ȦFLK��C$�_�A�m�Oˆ�*����~�+T�S�Y^:XI���VH8���TD�jP�f-���H}`u��N��EesFs,��^TY�T�(L 񊦖���_���>�`D��x���;��Z�rdq(���#%�D�F@b'��6�b�V0�!���jy�|�ާ3��n��>�/;�
\t�Ae�|���F{hV����Ocsa��2wzRX���y3n�k������ e����=}0��Y���{M�:�u0.o����Nw|�.���!Zm�Z�EN�d'_{��Rq�j�<Z��yw�D�eb��><�.��z�c2Sd��
�4ܰ�{�U�p�b}�l���}�yΒŠ1S�:��So-s�!_�i�&>��$M~u+|�P6�!��$�b@)6P�U�^59�Θ��-RP�Z��������G8%YSK�(2��#-c���xZ�5�"����z�%6���y�t_�`���Cm��gF*�xN;�<o-�f^�i���B��z<���E��%�2�,���!����Z����Vh��e�D���	�TD��i��ѫ�3=w�S�g��Ή7`�E(�^e*2I� Ad\Xq��7�j�%Ș �Y�?f(}�	JIk)����D�n�ѯm1�*�����	���f�pj���tіx�E�d%ޛ��C��󔏒lP�4t�����\��+�Q@Ɛ~R��MƈV�1�TZ�fK#GA�,D