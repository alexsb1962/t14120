��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����t|'�dWJ�S�ʳ���t@�~�B�a��f۹f#D�H)����=�l����E�����'" ����o���a��v]�|�}h+�#���U����%$W���m� �	#M���8�>�PWޕ'��U���<��\�T1Ua�M��,�A� ����Uq ����sHt�}���6M�jAr|y�$�
R7a)�
���k@��_d�%Ǐֱ�=Q� ��[���>�3���Q"i���I����oA���̒a���z���Žg�L��� �M�R�T`>��EO�x�G��r�d\����y���ߐ.պ-�~�D��^���
=�f����[�Y�`2%�W�4�o��t�"����}#����=���?����7t�����g�.�-Q�D��{�L�'�K����C���-�o�X�=�|��vע���_��U���?���n#�P���f5�ϣ�s�V�fӯ���7s`��tt���Y�54�7��܁��hql^;���7�V`i�8�J������H�=��JT!:�$IVSB��ȷ���s���sE��Xt�tk��z2;��ޙ(l4z���Tr��Dr݊�����
��ճ���/Z�>�j9>d�<H�©Z���m�C",�21�[�,����,�s7�W��Q\D��1a��+�wGu��s��f*��B�b�w�dI��~��h�B���N�I�q�_�7+��M�[�|-c���ɤ��4��o;��l�	��?��d&in'�}J �o~z,�q O��R�i5�
���Mn���<#U�*r}��vq9�p���͵�����)2��rp�� в*����	D�e��[�W�{�{Vox�����ŝ�v�\�V���~&'5��r|�Z��?+ǔ=�.��u;�['��←a���vs�!�lt�����2ew�q9�ְ)2��rd���1��?�B���=���R��Ct���1x�	wYYd�7�Kx�/���}���@����O8z@�8��n���(�����o+Y%�n�Q���г���"��ն��3h
R��8�<fn���6c���!�bӎ��QW�Q�@��m�mx"����Q���W7ݞ�a���FG_��s�����#C��ƃi��Uog�-{q-�U�_�����~wl裡v�U��U�SjD�5).��қM��?s�O�=	Xw�������.`���Nby���|�$!���kO��n[�����U!"Ʊ�ʵiKң�Q�+�H.M"�.$�:��w���ԁ$Ґgx@�@�6�p�>&�a��
E�eln�h�v���P��jYnb��-	J� ]<A�Hu��[�S��R��e�K�"Z�#��B n���xU� g�R��f�+8�IHV@��:��*:
�^��4N%��H�ʭ)�Q���cNǗ�Z��$M�%�}��7[�K)O+��f�|��%t�Rou3��AI�~e��3z�˜���]�>9*$"n��0����e�:/ܶl6�����EUf�%��٣C����2 ��`T4��F\��[��.���(��$�^��IU�@�|ʵ�Kj�MT`�'D�B#{|k&YKSm�x#=�c�]k�L�Z���#U�%;��V�L�|�1�K9[sFu$�}�F��ER�SV��hL����T��ӹ�I(�����W}!��d:
��W*�Ý�e���J?D�ĺ�����98��zQ��{�ʪ��Qc�s�����X)琏?1~�����X@�9$���M�@#i�W��vU� .��TbRȀ:�[�"P�0S�^
E�r��j:�-�+Sڧ������R���!����h�ǅ�{`*=T�s�-�K�����b�j���d'`��E%���x��Hy�,�����o*�����0!�4�O؋�F����k�����õ��\I5���$�q�]���%NW�l.��P(��x��"�KXy�Xhbڭ�o����>���B�|Ǧ:��wګU";��j�A�֘t`�k�b�����9��6V��	�r�
J�=M@B��U�������"�"V�Cy�Y2�rD�g��4�<�����q#o]�L�g�蠿u�
�+5�ߔ�iZ�E����FӪq dƜ�>Ҙܸ��:dr�.e$�0j��V�cT�y���b����0u���p��9Ò�Rl�!K�Fl��p1Uf�B5�x���
�Rm<@!�J�K8�y%����G�锁�[�j��pHVk�G7.I.����O��@�+Df��"�hi2�.����/9gzq(6�A|��k�5�c�,��$P��Q/���隱T7F�9���z�l�f�`�Z�������~��k���Q�M۟[�Q��  x,'�rIS4���/N���G�{w���(�x��(���	��+��v��c��R�=N���^���V4���az��b���ϛ�Q�s�~5�ٲ�+���f��>zz�w����0���������>�~oS`�ʰ��Hʰ��XJn;Vŷ>W����P9����)��B�r�'떞���һM�0�D�f;��\e�m�H�������^�T�0����wb=���ҳ�	������ݘ���Z�~S���-�M޶Ͳ�l�ai��}� n�'fT��z]G���}�~��ܬ���-��0&+m�b�$��b$��W�jvK���M���<��pK_c.���� >h�^��B�o���ǥ���E�0N�`�U����R���Ŝ���<���8H�K��?�|� �8$U�<���J�R�Gn�C���B{���������`>`'����j4���`R	��>���Zm�%(K��`�+�+�eP�[�^�>��z��CN'0��G�ׅ���vm�=~�|�)k���o܇�I'7�8{��5H��e��XۆK���(�3t��.�7��5󥯁��˒��;Ga=�]��a�\��ݘ���2��p��	g{�Xj��-J�~���`���ΚX�!}A<Ae������Y~唳1��ZJ:�5!b�`�_)zQ5�&4�\B�Kۋ9ލ[�<��	Ę�ˎ��(O�_t?,��.#p��o;��$���Լ��̦������HBI�$��ne(�qQ�A�k��D�׹��bRi?��`n�WA4�$t���T��, �!��?���T�����60�1ƈ�Kjҩ/E(`���9Zlk��X#@ƚ�h}5Y�����Ɠ��?w�"�,۠��n	�'�`��Xԑ�)(TG����F��؎�I�D�Ϙ��O��U��Rt�!�Ղ��i��=�U\o\�������{�PH���q{Ue����0�32�f3)��ǁY�{�������U~��Z<VQxl̦�1%�G�J�:9y���τIr���-Ŷj��WL�N�����y�=Ɔ�� �R Q�ʰ\
>w-#��Q���Jh��ku�)�XwLq=h:R���18b!н��Y%�?c#�r;����3�r� ����)��N�s�.Ka+P���m& N�B����>Y�>�iG/�^�� &[1�ƨ��.(r��&��v2�l�:�%�9����AɌ�S'D#�[/=>G�!KW��A�,�>��42Bo������^�0�rZ�Js���5��I�_9\�ox݁��_U�!��D��h�<a��k��d�FW.QI7����	~��/%�{}�;��:<�Ve�����z�YgQo�S4
� )��~0{�_��}C2*���}��M�"�E��Z��Z7m�<�g�6��g�3~��1껯,ðd�i��t���H�5>#��K�BU'��Dk b�+C���ͯ�� F�u���ut?�v,�����@�V<��,3	�����\Z��wc�j����ʑ�A>����(Jx��?y�:�o�d� 5����t�`7����@��o�O^�Fw|�	�mY�s��h�4��t
O�g3����g8Jda����zv8e�N�����YG���枞�T�tyQa��i,qѴi^% Y�0�2�3�Ap|��w�׋x �,��.Ň9q�k��y��5�hx4�x���0�X����W���r�=�i3&�i��E��#o����i���7�\H�Th�	)�~~ 9�;=���	O)�I���G�;Q�b��/nr��r���A��8'˅ݢ��H� �8�9��/dq��U'�TK4���;A�� X�y�9������}��0�X��c��
�1*�-��羉s����wY��j�)�tX�	���+��{����+`�=�;+�ؽ-�,<ܢ[�.m=W~�0��g ��=e�#7܀����rzd��D�H����Byǐ��x�mRV� d�?����F��mg��bb
R��ɚ ���լ�~����˂��y'+~�D��J��p���d�{f��|Px�f��S�.��YO���")�5�W�O�J�>B|��(�Iq}�l>E%O� z�g�$چ�:�M�k�l��si�SR���EpL�1��b�{si���X��1׺,��{ٯ����\��&4iC�5G�1�
U�@Hs������?_��կ{�!��e�m�.ﰱ&JЭK�Kv���cjxۖ��V����	�3f�R�!�hU4	GH+p}<�^�k$Z�r�=���/�R ��If���r��3���+�ȗb��[�7��M.
�^����30@&$0��P���.�O�����Ѝ�ʌ}x�De1��t2d�S0?�.;6Kfb1��\�V2�dM�U�ϋ3��3�II�f!�[|E����k�E[4@�46H��V&�o�\�J^Ʌٟ�	F�2�"�-D��ԑ4*���9��E+7�Y)6_�д�n���
Ņ������[<퓏�F^����q�X?���v���:�oGDTm}��"Kfi�_�.�O���6*���A��A�]�����_��8uq����^]�#��7Zp3㞐y��q��t�������S�s=<��FP��J�^���4��u�ʓ�A �V���"9����#Eł�B�����z�:ȗ ˪v{R�W�ZM3��f���
5ǿ0X-I�M8���A�	��������s\�Rg!0u�>�g�{�5�\I�Lj^Z_���U�����&�N쒡y��c%�aX����n������0��0�t�eFwH����aTơ7u0r���2
#M���C�/dۺhRS�+Y�K�"�)!�h�?��;p�݅��d,��"��f)�f���^ǂ%����9�,>���[��-7��	4!Ʒ�"��m�p4��_�	a���`�(�R��;KZW��L�J?�Ԕ�OW�,^RH5 ��CA�b���RSG��A@^S��k;����6H6�x��f$����X��{��d�S/� E�����y��~�̀�m�AѠoM6�l���	�1	�Bai���Xp8ӻ�|�)B7ÀC�����Kh�{�b]�C:�-t�,=(Ľ!S]n�����_�XL:0r#����罏�^{�ffn�ɞ�qP�ތ^1E�/� f�ά��t�X�(�6yx�$գ̴��� �;-D��ęYOX3a�i3�Y��G���듰�D{�Ŧ�Vs�us�V�!�����TF\���ǭr���J�X08?{v@m}L���J�	�D�[�_��"�qS_~�,L�~�+ 	���Z� �zF�y��`J|i���sb��C<��)ݏ,���4)F'��;𴖼�Ԓ���_iY΁�'���?�al��& ي�2�ݍIt�,ߙ&�k���~E�	р�dΫ�}O"x,㮧�|)I�ݣ�?����	=�4���4E:�\E�>/V����W#î�m�g�aWi�3��^������f����F��ޅ���'�U���:pW܎�-eNHd��Fq�k'y�uPJ�Y�?�P!����rzRy�"�L���˞r���5����4�,']�T �,�߲�jW��Ր@�3ܫ^��H���~�$@~���ng�ϴ̣&��X1�
U�(Z��8tā�������[��8"Υ�Oửg/y]s�a��jpz_��ԗ�iХ�'P7�C�n�T�n�}`υ`� ��Fg �7��ꕏُ�i�'�R�7��o�X���0����ly&]5
p�(��پ�Vt�g��r��ѦK��M�,%��e�VI���}U���R>��H}~�~�{�8��p�DR�Z�wkS��D���=����N~r�S�X�<P�!�Xgr�	�?��������!*c���}��j^�{�<D҃� ���m�;4̟��������L�L�@.wߞ�A!A׀���okVG�2b8��%�jV��
!�5��̏/�� ��<;�yI\#�3��+�<�����_5����;|e���C}�/���W%��5�T�9(T��q}�L��B$�vI��K���8!xԏ�}��\������,ȶ,���~^�#-x���xf��+ӽ�����v��t�B���d���:��M:h;y��6������[�!8�m�L��.r@7j��/�F;� ��N�H7J�4b�3�;�V�����&�4uG�4|E;�|l�G�c?ظ1M���]x��s���Ñ��zp�9�����ǩ�V�o{Ķ򌋇m���:�|7׸t���Ʃ��s���/�~P�yc�`-��y�GM�w�4��������,UUTn�ϦH�f�բ�Lʽ+��P�:�8{+BM���m ^�S� �<�ZB�P�d�#��n�R�%�:ܥ� ��*f��`�Ȯ�]��h�|��W��]�]ۚؤӹ���Gb�S����^��;V���8�B��fњζ�N5�]��`e�) T�L�2��jA�G�>2�h�^�����'���NS���sO>X�_�IZɌ��t��F���E�󹮰h�[4����R�*�1�-�"����-(Y ��ug��R��3�=5���Z��o :0|�����SH��U�:��QXRſ��8ef˄p��zn��=���0	����&Յ� l/)��Y{<�ٍ��~$*4��C�H����1�՚���D���o�ޙ�z?�H�9�� ����$���}�������u4a�h��L���:�]��_�鯾���e�'��+Sj1u,:\�I�	2[ �XniCԻ�F�qV�k7�p�L,/�Hu�򰣸A�'؈h��U�)����k���TL���L�3NtH�R��qyx>c���ͽu�7c�:$\�\@k�T��]�,�բ%�d}emU��檹u���DW�q}^��)]�}��`�h���}�%�Z�N���TAY&ʜ��Oj���J��@֕�	���:4h�me��^s�-�����#>����u�'K� ����?04R��ݵ� [���8�p�ir`p�P���^����X@��j[6ɨ,��U�B��s
m����L�l<E�?]����7*�l�z�]��J�k�9��QR8&�G�.M�ZI+�$�V���Ś�ۦ��S)��6���!N��.1pA��w`�b����m\��_'G�~�J����QL?h���b\��8�d�Kc��5�cd�r0��'����Z�<J.5�D���]":x���W�������J6�1�K?�F��8�)�z��_t�%\�%�-����@�Y����%��OH��«����pax|�<5�̀�-E�	���u�f�AyfͳG�k����4�V�[�F>��d}yz_.<dR�m5��Ç�� �HFH��	ʵ��jK)�t���nګ�$ҋ��lPw�y�M���gxq}3H�X��}���4�:X�-WvcγFHQV)�����Տ����р�I��a��̥�����x$��YBC��+�]vٔd�S A���0�{�8�{��Qe�YRv��׋�:.�Gql{���ܺ�/�}C�eTQ���9��d���J��x]1Hhd"ve��v��g_�KKƤX���>���0f��&�K�0���n�E0��ܮ|gǰ���&��go�J���슨�����Fr�*r��|���?�%g�
D|Zs�8M�9���Qr�?XA��o����f�~wյ�~�Z:6X��{x�y�<|zrw iM��U�zy@28��� ���S��O%��q�#�*�|���`�e�W�eJ4�}|Wӎw!Âѵ �+d8)Ft��&8�˼��7.�FPi�l��l�K�?'_3�F���ٞp�#M3�E�Uj8$�'H���Ƚ�m|@6�,l%�H�7�=�V���{�8��6���V7�h�E�	E;�m����dW��:�M2a��l9��E�	O��G���e���g}�K8�n�	��7k�f1�Qi^�x�ܜ�D�~Q�ݹ��$:�Fl+�D=pӸ�J�*q������V(VW/����Հ ݢu�7q�tTR�@J�����t醃d!&��v�Wm�pp}V���W�����W�t-o��t�QF�G�h�n6��vC��;��$:K� C�"����H(���E36�����@�%�o)�ό���\�?WR�Ad�`#`a_Po��$7��?�+����U>ӛi����9J%��q~Q��O��k[�RP��xD�R��hQ�k<��q/����+�EV9�v���oO��\��&��툦�
�,�����n���_�>(�W���n�T*�TȦ$ ���j�Kt/�w&��Q �q�l��N4�}L����?�_8�yVf:���Q��<��I�Hb)�JǍ���:��,�Lk�$�^1�W5��4<�����^|�޹���v+�;_/�B�XG/pulI�o�v�	<������)���Yq0�"���ȷ���Įec���4��vag��yM$�C,���C��݅ട�����=(5�8:�8z�I&R�\@����m] ��VO����]���s���y�[�GfSV��d]��)~,���"��}5��|M:v#����/n{m��O�?�"4[G���龽��4Im�}5A'�x�S�ګ/+[y��5�WK��h��|D�\�;Cp��h%ĺ����8%��5C�����or�J�`�s��ze��Io̿��'5ks5�đ'*����DBЗ� �S�z�.�uݳ����f�IrƠc�6�*)�}n�"L�1�@[$7_df1��NwKz� F��?f��^��w
�:z�V��A%��)#�����h��hP��rzE,�?k̽���)%C�#�N�Oӛ.�IޙС>����+�� �'�:���2t���ԥilf�Yq���r0�ƻ)l���|mdL�@�yq-�>�z�k|��\p�(�L��)q0wh}�I��9�y��|iHE�t͢�����O`���@�ժx��K�r&MF��=Gd%0h�d*�l�����|:��v!=I�P�K�
�n�Bl��֌_B�DV]�bk�#�V�x!YS�W�ǎ��}	�tkZj�ۑ!�<Tv۳P=07O��4"���� u�V�ᬗ�}_Kk]ּ�wk��NӋ�1C�p��?�NS��6_WT��	|�]U�Tf3K�g��\��d�i�1���<\.6�|�@��ʻIv��!��@��#�:��jř�n΢�Nf���sbo��դ��I!����W�U͜�E�!����ō����,΁|!���I���G!߷�Q�����lԠ��*���&��U��3=?\K*�B��[�3�3-�}�����t쇃��:�j���>�C1��	�������?Uo��pa��=����cItߧ�ucn7zu��P��>{j���׈�x|��W�͗3���i��y?q0V�ܿIL��<8m_� I]T6��\��S���U��a"�s���Kk�ML'#�u������Wc��vÐ(��Σ�*�޻x�ow(;3W��ixmLB�e�s�M���b���p����2����N�r��U@��=oQ���^gb�(���ʀЎU�V��@�0�+WJ�D��o/X���,l ڎ�ips%s��d�|���G��`�x@���̗@�"=�hB�{�X��f�N�9��)���iw\R��T�;x&��7��@فn�[���W��Vw�ȴ���Ԧצ����l���!�)@	��⊴)���k6���Vm�Rd"�X�p�9��}o({���@��,T����S��W��X�����^"�ϴ��?$���P��Y
p�/ ]n��[�@5��F����K�O�#��`n�B��<���&�V�Z��u�:�2 �E�h^2`�*I��zv<����2��H�l?Вa7j)Y
��٪?�0�ZJ��v��� �c� 9�^��>��W���N�7���~�li\��?P��/��������Y���h��[x�h�z����}H����B�'�ڸ�D/�������d�����ވ���g`�H�4���$��1��"�$̟^!p���iˍ���oX��E��lv��<�^��]M,��lڒ������-�����Q4��0�U���WM�f;�_[���O�C�ko�TZ����k�Z�s�q>�؆��F��A�ឯ�l?��>O�g9n�ї҃Jȸ���|p��Bv,���iPD`�8��t͛�!��
��}1<I��߷0�S���kn?���u�	pL,3���P�ּ�'c�0�C͜�G8��Q��}a�Nv�(�n]��<��DW� �:��1���0c��X6[�0��&�a�y���m�H}�#�Y8�R̀Y��KipGS�S���OD~6��Y�}�i�H/o�ΚȎ�1v��ƾU��m�m��g�$�a��k8�l��t��%]mg|�1������ǌtC~��DɏL
zW�.����s%#A�]D��W��),�5e�c�ۜ�cI���M��&��zᓪ��K���ln�M�\��/̿=!~O���%�s�B靨X�{Np���HN���ő`>5<:�T���5�\��4�,k��B;o!D���A/�ߨ��-�= �o��$m.28���%��#z��O��&ױ(&�j��.<��'��}�&���t��/~'��f	��c ��8]�m�����0'�'F�O�Y�(�#t.�b�?'u���@s"�fӘ��m��}a�z�2NG{^�s`IdU=TA��p6��ǐ�16���7,�w͖f�k�l��.0_@��o0��Ų�'�90�4HxDH.�U@�C���