��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a����"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!���Dꁖ�0����/L+�	e7�n�g�ɥe���������/��6�5f��ފ�g2�H[�+�)�}>�2� 	��.�� |p:8AU~���H���WhV�Z���</݊A����`��׋w^u`��+�u	z�Į?�{_/�W"���|����R0�
���\���>�r�S��?go��?���7`�����LY!�K��3�~-���,c��	���6�(`�m:���T�(�e^+s�#=��b��C|���Ry4�*��e�j/N�ٰ�,9�$4�+&[s���>���r�+���Q�%�ƑW�/À�K��D�E��X���������^k��Q sv>���B�	QL�k�D����i��N���G�04Ƒ�P��>��_5s�72���S��ǿnW��Z��W|�x4�_��4��ֈќ�d�V��;q��/K@�|<�1I��0'��caӵ�>TP���'�^�I��A}5�%��t���YS�Z��S�+�/�kr��{nɤ-GFz�-�os�fB�\������l&{�	\�e;�p�%�8RI�E����e��Z'���)�`M���z�G��v�f@��.L�c)-q�aI���v�����"�T�q` ���zP���N6~�l$�Mԋ���,]��މ�����zH���{��(�7 ��o�����%����������Y�A$O��n+�d�I6&g%��3��� ��mae��bg�*�1��M��KDEPh��JL_DF�hg��G|�~��Y��U>�[!��fi\=t�������ﯳF�! �7���/�5�Hu��#7�R�lhͰ/�3�9�#fg���e+�;/�H3��8��#�1;�mR��`���Ʒ��"PT�� >A�OYZ��^�5Q��)(C3�pHo�G��m��TAI��=���pƹ���$���Mբ'3Y �� e\�е�b����>��{8U{1�H���Vx�1~Az^��5�a6�l���������'���`!��ie��N0H���,���|6�0>8G&=���ܼ�[�������XI�IY;�M��Y(�qڈ�ڞ�k1s�&�^fu7�K�C��0��i��V�l0E�V	�	6��_�ʩ��� ������+s���ݶ'5��?W���J�:�bÜ ��A6Ǿ���Y˜��cQr�IA���n�[�b9�D`c��ם5Pg��;�MPޚ1.���s����^���d�f!���
J���)a��{i�(��u(e��A]��I-Ő���z �'؜����MV7�Xsj���u�fU��.��0���	]PV���4�C1�^�c-���#���]�i_����7�)���q�����\9�ޛ�>�y �`�p����ELK�7�I��� ��\B���Q]��S c@NX~z'RM��k-�x~V/�O�����̏���-�$�!/���8h�����`9*e[���(-�+Ta�0� �w�dH(2ϿȖ�Y=d��>�X�Q�K�hxe��[���8��R���w���c3R�c�i�Q�(j�zI�"H���؉h
��]k+��l,4�Ey�y\��(�M������H$\�� z�R�`�E���8�6@�nz�Ğ/�m�l�E,�5�-�_�|�O jz�
�/S���Z���ĞF�Lv���7b:F�WP��ÿ^I쨃�S/K.�GR0�_є?UE��|� ��d9Tؘ��M!(��~�[&I���s;]�_��	>Ź�^�⠛��)�/S5������v�,OR'�^��4?�ގ�Z���8輋	0��ڷc��ڇ�cM���l���_rXT͡Օ
�����T]s�*[��V���.� ��[$�[��̿>�M�8. oآ��m^�\��o;�b�2p�����Q��\����)�9��m"+�긃�-\�J��/��~].�+����݈
,\��Ģ��ăv(�zX�z���w����4dPa���2��ك��y�m����O$��f�R�M__}Z��Ʋ�|��YB�,�y���<�t���dl��@6p7�4�:���R�8�!��eԮ�@�w��T3QT}s <#XH��k�R�O���չ�S�P!d�,�"��UZ�Jʴ3����63v3Meٝ��_v�&�f�@'Wm��l�av�j�0���p��
F�d�1�BR�?7�%��Q��N}�L���y,�M�'�<l`{��F#(ގj��[i�@\4]�Ƴ4�NyxX����r������[����S���41��"�vbyB��*�e�C��Â���U��v���Wx�F�����"�34q�c�WN҈�h~�gE�����O��G[��#�=*��o�;ߏV�	�I���X���`�����3	�����6�yQ�8���7�{Y�,/��M7�d^!��X����'�[A���5��A�!9ʌ�8/�/��Ҟ�����Y�����E��@�q������Zޥ���-��O��	CL�7~6�����3���#�;�)b�\M��@����@u����B\p�w0+خ�� �`�dfy�Ҧ5ַb���;�/���e/GI�t���;����`���D5���n�G5G�FD{Y�ؒ"� ({�X�P���v;&�k��xF��x�ѝ�������f5I�9D�ǥ��T��u	�b�����.I֍�]��llK�PnL�d����O�ާ��Mv=����n�� �{��y�x�_� bw�!�mN��� ������2�^o�9�Spqy� ��hE%�����,�oJ������/A��dk�I
�`�U~r�&f]��d�`���^�8(�}�j��ve�U$�L��z�}�\>��@. 6�Jn> ��T�MaSܤE�ӝ4�a�]ώ>|�P� �2su=-Q�->kD־�D���$��׌
�PͬS�@}V��AL.:Ͳ��u��?D�ogѓ�.mJM��(�uXo���+����k��n�,�x/L���W7H��A�R�.�+HL/H6��7���-�(*��v�Q¹|����'誨��[Q��g��A�#�M2�]W�N�(=.�dg��IY�G;<������V���[��Qpu3��~gg+���11Q��n���� �Ң�+M5���M*L���Zs�Xy�(�^z�t��J�_!$�&����L����)*pRp�kC��z� "xصkt��M��Q�ٓ��>��zb���:��N�-��w��r�o�Zge&���"�h�1'-�]��^k��2�x��PRC��L~@&�Z���ҹ�W�=٥�u�ƑpHp���@o��qll:���qA��5y)1i3`�-y.�pVW6rl�y(��^�col�\}*����[�qЗ˒T��.�	}��8�j��0�:Q���n��F[��e�5c�wx�$k͊A����|�p�1RMuaT���B�^����9���e�;p��ٶQ�h�.76�q�5Y��� ƭ����.K�{��s;a%q�z��m�<����kp�����z|�+�~��5�C�_C��M��mע�(!�ػ��Y����&�����tm5��	O��ɗQ����X=Q!) ���(��]JɫǷ�Fdm�tm�Xo�ݪ�)�$vi�H����
�Hr� �e��e;��V�x+p �K(��"/q�:���o b�l�*��%�4��@G*�������`��g�����/��N&����ޢ�b�xwO���K��P7G�}�m[ޅA���������œV�8t�C�|�ϝ�����y>d3�4KC_(��:q�b�y"�N�Y g��N��Q�	h����U�5}��ˉ��u���V�	n�u�˽7���9BO��=��������/!�`��J^變cm8G`OШ�fF� ���Od�v�l�(�۱��2i��G&�Ö���g�c�Du����4"8��ci!����x`;��V�{L6�-�hiy�J�7�
$~ol]�u���ӨG�@���([Q:u�6q���h�jژ�D���`�j�t���8�ۦX�-�X yrիP��B�%��O$��
��ڬ�)x��G�4�0�1`�����y;u�ZV�a��p�N �B`%�Mq�ǉ���@�~���1��;�G��P#ixZ�' odum�Δ�-T}ڧ��5劍��":$�����cD��U����Iλ�ɛ
�tQL����ؿ�/$A���Q���N���|�1an
=q�o��[�>p�:�q�T�I����ž��݁�9�Զҋ�a��d����	W�p���ɷ�H㩖�\VB_Au��xc�/� s
�h��ሠ���8s[�Qhf��_��KEfeC��w�l�W�/���N�{���Pے2)�!�{�{?��)�k��	����_,/����;D��b�~s� S�T{ڠ��H:���#գ3Z301�豬���a�8H�_��	h���u��i�^��N@�@mٸ����m�e�nm{N����"�iejצl^Bp�Z��M��m��U�A��]��Bmܼ�$�j�|mW�Q,��際�n/.����"%�lO��*�RO���׎�8Я���/���V��2����/W=w�B�i�Ut�snaG����Q�
�e�<'����aB���.�G�r�N�`�ǣn���{�#7R*���r�!ȩ����Dj]�D��[���_߾zr��2 �q[|�@��\����W�du�Onb���44�����(\k�o�i9$�e�*��4��YB."C՜!��IH�"0z_�龱)�Mn�ki=y��f��w�;��n�U)�.�.=�?PGP#TK��h~E�֟|xc�m���9ܑ^�HV�m�z��nX�Q��wG�d��hZe0�����Y��m����ި�nW^����f^��p~fPKv���w�ʤQ��=�$u���$p�*L��w�]�5��'q�'J�O��O�"��!�	�C���+�x��Gg\�&���k6v���ǘK���;�\�f���gA&�����^������p��N`uR��Dd[k�N��R>J�L�oGFb��mJ<��a8lh-Ld ����xcM-��תJ�[�&��r�Ś	o|���)�%+��_�Cǽ��]�z�y�!�]q�|�о�c5�	���^ֵ$T���	0�D[���7ݛj��b D��:�!��|V!�����y{�b���1�3C����<�.D�<G��w���L�����p��%�k���#�x�
�H&��e.� �����lU�7N��mT*�$�Ŕ�����l{�^�T��{_�Y���#8���"���o��n�|�jE����;�X�>���A�?n�ł��K��^�ƂSW9kP�;#^��[q�9����8��:�ދ���>i�+�}� ����'�Fn�7�1����f��5�Ô>���5�OӋ�@�o	�>��k��G�of"I~Q�n��:i�K�ؑ~�p�Q�i�.9�2a���̭;�Y�w���oj,�[e����^�y�O�;h+}ٓv�0$K��?m�\�(j��NF�p��Q#�s�.��!�/K�3�x�����E? ��䦴��WΓ.rѯ�� �y��9>��Y�D�s�a.g Tvށ�����������k"���h��jC�U��P��<z:�9͝���t���MV�>˙9U(ﶾ��j�#�:�%>�Q���e�B5���� ,��[�K���7Di�%(Fl(�H�}P��q��Q �ī��G�L�U�fRj�$~�-:�3�Ү� ���7�<lP���i;Y{�	���vZM��R�\��L���5��!Vܰ�^\� 6�kBR�xs�Ԧ�]U{g�d
�����!o2
���g(CD]Ku�5�����kY0J�D1�������s����:h�Te#��)���r�-��UC�LCJ��({<	v�+�h�-E�ӣmƫqC߼0��]CjJ�J��+���P_`�z7J���^����4��T��Q�K�]�ë�j�� �Ao��^%ux���:���z]��l}�b%9E[Z�**��g�lx#}y f�t�5R��e�󬍀I<����0���sI9�]��`��vw�L�T�WZr�轣� �8n��>�NI�@I�#ʹe@#~���ծ����B`��n�s&���6[�7�������ib�����$<��B\|gg���Q4�n���ێE�����W;ڙ�U��xNo�^C��G��Ԧ��ų���Z����Ց�;Nv���|�[M:�j�읐_�"=�:«�5nv�u�ƹ��V�M����o��\pm�i���"ǔ���+�A!׾
韉�-l�|
Il
jV�����^o��+��ၡ~^C
H<:���4�V>߹u=%�ղo���X�7��v�me�1�*O���&�[�&�C�����((�j�`��v�&��P�7JS����W�!�Z���h~�Εh���՘Y�Fl72S�f��m����=d?�5��u���U��fH
kݲ���7��h�潿�CX�D�nQ ��m�2W���E�|6s�o=�b�93]8�K�Zn�<����k��Q���,����[W؞�qOv�~��mP��y���;p�3'�u������ߏ��M�1��S���ȯ#�j����;���e �j�5:F�U�� ���r���I�w%�r��
rL����]O�^�	 G��3���7�-M��'MUĖnbz�&���z���������8>�y��� �Ȇ[�>�j�O�ƐZK���i?��ud��BWRm��B�� �.^��0�rDPeX�F�4˵9��ru&��S�a��D�!�9[p��ԴG:$�Z��ܵ�͙�i�ǅT�$���SK![���q����p�)�4
���_x�=$>�u����z�j  p�\�w2gmA��~�4�kX�K���.�x��|ϓK
ѽ5��_R�&�8��ݬ���Jh�����c���1B@���%���J=��<�I��#��f��7��]��lE� ��,]��/�e�a��wQ��u��+�[Ô#e���lRq5���"l���W�i5�� cr�&�H���R4�/�2��ݚ�h�OG���q��3g**����M�,����s����^2k-2�'��=h~�x�2ãbTy�
S��je"�⩶��p��ro�4{!1����7�p{?�!�:ou��`��g9��0&�����8���qI5��v�)����?��5kD�a:�Sx��f�Etqv���2k&<i���k��7�U��,�Tb;� �rOTevI��z�@c���Ґ���-�������>:���.6>*ճ$��yM�`-��~��T�!1�ݸ��vV��c��I(��Z��R2#�ݵ�^5�[2���]!LQ�!Py�m�I�~.s=�/��n6f�����'��Z�?�xB�lM�����M����b��L�{XN���ʻ�Fٗ�+!�0Vc���q$\a�������;�%�:Hlp(o� 4΃�y�]�ZF:x�t8+���9�>c��h�fM+;���4�o���~��J����S�	'��^���'��z>����^���_�]n�WDܯ
�M�i�8��&Vʦ'�I�ʨE�,�͎O��r�*�.�L�}zt��'wCXD��:�ϙA�%��gKjkF8^n��ۏRd����m���~�_��h�z=�e��Y� "�71\�~�ݚ�;����b6���ժ�����P��_jl��� �҆����d����3Sr����
UDC��JGI�w�#[n��2��.��/{��E�"rcY��ԹA`���9BM��l��
��69�����:c�Î��C�pC������:�h$����/GΜ<��a��^�bP��&0{��+s��.��N�� ��rp�`���&D-�&Y��',�]���9t��Ǒf8�����{y����=��q��`�ɓ1l\�Ti|�녈�h�}[P�Y���r1�C�#�ofl'��u<����<��-7���*K�3
�����je:INYzcY�چj�Q`c~}i�(�V�˲E*$���$�=��#T�|u	.����_�'K��A'fU�p�����
�ͨ�G��
�w`�Oy���Kj�b �t�MS�[ҹ*�&od%�=���2��}����R{�&�i�/�X���>��:n�q��s�;K�,���מY��h��>]b�oe�[G}9W۫Qu"�O�^YA 6AUMA��Ido���̒uTa�I�)��ÿD�u�-lU/�['�:��J��"�Qww��N�|���@����r�}P!;0�o�.��G�.M�C�Ѯ��AGڍ��4R��nwf�>���D].��5���5�<I�����ʂp��H�MB(���=/�#{W�-�y%ƿ
ů=rfؤ����au1�U�c�7f4��]z=9}�������-dd�zO�#��)h*,4'�DF�������Ӕ���ێ�͗�������P񠺌��2�,x��r��֓�LcwE�c�����W^yz�c��`H͙�v�Vm�*Fg�0,��^�S��i7G��h�bn�zvu��!D�g�4��щ��Kru��i�Y�*^'��]�`C���x���i0%e����ʽ�������1��v�G��@ȿe%�lFuI/.�'�Բ�������AV_�&�"�����}��N�����+��^zTȎ�dN�=���n�Ŝ������
�\/��np3`�U�Ϗߒc=+$V*6e\R�z�(RB��2:�xH��>������o�"��Xj+et�~N6r��n��?,{~7����E'4o1pW� ��4��aq��A������8t�eNH���za���[���7r3�%���8�8��@:����VAA�A��U	�l� �*B��j#Sl�b��2\;eO`�:��V�kE�}Hλ���g3�߻�y��K�>� ���$q����X� ���Ƿ)m�SԴa_~�3S�ډX��IkU��?���?3��� ��O��8���bs��W��U��l@!��J�&↱���̼�MJWK{v���H�Ǚ���c���CEʺc�WH��(j�"��w�!��:d�d�;*�r(��/WFϬ�TS����8?A���.�X�]�b�:����K:��́�����0#ۗ����L 	���.Z��09�>�~�F7�����~�37 q����6	߱vK(������@���-���Ԯ-��0�-��O�<�1�f��l�}�����W��l%��M?�l��~����l/Ҡ�Ľ_���@�x�{�eÀ<(^I�cƓ�g�l�ǭ9x���S�_��e���l�=�:���X*�p4�l�!z���6�Y �cD��|\�S�1�8cZ�7ﳾ�@%id7����ġq}ɴ���:�ź�=�B��'"k�U!�B����:2a�au�����u*3ZL�:��W�?�;���������]fK�&�rDr��J�����'~D���3����CGA���3�[���w	��h^���%�7+��u	s�A�ab�r��y>�f<�ń���Pc���;h���"�ˬ=�v�ƈA� ��2�uwawTq��>Ю&��n�w�i�z�pAݮ�7,)f��0m>�B��Vr��x�������H�D�;�u�vȆ��^�2�� ���7)6MI�?��x�����A�Fx2��պ��GD���}{��nyF���u�r<S8wU��wMZ�2zX�<�UBUh�R��hZ!�n�܏O.�A:��D>K*`'@c��I[|��=�V��{�{v\�y��[��պ��6r �umY
�};���?�ľ��cy��?whEng�BY_A��(P��pu��jN=��G��#�8��>�ߴ��Q�=�};��D.E��f�C���Ue���Dq]�iQ'_����Гdi���j*�����1����<�%�TC�/t%T�w%<�D"F� ����٤���T�_Qy������A��W�ŋ�5T8���j��M��K��� �D\���>�-+*H��B
�oQ�6"��R�_7]��!9=����z|�)��ϊ��pMN/{��AUd�gb����V��g��>mQ����FR9YВ����~i|t�K��|�k��\w���'���V-��3�޷�@��,���x�����v�&�3�*��قx�g_
�����/W����q��ώg' �v�l<h�5P�9�	��s�cl#P �9���쉥S#����aYR]H*'*Bu��3�hȎsn����MD��QC�O��.��������oH�d�p�J� ρ��	T�Z�(����!G�7�5�A�}��jע���	;������T���[�"��(����'"x�ŋ&��q���,�\����r�b-sqɄ`,���R܎�cX���%"U9�Yz�6N�8t�B�Fiw>�����
�=CiS��udy�*[d��ْ!l���t��t�7\��R�G�PB�UZ?���>(�6۝�ac1�+g�2kAafeTΥ�cu{Ƶy��'8�h���{�X���ѡ)�m���3��%$D!��R�0��!o�u���J`U�T,�2P����-���Hkauݽ(��7U���N��fpSG�[�_xjČD�?G9u$�V�L��^����M���zʰ&��׌v�*��	��b��ʩT�\q�X��!*r�X��0��5p�v��]�3e��I_꒚3���JR��LiKr@u��نł�}q�QXJ���D] �;�RPN�N�����|+ra��~}����E�.���
���Ǥ�*����<jVt�3����Չ�f� �Cgd�~��`��l�����kO�%����"�8a�`�݄�&r:�78a1��y��$����撃4*�iLaYT�Iղ�K:j{��׀�>�\Ѹ����̢5���f�����L���A� �:I����A�� �۟t�aӵ�p��h|Ӭ��+i��ft�0����}I�I��(LO�&����c�Iy�xJ��J-.��ĵ'[��?o^�B���/=R�kVX���z7������',�>�����	�����9��	=�ԐT1޲3a_t>�	G�0���#��{՗n�����;���ͭ��Pv�O��B��}T$v������1��֘�����F3�����P�c!��p�eM&��RM��i�!eui����_B�rEX����:�kQL�x�c"3�u+Y�\'�tJ<̓u�>j+b-�w
اR���-[:���k9���8�t2w�e�q��rݚ� � �C��ڗkOu_��л?+�4&����~vR���*��+L
�k(��2>#ʐ.O��v���ָd#����UVc;T��q(�}�`�l�GDw�������N�nӘ����qT��1	��X�eP8�^%y��`5T�9	�\���Ƌ:�*;�$ ��DϜ�H�{�Զ���d2�8��?��o���%7=�[��u���p�"b~�+�B�`�W	AɊ
���"���kyK�j@D�ލ�֤,&ʶ�˒�L%��#��3|�W�N�$�4��oI��Bg�����9�[���]��V���/�L�#~ɷ�<�����_=��Qd�\fm�H\P���Pʣ9DCs ]��o�XW�ZV5�{�9�A	=y�FX�ņU�ϊ�HDe�]<�Js���Z��sG8��{=ث�M[� �&�X���Z���)��^LQpʭ�o&�#UgA,p�Q�Y�����!�����8����/�4KA���L����I8�R%b=�:�5 ��M���m@����f�,��6�E�>�ŴBo���,�Զ��&`�-W��i�)i�Z��:�~�>bZyRG���O:ǥQ�.��im�A���-��D�J���_�q.�����S��fl����.�4}�@�Y���&`,�����B�gmNX�D0xGx���� �\8˟&�/^��u��&�hp.�A�|�a ���(?YZ�N=�bT\Z�q�W-0R\��<Є��_w4(0��P�A8|E��v�K�G��/eC��D�����^�"-)����90����n�_@��f���=n۽�7Cnċ�C�^��:c�c�L��D�L٘����d5�"g�=�L�'�A���dӟ`ۿ��W��=UoB?Ҩ���z�E�����]RiK��F �!Ļ+��W@���쭮X�M��d�D�O��y�p�ݪ�c$�Y��Z��<�����֑6��*�Rԋ�_�7�=�{:_�|{�"vqbm2���c<q:L�}�5��m5Mi-y������tO��b��oi�
N['��K�D�I����x9_�(�'�Hj$����è�kb?��$�1}E����^:��܁�֕_y�u&?�Kk�u��R�J�34�"c�ݺ���2�ϧ1{�� �v*�:,�����IN�I�{?�+~Ɔ�u��c�� ba$�zI0��*�DK3�gl]�+G!C<%(�p������nE����4u����D<�zҝ�>�8M���O>Et �A�� Gy���9��
�ҍاm���WT�,��7.�O�q��ϟĪ�ei�O�hWa��镅� �v�{?�^�%�����(�Sm�$y�w:��u.'K�Ѭ��v�D�BPnGd?Ff���>Xn<Ϣ�N�g4��h$��n}ѻ7�R��ƃ#�8�+���+��6P����e�r�A:���]t ��(�O+����B������Q,�ъ�y##"[:pf���ش��~�&��������ኪ��
�(�<h��d��]�@�&׺A���;��U�XH�V�4����U�L%6Q�آ�ֳj�c���q���r�����nu��ȃ�T�	ku{$����t�&6A��ĝ����R��rxř?/�-g�Ƕ:p=D����Ϸ�lթ*)q����AP�Q���	������6�:~C{�C�^����i5�cF��C����'#$��A��>���86�R���b<�D	�1Fj;��#���H|/�^Dz������ђ!�>�.H_:�h�9l��k����}xu��s>-�_F+)��nh�{�Xoj��Rk5lh�-�׶4�mT��1k(�M{�k��v���:���l��6�`��2)�1�D{yk>j�A��]"�( �a痘bj�I�S ��_�+zK(X��ي�xZ���*�3mY������W�hΆ�W���u��1Hp3�zk?~��s�JX �d\1���҂w�
2� ��
�� _�'��ܜ�d�,���ҙQA�A:j�����pl"�w�����tp��ޙ�-?��x:Y6&y�O�PY�p��c�Ǹ.ta�A@(�-9�2�;�w�`��<�w���9
D�HKV�sp�|R�;�z�*�謼:����" ��4A��u��ys���B���.w����8`��?�����;��/ta����T�,����Ű�Y���`X���<��4VD��mF>�J�;��� �čb{�=`��C�����e�YW�	����ʓ܊U��6ב�7`1Η�j��l����T9���b0���:l����LJ�h	7���=��?���TN1҅gMRyr�s�<��R���h���=.��%j�h��X��Af�E�qE����!3���?&�y��7'�S�5)����]�$bɆ���s����iܛ�*D�촸T^�둜sh~� ��;�k��Z7���f#�K�̕��F���ry�.�H�J4�A�Nk��Yt��@I�
-��~�8���A�t1��S��p�A|�K�����	�sGA֏q�~+rݵ�BBcQ�JK&E��tvh�'ڤS@ l�s-����u��P0؅�U�4d�}�6�߶�Sv���M�ɭ1�<��w��D"¯�������� [v�f(msK?O;c�!�	�'��Z`����������J�`oiX�7چK�C���)#�z�u������F�J|6�1�h��sZ-��(��*���	�S���N=��Y���*$9?�������r�+�!���|�ӮP7
;u��שֻksc�Rcn^1[9��8Ĥ�(�p�f�,�
��� Ƃ�j�n�.F��q��a��WE6L��)�o�l�l>��ZAkB>	�zo����/�/�S״���,;�B���	��z�L�և�� ꮰ8y���Ug����ő�}a%�a���Q��=�Ӵذn�s�Wv�[���J�Z�f��ӂR�:�>��<9t�ŔB:J�X]���.߻������*�Sʾ��`C���j����d��'�_6�i�_g��&�
,�J����1L����#G?�:�#J+��X��zW�V���zBJ��zw�\#��71j�KX���3�T�@Y�a������1D��w8�����D�� �1a������]�ꍄM>B����}#D�td]�����_�\-��q��h����=z�`�����J2*�w�=����j���݇dd[}rI`����|�����������T�״�ח\��>�܍�E�Q���[��\8��:%��ӏVg�%�V��`���mH�mk4}H��N^�ſ����n__}�Ch�����#�W��ޝL��qp��m�3�t���uX_)'�C䪋��s�?��~��g�_"O��P������A=,�����L�d�# GQo���?'"�W�+���FǬ�c�G�����������L���
�"oD,�|۸������*$���X4 ��S��س$ X#�"��jwAp��_T���E��@CH�V�R8�)-x�	S�Pa���6���q'}�OS�&�e6P0��V�����tTJ��#&��ƻ阐Yc�;X��8c�md�>+����N��2����B�(��!OqW��:�|���i�	!0�F�r��Z�ڹ`5����ڄ�(xB�@(�]� �b�͡��s4�ź������p"�l�@����E��
��V2�Uy;��8ׂ�w���s��6�uIt*SYe��8K>7��z������LA6NC
���]9��0�b�fa^U���L;w�b[��I��^6���x��@�?�ÐK!�%�W��(wQ�Q8�DC�����1�#l}}`tJ�OXE��g�݈r�;e������8�D�
e��I�E�<E�H��o9���y�{'�<�������Ϩ�N�K�v��J�B������v�=t�=z�@�C�"�Y�x�Hx��̬�B>V�ȴBg)�dͺ�m�le�k�3 �Zp
?����B�~���D����u̸�d��`��p��CBM�Ѵ`JA���9m�����d8Q�f�����~xy��ߦg���俺�=�2���цb�	}��5y�S�cKJ�f?�0V���O=�߅F�4�x��]@:hv��ڑ�o�t��{�ٚ��[g�VBŜ"Yď)w%`�
�l���ZuFK���&�� �uEϘf�HC�!�樓_I���wZ�]:�����n)�~Ⱦ0Pjcb��?�%�Y'�"R��`RT�d6z����tmiw9n�C��6@/���Wk�I��Z�R�@��;e7�A������ص�,?�j��Rċ?s׀i:�#�dI��H��g���
��a�ꕎ�
�(�<�2��	��[�	��뿱��Ԑ���1�C�O�H��V)��M�T-�;m(�B�d�a|#��T��6�5�OS��Z��cc�ү%��z^�cM�f� ��('�*�.��0w�qȕJ��L�&�腘m^:M��w�6)��tU�V Ȧ�ƿx7����h^S���H-�ʝm�`|Ӏ���X�K��=U�M,�@�0Q��n���t��d���+k��$���6��o�M��3^=��V<����t���t���m�Aw���R���v��>���$`u��8a8EC�F6��p�&�78>���k�k?ľ���Y\y&wn#9�Hk�2�p��J�,�N3t����N&�)Ɔ^}�}����v��z��Cf��3న���:�3T����l��`;�=�hQ ����0o]�7��u`��6Wp�� �霎]��~�� ���	�,-�ʡE����tҸQ?�v�(��r�u��f�;l���ʂ$ې�D�q���(�C��\c\�(��2!5��<�4���M�8Q��M��D�+�+l�픢5�i�vˠB�2���jv�q^��Y�zP�[U�f
vc�F����,����|�	�P�$� �g�� ���r�>�A|�i$8|�A�*{%��Oʇ/�)+Ļ��Bz��"��}2�zL�Y�V�����.���G�/�Ҹ��Qive�.�2� ���DHx�4Gv���wpE�� lrV�Uaj�g�U�;�;L^��m�;j����t-"*z)��cڜ_t�i��l���ml���a�v�o�)F>GP�k�ڙ,�/�{f���*���ђ�� }>l�\�Yp�G��O��q�'�sau�6�_��o+���Q���%T�C���y9  Z4��M�yu�v�˄��z��4w�B��M�9b{H�7H�'�ɟ���uZ0]J?���A�`��X�"�q�n�J�f.�_������θ�q���Y�o�:��Ջ��Ͳ	�a��UM��Fj��(2���lŷ!'/Ҙh�/M|���vug�6�V7>��?�3�P����a�s�&m3�c��6��c�;�I��êu�֓(��o�}bzxh$Ł F��q�i��_鮞;B�M0��3ήqB�����{��΁����~`�bs�v�xkq;���'��jUܗH�*X�؄�������:���`�Q�h�y������t3FUv�E�ؿlזq���	��xRo��ٳC�q��dG�R`��1?b�&�fX��}S�Ĭ��7dIJG���Y+�IlB�]+)�t圼::%%��RɅ%����+�pA�ID3pNkx�ᮺa ��^Q�+=����(A�yO'��E���d�`����_�b�	cn� c�;�2?����S^��� r��t3=����J�[�Ҏ�6!0�lc#�3����p��� �[xL���G�%�|M ��@�A��S���BC�g�5-�0�ƿ�$S���B
�p�yv7d$zgoo����k�J�O�bTPN �#S�� ѓ�8�R�k��%}_��[\�+�1��h>Ӵ)ԗp��ev2-����=yJ3��3��i�PsBs��1��Q����"���N�7�+êN3|O�C�hT|ېG�" �M�
�l�~ɄM�V��z���� � R�&�lC	sKQV��O3��r)��؃cȽ��m�,�<ԡ���M"~T�4�O ^��T�d
���qW��v�D*�v�5sRň�m��;SD�Jw^�X�.e�,za,#.�Faߧ�];��$�
 ���'�g��ލ�����G���ּ%�L	�6��A߹�i�bK�P��#�뒃n��m��Y�a24ά�7c�7�
�3�VR��1yYs��M������> p'�z�E����u8��&�ڦ�l������@�`���(K8���)*����b�lZQ=FJ�$ݲ�CX0�&<�5�Ro��V���2���E�!�9���U���RN1�l !=S���ԯ�A���g�vNn�r�|��U�ݧ�h5,=J����Z%��},�c���F�1�ɖ������ɝ�C�+0�z�r�_�y�4 �o�L�׶�;SV�"N����H��ޔ��5�]2�������&Iw�������*��= L#��B"vP���.�Y/�K��i�6Q8en��ԬO!_��~���Ǖ�6���������1K��(	��<H�G�n�Y��owJ!�ʂ��Nk
�[Q��D����E���h���rB�i���/6�-}��T��#�"f^i��S�*/����KZ��.g����Br�����B��o�d��BalyPa���@�>TM��T3+�o�ө��O�'�#�Mt���h�+[0;J�m��E2щ��v�|� ����5�!R@�#�1K�g�Eh4����eo��'!)F��U�kDCIR�twig-�-��@��s%,~Å��FZBm�}N��/�bY|[V�nK�|m��-u��Q_�]�����u0\LR2q]�4_��p��F7��cL���C޲���`���#�a�>����g/���"![�@`���6@�t	��v*?��BV� �5�yh���r,�LT]Z:��\�@	����U,��*ܟ�L5�!sy����\Z�S�dZ��P�f��a�ZBhj�(�k��.��홊,��cW~�)/�yb58�J��b�TG�ִ�w$��	 x�3
���~�}LIi7/h�IH��(0�iE��.�e�Ay눂�{����+[�<N��;ƿ��$�{���]�A�Y18��
�a�U�O����� 9,/�N�T~k/�J�j���|�d�a���l���շ�>�y��<Zt��&����Ċ$-!p*ZKl��U�O:�!����7��4?8�R�W/���������d����p�����Ojy��i��ǖz��m��{�c_Pm�+�v�~0�ݺg.�7(u��>��]�#��ء>4�춠~�0Fwa����Ȣ�������E�� ����}$wi~��� y!�1�`0�[F>j���j��]r!�5�b���s�3uE)($;���]J�ϩY-)R���ܨGC%o+�S�?4�������9Э��l�bC�&�9(y���"��O`�c2Xd�P\�	�ƭ���w�����T̛��8��@G�7�?��>�w]Wbg���6m�#_"'���{��*c8dSg�uD�FP�v�v�Ć9R$x\�9�S^�xm�.l���h<���Ɇ���᧎��C�8�{W�N���G0NĠ��Օ�Y��	Ž��ې�
�b�Y�K'�|���	��)�4@CN�������c=�:�\��5L�~��ю=��ھ�h�[�"�`�C/������K�)ۼ72���
/>=����MR��,��#'E��~�5M�{�p�#��*�M�y�<���Ms�'I6jTRpżj�6GR���2]��n����"g��C�����4/��s�I�)�6x�����]������uU(��_��-N
1�G��h������{g�3�!	�f��KJ]�{E=ڛ�+`�h�沄P�9)�h���1ȸ�� ��/#c�����D�G �X;�"�]]�2|֝b�)��Dޒp�7�9��MN����.f�����B�6+���a���WL�[�搁�ߥ�j�(���	�2����
�����w��� v��H:�B�!�1�e7D��"�}�(�/��p��ʻ<��2�M��0���e��%Ԃ������&g@+�����T:�w�W�v��טPƭ�gTjY��m?%�	�d����T;���7�$&<o+�p'��p���=���Z�Ԅ�1�o�C�𧼝�z{�Vk�C��[Eb-Aa�%1�KCHFx����<x�$@���0�oC�ɨ���mmC�#�I|�����y�;��h�\��%:�� �%���lѹ.�/cM
sf7�
���/�������xѵyaK��|�i��~9�ūm����֫� ,�W�q�w�{~1�_� �32�0�ȫ�N@���N�����o@����xC�F�\yR�[�{�,�>U$�~�CB�q�#ILo0����V��~�Oĭcw�Gm{��R2�n7��A��l��l��	x~�6r ���F�tX������w7���Euѷ����mȪ��K�Hә90 �	�Py4Ygl�U9�D}��K�g���Ad�U�hY����[{�a\&uA�n��]�r]8��4I-�G�`�<��v}��14yD�}B��C�P�4�"M-�bn_Y��9to�D��Hڰi�`~|�D�q�]X�+ 7�a_��h+��M<%<���A�H;Da+�_���Pߜ�����ۦ9D܀L�f-�6�w���e~Ӊ9l%��&��
fc��|��r���-��s��,=��Mp���.,���(�2��Wo��u�����|�g�[�#�wA֎�O:�2����T?��65�r�I���3������9V�	�p�?��~7Ҟq���ڕ��ou�B��g� &.��#�Z�yʨ�ǀ�z��.���P1)��.�X���%�_3Hk�p��Q�k̸,��t���],YA�˔���7?u��Z"[م������9�`��^��s��vi2���ϟ��?�N����Г�@]��xU�����Yu|\�x2�d��
v�4��U�s��WmU�&�11�� ���n �R�X�WD���ۏ�ey��v\�v&����l
]�������`��S�?�ǰ4�1[���CEQ�q�-��:lzܭ]���3UgM�J��q�U@Ԝ��7�ލ�^�
ǗX�|p| 4�L����`�"�V�"����a���=D�q��o������&�+ƛ_�T�vO�r�s0�����]� �F긕�c�|6��3kt���\��z�!l���a�CT!�$a�l�&$���~�}���l6t���J0D�z��/\��