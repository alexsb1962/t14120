��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5����Z�Q�!�&��^�����'Fdf}uQ��z����*��>1���	��k.A_wa���Dky�G�#�,��*W(<�����%����۲Ȇ�������J0i�}6(�� ?Rvt�=�8{����dR��冖�kx�BZ{��$̐�,�?AvvR]5�Sڔ�\�4����j��>,�5>�-������E=���Q b���k��s ������c��Y��E�̒;�[����5������A�k�R�U+IM�"�JGp��w��Q*�|H��2�c�o��MP��P�W�-�0����9�Y�� �~~'A�wёO��/�ϧ{%+�)�8�B�F�H��l@.��Z��!;OJ�R	(� ��P���P�C���^���J�yӵ�����)7�ߦ/�L�������vO5ك?8=� �$N,�N����C|��(��-����l0M��Hs~��d�#:/ ����HjAEMi���~������1d;�m	��ԢvO�|��H�R���v�ta��;��j-������6�,�Fj�Ͽ��9�Q���T>*���	��B�\w��������!*E	f�z���݉�8̬\	�v�ܥ�Bf��PO5d�9|�.��e�E�]��/��F@ķ[��՞�Ƥ���RXYb̹�}�4c�:{�U�m	���	^�.���o]b��BZ��E��V0��+���R
��6��������פ���N͛"��O��	��F�Z!ޢ���Iȃ���B���0� �����J�T�2nu�2�M�)�!ł�n Ŷ��t���t�����M(��'�sg���g�]j�z�ɿ�e�얱g?ջƝA��Z��Y�4�d�]�"1�l1�����:�Br���4�d��7��C>����^��N
�7��{�����e���s�����1		#5Ȃ����o�����(B|#ӑ���{�I�~�_��U�X~f�����p-�4�%���Q-�Q}gp���c^�]w�ܶ&쩜Q��X�E�4�r�^�1��Gc���dqƦ;���To涊�0�3�@����\gr�xy�&:�W�6!6���!7��Mk��U6���.��c$J�GMW|�*��C���Cꨛg�#P��!\hdii�i�\�!8���Y�t?�f=�Օ +�-��*�4j���鋽�Bɓ�o�y���D��Gz�cʕ��%z�O����q�~�@:�z_��
���n����!�:yh*�TY��Q~`�>��͙��z	?�����;��< m��V�A�������+^���g}�G|�M��~EJ?۴6��ݹȕ�8���{��0T
A01�'��z��K:����V�@ ��F�T�!`�M���?�Á��[q����@�ޔ����*�h��5n�'3n@�<#�V�����-�x�Ҳ�wYoq&.	�rΰ��|y����L���T!�{B[�'G ��}S .	2���ӝm˔5��,Gv��LrZ���+��谺9�ﮁ��֜�탺�l��	�L8�,�����Csɩ����ql,n�&���/9��f��G�����e��F��ז�,ݽX����]?ʾ���m{Q�t�t�>��-kMAY�\/͔�2����Ő��86� ��	c	�y[p.��h�$��x��E<�ݴ�_�o��q(�E^V�f��M�ĀH]�k]!�@.">S��4�S֠�k� �<�+��Z�[�Sr��#�}C?	b �����@�!�	$ԟ����^VÒ�+�s娣�����P�m�'����v�^%�JB3��7��^Δ>܂֪Z�����G�}�1ٝ7Jf��̟N�����^�@7m��i���X��kb�!G�Z3"��f�H�y	�))~�2fl]���YTUhS�%&LӲ�	Ii���n߾Lmv���9Z�>�e$_���>~��yHi��s7��Mr�S�~���_9�2b�����s\���˳������n
-��t�+�& ����o�Z�<r�n^������bV��2�.�\&�`���(Ѹ�4�+U v;��N���n&	����H�N���� a	y���r�,CD��&��QC���uڧ�K{v���d�j�n6K���t�$�t��f�������~F����}}{�S�L�	B^~t�A�u���oYv���t����O�cla��o�;�B�����Ɋ,�����SK�����7jT��.+�G���2�>V>$"�e��k
]�����H��M+ؕ-��t��rd�������.��E6���x/q��W�s|B2�_��NGrU��'���_����Ϫ�`-XFP��d�X!�-�aa�p�k�ۑ�gA=� �_A���)��F�Ǧ+W9ԯ�G�Zo���m�!@�b�儿dy�!A�������18��������4��v~].�=ɉζ5>����/2�	0����ך���Qv���U��@�P�M[�(f�aBNh\������<���D�Q��]�`uE�l�B�(�_c�V��1�I���Y��0��[;&F�Uܡ�������BM 5�G��qZ�&���K���u�U��PIhF��w�i���'���p��!�)VX�	��c�v�E�Y�.I��I����w��3Mk\��g4{b����siǗ��,{����Aзz�&�t�m���KX�B���[���eYE�?�l5q2"���쩕Օ*9��HՏhn!d����S��c��p+�A��,�o��Q����6zP1���\��q��]��!f�b��n�()?��HY�T��k`��,3GϵM^�4Nf�\�)��Ndu)<��ˢ�~zS�ӵ��s"J�ؐj!E
�p�M\;3FN��iX�㥈��iCR��#�HwP[Ō�
�a����d�e!?�T�!l�"$���3��0�Q�,K���+�6���<�,An�P�o��PF�,��K��GP�~�SR��S��\
��qk�Y�y��VQ����\���ߵ��&[��w���wG�}*���Ei����,4���1�''ƥ_@3�
�ju;|�$h�g���u�^$t������6����O�֗�r�@�Ie����#0A�Qc\*����&ۡ	��E�=t�,J�7�dV��� �J���y��o��ԝ.��FN��T�)�9Q�P%�Z)�C|~��P<Q�r1�ps���XlJ򄺧�C�eD�pn~�`[�t���Y��ɗy��K�{h������BD?�V
	ǹ*)�+H�#Y�
ص���ѩ,sl�|ܕ��c�7�NAQ�&��R�Ы�h-���= ����b�j�C����s��6����U���R�ՠ����z�-�����Ի\q�2CEն5F� �o��0?��F���ˇ[�(�Cv��jre�n���r�ֵ̙���j�q�rn�ݣUA��P�����G\k�4r"��(�h��c�lo���ٝUр�.�A��Ҧ	�qc���˜����Rr��p�^��s�z����6\�!��ơXOq�9cU��# ���<D��
ffM��␘�����"X�z{V|��e�nt��{��z��7��!�Wd��&<��A�yDĜ�4�i��7.\��	'��VО�Y �\��k������F?�ϋ9������J'�ϰ�u��k�"��]D�q!}i���L���6!qy&���d'���������?J,�`V�[��v��&F&)#�Zy0"܏a�����f㊳��Cb���}����)y��`P)Bo
�%���e`磽
���OI��p�_��<03l�y�����s�Lo�cTpwa�����SO��_����x��	���Q�d��)M��ۑ�O-Z�$%v�|�:��I�;���L{�6?>(��a���lv6;ʺ.�����!�&pDsk������r\��L�f]���KF�+6� lI-$/�q��`1�-�Wmt��)�9�
�E�ʷ�ǅ-Pp�e��q��z�=^�6���P�Yb`I�0����}KXR&:�ެb͔�I�I`�?�T�񹵝+�c}�A��kH�|N��%H��
������|����g`ue�qBP �B8 ��o^2z��ŋ��ٛ�����vo�$2�΢���lW�V_�^���	�Y��c�K�BG�*��ˆ!�,aB7�<����v�d����sb�f}k
b=�y�v���W�ٷ9w�� �~{��B�fX�x�I�M�W�L����xy�������������MU�1�EZ��W���Ɇ����a��Y�p�[)7qCے(����d���x��{h$e�繳*�IQ�i�4�C�m`�ou&z�[�,�f6aF��s7���mL���u5�H���8Bx+gxe{ n�R��ѮT�;�e2��!3���n�Ƽg%~�<Ĳe_]&�L3�$6��y@*���9����WX�3�^���q���W��Ei�4
 .��A����s����W�(f��} ��Zn,����.M���"�2+/!�N^T(<�Dg8f@k���Y}��m@�T9�lH-z����#����4�g{fw$�&H8�1�:�y�K�����@��Q�����X���8n���#*Ym�
A��L���i~�� �&�	9�i4���<}���y���jHGc���P�∄E��QO�v����|/3���'����������fה~��ۮ�E���qe�r6u�DnNT�G���������z-���#�h�-\.�x7��/y�-�y�#Vy�cn�X\aN-<���׺K΍�����#�rl�ĉk��;V3�*�YF\VI���((���]�ܲu���O�82�Uk�{�����F̒ *��w�<4�\�u����K�f1𚵤�/�	5$�^������g�v��d^�o E�0�rʴ���dXѮ%��^���LU�-"�^8�u��mFL���>��!�:3��o�כ{#�W�i�	���4s�dB��B���o�#F�%LiM���P�o��>�Z��e���&����4�SG�8KJ�z�|Tf�2��0o{�Qo�f�����Z���iA�tj���Bψ�),7۹
�k�pֶEv��I?��a9:�~L���3'I��vO�[!}-������o����0�,�~��d2KFpngK��;�\9u�6��p ��g�#�rv�����HH�I��������#f��a��d:5o{���Cl[��I��eI�x7'��,��\wA/� ��x���j^��
�M�M~
a���W�ݯ��z����>����s��@[0�h�Fb�ti�����sl��e��))i�Z)�*�����H`�n�fb��S?���b�?�-�)s�CDx��cs��^y�&��k� I�='�1msk����,����c��HŞF0Sx���6_���|���P*C�k�4
����o�m�)�.)�K{͐zڈ���L��ݬ��OJ�_��4̭�ʂ������5&�u?���A�Y9!]�����/IW}D����`洈3�PfE({W�*x������C�R��gת8O�
��$�ˌ�?i���� �p�dIE�SJ�͸3��z.��	GCj��wA������z�T�������2P������<\���R0$nQO�s�����X&޽�u;��e�P%U�����\u6�����K(�R�o\^V.X���o��Y�V'1�(Ѳ��JH�>��P|����#Ab)���r`���{-`��S��uW}�Q���'ksq������ՙ��s��sa)�'͗=��B*��B.�Ǫ�v{=�j��T�Ob@��r�����Σ���Y�'�vȣ�� 	�OY;�@�-Ͳ�乊2�N'����U�K&��a��u���@�?/&k�R�·�`��	`p���~E������y(Hԑ��o�Լ!ObʧDąݔ�0�ɰ�R��c_�jx��^31��I���);x�[z>����py# x
��]�lպw(3+VP���������7t�7��- ��|E��sn��-D�W<���PI���#���!�+]~,K�����ӗ4��Zz~���7\�h���1
T�\�|Ʊ8w�(a�@O7@���v^�P�A_ɢ�nŌ���3�W+��w����A�r+W��L @�ߨ�1������� �u=F��d�3�z%�Ve@�GU�
`]��<Q�&=�氲#� ����&s܉�	MĠ7h�W�*�it���m9E&�6�2���V7�)�Ų�F����0�hC4� �#-Ѹ����Y�X��#��يp�\�$���,��+pvh�`�XN���p��k��#��7�~u��8��ϝ�,�dH7���m�l㷶f���
X4������huL���H�{�&�#v]��!5��&�������{AU,{ N}�Ӥ���"`{��W�1(���Qc/�U�0u����1��~�����p�í��Fo��k�ե�@e��C����d�N�86�����8��p��N_*V1��/��///��%��lLkeX�l���m�U�f��7C�
2�5����u�Y���j��F[8L�)��寄^^cA�u���k/�V��Q"���;E\��w��ߎ{O~�?�M
���h�|�H^�cY +ݝC1�a�B�5�O�c��h��(����L4�b�V�!5٧�Ed�|9;Z'���jv��4��r���ck\wȤM��$���Ŗf�lē����er��_� ��^�'�M��K��):�t�����SО�Uvr� Ͼ�h�rZ��y�A�����W,2y/��QE{`Bٞe�x�[�T����.�l(~�p�bz3�T��am\�b�<���/�Ex۟Ŕ���1�p��ߠ;�M�4�j
7�dF�Vȑ2���AF|>s������x��gy�pͥ��^W*�t�1{䟲#�5;yvl54i$�ȹ����pqŷ���ھN�M�'}����ղC�v] ����Gt!�ѱ@�tN���.���M��!�z<(����c�SnRq/ެ�U�(hg�B溉(E'�-�5vs�oa���}~hBH�`Y���?�W����^��,�:�A��ߔo��D�/��Ƒ&�w��SE�
E��X�F��A��;/5�c.�E|�,�u�VD�v�|b|���X��vdj|�p	�C�=�͉�p\��l��w���zr
y��Q:<�N����[<�(���l��^�ܚ_�/=w�h�m��~�X�o��D����c9Z��G��/�[�~�߿~��h�mݹQ�s��u��Q&#��ZE���:4o�]����B��%pw;{]/�PgԼ|��1I;:5�l�sw����8���z����z���k%�c(���`��
��~Ѱ��hУ�o����(^&K�,j+�����Sc��D~j8���׾��Kus�O��#C��=e����av���B��} �Z�1t�l������7�jʃ��7�A8�w/���\~��T�'���IK��?z<��W��#���O��s��2�?�]-��:� T��5s�����Tuj�����y��7�b�K������N�n�tiW�H�كS�D�S=n�{���V���eW���[��oAA��;���:����~-A�j��4Qw��R�
�97"[�~��*���'iO��8N��w��K�%m�ED1�m q�xL��xI���)w���W�/ં<������5��=���-���d���%N�TU�%�% N�o���aQf���k4��6���oI�3�u���`L`���(���VU8p�Ɯh!��s��	�pe�iߌ#�Q��M�*��5T�c�f�E[���%������PA��T�M�%$��7��[����A����{�2$�zY�i�d+749��Gd^�޲�ʑ8_k`D�8m�v�<寄�'�z�<6+��|}-�hCEF^�%j ����k������M?Sԥz`R�c�|��X.v��}�����Xn��[����a� �pb�QZ�'aR��h[�7oW�������Dzp���g�8a�GJ��[����>�,���&�����9U��Qk�&1*s�x4�y�@(�-�nŵ�y�\|{�x#��I� '����˘+ܳ�vS
D)���9��M �m�6i�Yec���Ԝ�hz-2R�-y�jF㯭�`�%诫��:^�Ң�`�ne�L�-�������<Q��m��<{����|W���nnAɡ��-K$.hْ,�k^0�k*��B��d8��z�OR����*�e8juj'�dQ��Ο�� �ڟ��l��h�Pz�6`Dv��H�ųb�p��3G�_o�a�ïU��޽p}E}�[��L���{�0�.&�`�O��Gv��i�>8_BR�B���2{�YK=�H��ErL��T�(gN	X ._w�t^�H���*�:P(Ƚ�?��,��J�$NMCL�3UH�%���B���n,E���U%��>�� �IƊ:�s2��"�����}�֗uV+n΀��2��~�;<9r�'�y�3o�� ���K$�f�O/�ϳD�.SF	��Xn�x��&��	���3�N_ۖ�����۪ ���:��~�0cI"|�`H�g��;[`P&�p���>h�N�]�����G{b����Eɥ��j»���cJ�\5��..�g����,;E����M󾭣��.ZR��r�1ZE��� ���I��^(�c����
Φ�$��c-�p̖����⃂�ތ�wO)��ݖ���ZV:�9�kܔ�2[���
zB�y|5���4QR"��.˙�D�8�O3ZY�)��m�_�D,�w��n��ڰyF�6(�رW���+;*ɕ�dL�A��!��R���A�O�@�_�����b9��k��*���Y�_yز�#x2���d���|B�:���� ]ްN��㷲�z�_΋������i��ֺ�q��:}Ck�����ؑq{��D��(I����Z���K�,q�No�s��VQ� N��D�|��y�9����|������&���;�T�e�S'��������8N_]��mcͪք}����Tb���'�4��rC�m,WIE�B)�:>$����P��^��8$H�xõ�w��V�Zn�.^4�
���_����d�G
(�k��, c��(��-��ܬ� �/�Q��mj����/�l��NS��1F��Im�����YrdX�7T���[-���������@��^z�ΫC��P���ݩ��o3>�b�axX�&Ȟ����>şD��Ay�ԋ\y�����ģmT;��/3V��ݳT%�[�M�|�O����k�:
���M,JH�NKƽ�,P�ĭ�Q��{�4߅��]��.Q=ov��--��7�@���\�E�i([���ή�`��~,N�!����q\��=ܙ�{Y/M�����xU+�B����� s�c����ΤJ��\��o��zxǖ�5zlm��1{�ɶ��fՒ�_DX읾W��h��8禈�i`A�+�> it��>$��W ϫ��K�9�i����cˊй�d�W�&��M� +�n�m%������X���v���W���`a�!T)���&w��,��Yy��&Rp.��W��c|�q�����%��x�'ތ�L�ٞ�/#�"s��܇�"(D��~#�<p�/�`P��2$��s+[14�%�J�ii��~�Y��3�$�?+��V�d��ǂ�n��F5y⮌��\u��w,.���z۰9�jqBG+��岫�1�ݬ=�)z&�V/�V�C���� D0WO�4�耉s�?�n�-�u���*��-�O�&{,�?�
����z�)�ڲ��y�g��to��0Y=�7���i�X>�rR~�Ծ7+��7�TN=u���s֬����c@S��cY�a�[2�↢�#'�����׽��
'^�j��U,]X�G!SE���NѰ�h�x߰*�4:�6�t0����:��FH�mK2�m(�"��O,�? �S���	�>��0A!���ЦM�Ds@���Q2�����ω��] �� �~���R'�!}�*$(���WN�\<���Ұ���p(u����O1}�	�WO�{@m,kqY��}c2��zfU3��~�����5[:zYE�( 
��m�9ճ����qJ�	���Qf�{ ���[q�� <g@؞��e����W�t1��ց~?r�^Y�~&B�!���b6�q��_AS\,���Bo�O�i����'�3ܨ�
�Y��׹,���ODg�-�^U7��>C�u���~X�Eb9��S��Y����0��i�N� �V̡�7I�5޷��;�M64f���:��d97��s�W��o� ���/b<�`?���o�f�{rc�}�Ќ,[~�.0�32�<�Re��k�1��!9����.R0� ���_�R�C�Ԅt*��>�t�e ��Yq%�=�M��\}l��H1��0�ȣ�*;�ZrC�n�뗹g:��6���ֻ��k��ic�p/&vA�@�=�RtN2��@a�Nt�,{�� �ުmr�-��Y�<���Kc�	�g�E��L�B�w��P��80��'�t�|S�%*��w$ �g�g����P�O(VF��+#��rD�H4F�ge���x"`!��ΎD�6���T�fe9��Q��6�lQX�cq'�{������gFE.��<ok��=��3y�#Gո�X1�<�]C	_�Ig���'�ns��z���ʉ_�(�lи1F���5��uh6
e��Of{�����-�,��q�~�(-���+��:����bl�{q���>
Z����_q���f�=�:I�Kn����1��O9�{�B���l���9|Z�/�3%�s���8��x��s�-J]f��²��:���'.`Ae1�Tyh 쭭���2ɯ�!.����_"���	����'xU��	K�F�"�cw7��αl����Ù)�a�q�r���/Do�z�1E�WX����P!�
�#q=h���G�,tQx_W�!jS .�A��A���u�?�8I�7��t<�Sx��_RS����'t:��{k�ƨ>��a7�%9O�ɥ���-WW ��.F��E=��(Ė@���{_m^�sx�d��J�����l�J$G��O�-����a)#r���� �߽��,���(��)�:����66fp� �VQ-�q��xy^�K����\�Lz���s� O�/"�Ɔ�H�<E�!8���#��ky.�p]@�Q �]S�FX<�id��Q�D���fζ�=�U��1yI�B�gf�N���}�mȟ��Q�@5�s�:(-�4uT�ѨK�w��B�����A�(�ܨ҄���%dF�	�g���ɨ:�bhꨊл���ůuG�sT����f ����_�/����|�tm˿�u{J����l8���ǙxA_,
}�pl�b$˒��ݥ�a�	,r�Sq�I���'�ȭ-��� H��3}��eUe��X U�X<:ÒB6{d�C_�� ���[��8�t)���:~��f�W�y���r31Ɯz2�i��:'F=�咦ACk2�m�z7`�=d��W�C��Ԟ˵�����B�BQ�Ik��$C?. $��T�)8���mڇT?�j�*!ݝ�"�QLB`p�]���N�O�n�O_ӎտ��c�3���y�G-'i4�ÑV���+�}[go� $	�b��g��>o��ʘ��Vşk̬���=f�r@��$[�ުvKX���*���J;�Z7?�JvEb���.�:�����k��|\�w7d�ܵ��	��3p��w�h��ef�i�uؚ�6��c"
,�R����:k5!	��Q���i�z _�]�d��*Oa�G2T�`k�-X�Z�x�FK_�$u6��x�=/�P+!J���'��1���!�i�����\j��S� �\���n1NX�W��˛���WU �Z�Q|8���sw�+�	w\���2̅������B3�͗�h��@�aO��'���Rt��QO�R����L�����U��`ʒ���RRr�_�oB��f-���<�s����T���Y�]�K[��.�d�������[�ًB�r,r���Ca7�oFk�����S���]߿�l���mš]�=FM��6`I��������9 �?I/-2�X��DU�u['Ibv-���Eo%a�D6�L��� ;�jDY�����,I�x({|YO_޴I\e����,�h
�!CTS�	�v���Usy���:�X��n�� ���4{��)�j!�.�b�Sy19v^��������5+ׇ� �ǔ�4��^YL��.����0����L�u@0j]��]�>�~ֱ�P��f�Ӊu����Ӎ�� O�b�� [r]]*�v�bJ{}��#\I3�՗�G_�z�p����|��n��V��:,F����x�ޑ��(qz�y%4��H2?���N�����4D��#�y�0����e O�^�XX=L����NO\�).?�����T�8�§��1�H�qq`yn��'@�b�6�Nv�e:��F7��@�b�M��T.�$H�{��V	��t�+�5�Z�F�Ҷ�|���|x�E{D<0-����<��pqj"w/@胋����^���z��u<�k��W�AK<_l��,�ꥒ�o�Ī/���'rh�Խ��?�����
��9��M
�n7��.A��buD}��T�;%T� �9�����/�s[IH3{��r Ș�@��1N����e'lr��m<e_��`a�G��|&$���������L��Q���Ʋ�д���n?���Ī���t4e�BC3�$�iu/P���c�-��`�bށc�1c)���#T�^�n���)�E�a���4Y]}�9D�(A�x�,4�3�����Ny«i�X\h���	�>ofC�H�ۙ���6���1�UAU���,!ZX�4�#I���"3�8�i�y1@�q��M��J�_����d㒑$a=�%s�[���{M�uCdqK��"2��3�j��.�I3WnO��mmՌB���:�	��n����	�H�Hةd�O�o�Htlmi�N6#���Zp��:O�����}��y6
���d�^�ZJ���Δ��ٙ� �ׅ^	��:1�g�q�wʞ�Ҥ���o����lͺ�ND�ǫS}�;���XK�!�0$���n&���5��1�8Ж�����,f�d[�؇7S��F��*�A�qP��:�/)=Sn��O�v��9�`�ܑ�(�?I�l�<"���fD��Nh���0���y�u�9B�C��S�=`0HR��Z@�Ǳ�WEjp� �	{�@��N�G�(1ĳY;�(+�����D�@g� �WK��(8Ok�� ��A~>��V���]��U�E��<䗰��:�C������,L�Ivj^D�L>����*���g�v�
|6�-�q9���:�cvX2�*o��"����fy�/���7`@�HFx��
�?�9�����g���~^3ga�~Ź>{� �Y <y��.��Oآ�o�t4:xuZ�}�4/�'/o���)�kC��=8
�4�����u�_��� �PrO�Rd�F4��t�;Ɨb��K��Qi#R��X�-��q�P�-�D5�j��~��&�Hb��1-,A� bdf������[h�E��.�ic�[���b��M�j�@7S��R6��X)M�Xp4�0�BH:w�W�[��'��s��6�L��!%��Wwͅ% ��X]�pۼ��؉j�Y��'�A9j�گ4N=&o�	ُԗV#�!��|���sHcS�sD7F-�R/�S@�C���!ۿta]�����9��7�CN@�vܣP-��Q/�2٥������X�!������v ���W^aU���1/0~C�� �_��OcY�%�q��D�"��16US-�%�]��W���)�ܐ���>�DM8'�XqĠ��X�uj�����2�t	�37�4�^�t?�tTEr�/�qu˒�Ǻ��B�!`s��&�������2���	?��������@X+���D�(�E�R��X�qlk����m�%��MB�d���잼�w+���YN�t�x�et�&P�Ԓޥ�>����H�wԗ�Ɩ0yfD�q l�����6#^a�e%��a�����mm�{�c�R���=���@��`Qב���!\/�M��ZIk�әaշ	����q���M�;,��e8u�+��8P��`����-WSg+�����.�����㽶����L/l�gCx���{������ao�]�O�y� �K9ɿ?5E]�5�m3��i�y|�4 bR�c��t~�L�Z,�8B�	K��e3Qe��������k�v ���]��hF=p@�d>�9�Ƶ;D�-60�R�
�+UM���RgŽ<މ� _YZ 8Ά�i�\'dwl�xA|Is��l',����s�g��yO��QˤX��4�*o���ۚJ��� [��=���c�9�C���=�/���qy�i���Lq�R%/��f�x�X}���|���s�{��x�l�2�[)yEs�ݟ�`�Y|7��;�VY������O�����-Ӄ$�H2k�����Q5�?�$!+<��h1���� d7���ف��2�V�fsi���p�nV).p&��솠�/�����~ M�#�wm��y�_�;�ZX$kwe愔xAmQ��K�-��8l4�rdĮ����gѢ��ag���<�z���CV�ﱰ�K1�+Vj*F�]�t���	��6��0R�E��Q+W-���LzӤYqn�`�wޔ�4�9�!�ڏ���C���U|dK����>rjs,=��in�!��c�a̸��z�Ȣj��"��ps*4����s=sP�W��wkg��6��sF�(�b䵐&^�&�m�xD� 	m����:Rs3ԯ�r?�o��4^7�I�������lmq�"Y,���r3�*��B詠So7����tf���+0Ä���)q�8ه��Q�nд��q��'�L�wЖ�F�d�=��p4'��7/���g,D�'�foA�L����M���r������PG0� slt;#��
ǩ��q\(ĉzoU�g��'9�|�xTk<�F"�k��{��oY������	����ӀY^�6����-��I�h4�Aa��/�Z��Uf��Dd�L���=���O�_U��݀���{->ܐ�����U9��#\W�fd�ri���-���SO�`������!���1��O��� ���'�����&U%��n-�v��AFX8���u�bX9hk"�%�� ��7��)�}�E �e��؍���F��y�>Lm�ֱ*��͡�5+�Dq7�?k�A���K��"m�ԩ;._%%��	�ha���b����o��9#z�aP�4jkR�#/�� <�
x�!\�M�Zãmp��Y��t�4׼z)w�J�~-���p�-�ˁ$c�I�5؏��E�h�2b�!�X��u��=����Q�uuI�P:�
�1.}7�1���<È�/Uɦ���V�� K�;
_%2I�Y�@�tЪ�<��s� ]^Uc�	C0]K�'�%�q��8Kު�n�E�g��pN���	u��fl�gE���G�/�,YD�@#gNn�a�\��T`�{��ZN[֩��wΩjc��,��� �����;��Ore��|��]�D��;m)�����t��q����K�~G��]D��� ��3'�����r�玎��������lP�}�(�e�QXY��F�k۫#�rЦ�t1l�K�CJ���Ȑ��P��/�M�z�!<z}l�_M��+�Ӗi�A�x���1�E{�x����Q��dOF��W{Т����kFex�	u����Z�3]<�X}Z:�� >����Z��p�<��;L&Cu-d�����,<��rk�t4���J�g�=�2}�B���I��Tw�}$;���<�H��ws��`��|�G�y&#����U�U��f-haǝu���5H�;�|vV�A�Q���_]wbhd�L�:Z<��:	`
-���g0�Ms�ZS�7��`�%y��)�HM���mn�J��iM��V�����0�qi��ONTˊ��Z����d-�oΘ�\+H�e�U�)�&ğ|-J�ΐĦ��C{sW^�^��2b�w��r�
{r�w�o'��ˏuI\m���������1Y��R������� 7��H�7e��a�/Ӎ'�lw�H;Gl�H�1����	/���]k	%�UwtMҹ�0��P�o a�D��M?�+�Cl`@յy׵]6iX�D䥍��{�� �4���	N|�H\ۘV(��e�q�UF�"�x������Kp���MG�����q�)�x���Dơ�W.Á�rQFK�W��d;���e� p�Po�U�;?,jqY�I׷ș�=���������-�K�<\������o�1зLu8 |����#4ԛ�ù�`<i�h��>e9��8��܍V�:.>g�����A�-�l3/�W�:�WA���Z:�J��+�Qs���Ԉ.�j�g,�c�-�y1$��U����KGZ��nm�)t��%�yu�ZuEẺmr|3Gm��]��ڟ����.>�\�b#GJ����a �y0��ʄz
�_�Me�����/�>�9_M�]��}�r.L�����:6�Kn�zO�v2��
q����O��cbL�fP�+�9|_6�ӿSV-6܌Cs��W�c�V&!�44�K�B���[��I2�t�?uc�DĪ_� m_�݅�7D6��(���i!�G�+�d��^�ӑ��(.e.v�,�)hu�ё����J�����R��]�V(�wU���$�$��M,���Z��7�N���jBс͎�� o�#�!�"�{Z���>�e�E��XS�..1,�t�Y����^��f�u�_]�r�U��zb�4��T�a�7ٟ�\U�L�b�5J�"�o���C���u���X�\cg��eS=�i	g]a1�	)ofT���(�ۀ���̠^���:�Ⱥ�w��/Ui�6a�fO~L+ ��$T�T�&W�5k�ufUB�9i�G_nB�E'�0F9'ʰn�m4��"&���$�9��� H��S�U�$��#i��,������S�P�׹)IE3jb�U�?�".Y1����--����.9� �$}���I��V�>��7bSqf��kL��L;Z�Q�^H�!o�5���H������ghG)S��U�3�J�gQ�-_Jڳ�RK���4��6���	g{���c�&�p��;x/���D-�.\�'V�g�#wEmA�&��#�����R̃��?�I7�z%�����@}��^��
�ޓR4�|����/,���������ŀ�b�#�VM�x@�/D�y��f��L4���o-�;M�{N[x�\ZQ�?���AY=�G/j�LLoЫ�#�!�f�ǲ"{h(�k.*��av.�{&p�Y�h]3Uz�ЕHڿ`�j���w6 ���Db���(�w��Gσm,��������W�����4�w���WW��?���x�Ga^��9�{�s��ы�fxUm�D�/�9P�P�A��zgy����bʓ��u�\PP)7��Q$��}͘�;�j1��fP�����)���e��I�|z�z�a�Z�Ш��-��)!"x��`!`�(3���x��yZ����G�m6 'q/�v�j��J.|�"a�_��~��!�"`�G�[60�&�F��#������f$��:1��9���;{�#�jO��+I2'})��EHz��e:�T.���@��x�s�"V!C��������B~����Ͻ���H9�YZ;ܗ�N�!9���.��(¸^=��*�z�̾�=��'NDE3qq#n�	��B�C^��Llc��)�ױ=�����S9��6ܞ�W�]"�y��*ח�?a�Q�^F�L�~�]a��+f�]p՗�����7J��e�#�+2�2�����B�#
55�+��u �h�\�,���70��:��|y�&�x4>�����ĭr�؏qh��3��G�Ȳ� ȯ~v����N�9c��� �����kb5e�5>�i�`�Ot���<Ĕ�H�YO�wE0�D��f�w�������1^��pM�W�C�,P�ħH�)�j�d�K�x����̑�t��� -��o�%�a�5j�Uo�c;w8׽b�,�y�%��8���>��u9�=��NO�H�@�R_�=��,d�	�����3�!�/ �1�LB�-b���ٍ�޼����b��\>wv�[&��̏ΛjC��4~�τ�4Q�;%ԅ�vοLD@�T>Y��U� �0�:~�÷�D��`�䋩K�]~�#e'���BDp�^�0��
�%���8�Wb|:��ѐ��^�*�|���a��Q9s�{��1�!��b�� �>}�=�QN0�]'l7�*k8l��s-槊�+�����R�s��5E�#ų|��FN�,�G�*5ĦyY��ǰ*B�6����_FXR��Y���&^Y>��W-�ݧ<�A�Lkͭ�I?H�`c�^�儌�hF,Mf����=|(�r��0�*���kA���b`��Bx�?s���$�gmi���S�ȹ�����eCtG�2jw�ڀ�n��ڜ�Oa��ݸ^v"��z,"s�"	HT�3�똯A������Ep������ԝ��03 �bK���p�k�Z���Ҹ��񢖺�VM�;� 0�ekQ x���D?��B�誎�+R�%������EڑI��ws��b�����5�����a�)Z�-�E��P$�}��������@A|�n�+����#���P(��O:�Յ�'�VBr�ԁ�1�#o�cBt>+Eҧn&)կ�Γ��+1���O�莭�͐�\N���%��d�^�����>�n�
�`���*n�;��H�.}(�6��;m��
Y����k;���#I`cY��8{�`a��,� y~�"Ӓb�,8�	7p�1#,���׏�i��F��8o���7��m�@i���+�2���|�
���P�xm������Y�������q"
�i+J���}ȁr_!�1ݴT�N��Ɖ�p;#[$��u�b7U?ISR�t�f�,�>2�ʂ���Ь;eq���a����qn��s�U[�g'9?�o9es��+��_EEo���,2����@ʹ�L=�W�>��7�rBĸ%O=Ab�+�xI�p�,o�T�y3y%p@��w[�%��_2�,�R;];`Γn��m_�q��fd7���
X+ǡ�������^m[�W����.�\;��C���W6'�T�� �M�a4=M�;]	���*����xZ5�PvAR���P
Й�O���n��q��f�☛���9Y�CI��+j{Pb!QP����?��O*;�x����( O=?®�7����x`��2I�Y(ҥޏ~$_j7��wh��HK�]�QDYd����ga]N�f�	-e:a�k�$�y�;�g�&���
+�SE{���j7�2�� 3�ҁlʂ��Yú��4p��$_I5��������j�������W~�2��E��t��m�C����o�]�=�tj�c�ĆnV�G>�t�Y�~���j�l�VC	��OWz�l�B�`�v�89�<�@��"�.{ Fՠ+4FrJ�Q
]f	Y���
��M~w�h���և�8�J�~���~5Ēؚ6��ԖQ�x�B�1���XZNf~��(}JFW"�[Ѱ�g.���<6X5O��҅��������zk"�Q�7@� ���}J��W/�ؕ�V���{挚��ʄ���!Q�z��δ�*8S����
��!�^��![h�B	�Z�ؤ�:�
���L�S�|ggV�1<Fc5�󴽱��� H�jl-����(0>Z�Z,��aO�����[\�+&X
��.���Y�Q;��Qb����.-�m�6�!V� &y���[�Aio͸N5.t�KK�An��~�����Z��9�_�<"m:���ӵ���� �~c�m�2z�E���!�'�,t�#�xz��)��A'5o�J1����3>��_!õ�w:���þ4�;�ϊ�"l$y�J�Z�5�j�AāJ8{����eI��pCƆ �i�0��݃1cݧy���0MU/�ǣ	tr�����^&%���b}fO�yLf��h������CH	/�����%
�O�	��x[]�U�,����}>h�*�V�>E���UB1׎������e�"�s����SVaWԮZ��n��#�КF\X�%%LZn����
�(���H�|T(����ɥK9J)g��t���?��&_h��~�����Z$3��������V
a��Zvi
;�ń�/�+��,�}rqb�=Arm ~/\��YП�D]��B��ӕ�Gw���Oq��iU%ٰQ� .a9�\���ڙԡ��T��P;��|��ֵ)@�|��2gi���P�;x[��䮨t������|zD�3r��m�-X��6<;� ������pG�b��_ǁ	Fp��jY�{�h��NXG}�~Qbл$�j�52dȊ����_0�?�{D�D����NSC
����Ҹ:����b$�G�2����t�XB,�riqZӓ"��l�^��$�sx_��q�1v������
����^ 44�V7]��<g����F����wDC�?�ÕI�<k8���U4H6ȼV� �9�e,���'E�Z�'PFe��a7%}0��%�|2�8�t$��fFx%�5�`�?����_��f�m�
�&I~�.c��cy�M���	=�ȥ�]:_F݊y��,�-G����o���	]KR���0����𫹹<|Q�Nq�,��LxO*�����#a�g�[�*�����U���yH�r���H8ge��`Ԓ�F.�_�����Ru��vpZ9����h�:��,�/�mf{���lIy ��WVGc�xH�ؚus��$ڗ���\!��־u����P�g3C�=̖^�f��2JU6���3�B�0O�3"Q$.��p�f�1��7�8b w6�8wOuBv� �RE�e��Y�s^�"gđ�KP�?F�\��3.>'(�=�a�A�5��T��Li��e��&��-lq2��pefHHF*��W�Z�-��F�6�׎
�~�!=>��a`h�1V�~)�/
�w�SƺkQ�=/3K�׵����V�+������Rp5�̃����P�Ai[n3j�l��`���PP�f��e�����E飇��$�#v���@+���o�R�mQ�@����i6+�T_(�>���Q�F�sl �T0e-�;�G���N�٥Мǚ��ܿwt¼�4���8�u�P,vq��?p���<���d��9��Y�:_��8+�R~��3����-0�x��w�|@��$2A��O��l��O"��q�xa�$c�qOo_�ID�����z�T�_��ʧ��Q�c��U�I`ל�B�7Y�Qc3Ɋf��a�ج���2sF��2��Co����Z\���r�ޥ;j�6xP�q$A83������Pĺ�:��X��U�DS�Z[�)��g֔��g�T��� 4A`������`�#�����=�[�O�-�P{�	��]�DI��-5��P������ �Ed�w߷�.�S*U��s�N2�[�R+�;�j�U�n09�u��,ݟ��C���|�E�9F��A�@�#֏��6u�;�1�y���6���AV�.�����>����|�/�Z:��K	�`�T�~��)IVGK��%9!k,m���<���Q��u����4GN;S���'��� ���B���і�e�!#H���k��5��YE�doWɖ��Kr�EZ|�( H�٥�[ɦM����B��o�e�G���Cr]#�3��NF��tV���G����&��o��B�k�,�Y�cZ4<'pT4^�*q֑/�6����mĘ��#:H�m7��z�iw�InU,���&פ)�6�H��;����Y�n
O`�A�+wk7ý���?=�j��k����O5��Oc*0h��B�e���t�ۺ��u��p˲����6P��8��� ��L���g^�; ���`"y�w���`XLQǧq��r���n���&L�*�?�Ss�,��^|G����n��>��/�
��S�OJ0ή�	z�m���MG�.���pA@_6W/u��D�D�^�J�/���&�ÿ�vݭ��!#��qz�u�> �憒�{�C��gJ��/���_*.#��z�p��>��'��#-x�:M��sؒah�&4z�n�p��� �����ej����8&=�I�
�c�/S���ϼ"��v�(j�Q��a䫜F�Yϒ1�"�U��-Q�Z6?���|�@�+v�Q�PC���B:%A\/TҰȺ�|T�H���E��h_d_�K��2f��*�cp�̃�ُ�[�W�@��[���&�"���A�2�K���f�׼�*�2�����d8��K=�0���9�:�<N�R��;�`!s�Ĉ����]0�׌-òƁ�+}�zm!Nt�d�>V֘\H�s�=�	YX~���j� �t�~p!�[��h|{4�XX}�����	��AC0���c���D*e���h>:�RKI6�bi�/��Ű�T��h��KEK���$�țR��?�U~G���M�Z�ϐ�#G��5Z�c;�[Q�!��d�����T�U^R��O3#�z�WV}Ni�d��.����1�v�tr[�=��W�zhT"������=:R�V����e����ᙞ��)�:�#���%/�Z��(����Bc*�: G�ߘ��Ys�}8Y=����Ɋ�����s���_w�o� �>ڣ�]!�r��'�)���Q�j@��D��Ş�r��m'�v����b<�H�p�y��N:�
�n�0��@��L�j���O<frx����-m%)ᮩV�<L�G���ٹb�?�fo�rf*��?����W#��怊���*���V����"��:��ο�M~�����Y1���M$[L"���R�)�ɥYω��R�+�+�d�M�{V[[��&��Y����5����v���r�>9�QM�Ӻ���bxA]_y��)��vs�շ�Rb[OW��T�Ӫ{hz������ �]{����$�p�6u�����7}~&McW#��#��jR4d,�yt�)&����.��
��P����x�L��&��Y�U-�C1���I���QQ��N̠r\�[���n��ڔ���o���F�޾���5�ݧ���OL�O!7�z���q��ߗ�L,�8B-���l�[%�v[7/÷(��lf��~� ?B0xӜa3����j��� �{�,��F�|�;�*��J�X�Nq��#�!�))�ӫ���D�pK�X�h��	`��3e,�Z��#"]>u�ܜnP�����y:0�M����4hӧd�2�AQ"⎉�my�\�Z	�+1o�ҝL��Mx^�Z�ht�۴5��cF�fVX�R-�"a�wHwh���B�e�0D2�1��?��ki�b�F���8R�浽e�;��;D��)h9#� ?ѐ�|�S�wne�àn�c��ʳ��1���v�^�YJO��9�x��8z�A����1��lpv.�kCD##c/K����2�>q�6O��.��Yp@��.��jj��bU�׃��eF	>��V4���w�����<�Z��5҅�J�����J'��${j}/!�b<B���x"h�$ {"h��][����i�T��ҫS��F/�ӓ��4¤L<�2U���Ƨ�%���Y��~V��o�ȱ��S�x/9��j͎�BJ��钼,'bu�O��/��9��~���PC%u��@�^�/
*�\�Q�{� ��z�F����R��Y�֔�w񫴞����@�wn�����sbd�|�r��I�@!�Ī��B H����/�m!�j���i���m��#R@�(��.s�+���g��4-���s�ϥ*'��Ū�NE'���lX���a��UaB��s�>��Z��`8��%��]I���!��C�����ܫ#}�����\h�YV/@Gԛʪ"q��z� r�s!���2���U�P1x����"Տ�m���r����/<
��$�tܨ���3�c���u�����v����~l|�#j1������GW�����x��^c.[��|<2FsF�3J弣w�� �k��ߕ�&0�>��h��"����0�x��cpb'���Uo�B��K��J�+�Md]m�F��s�Tܒ��c�vxTK��@E�*��+�[�/��T���s���4_�w��R��}���Y8κ�������%e�O�"���'o�d蟞��JF^�K~���q���]�6���8C��� ��r ��Q��,��
"~p��D#�1_��B��(��Φ�������y�&�4����9���J.~�pH糛vo��t��Gqi�O�=v�	{�Vg*-WI�|�H��%$ϟE�G$n?�?/u�t�4�?��:�ٴ�n������%�a|0�#(��������<�+�Ƈ�v�h�Z
0c��Z���]����c�Ʈ�|Z��6���A�Fr��E��PL�ܬ_����W�N zL���^�m�+!t�@a*�tB�.�2C�v���E�fX��>/J�b���Q�#��ne��u�#��AD���+U�Q��<�>L��F��#�q�D��q�p#EXy�|�պ>�����BM�����P�� @�~��#�2���%!�8�P�����n�?A0&�v��\�T�[���SٺW�y0%8f��i��"\��
\3�I882�7h��{<� z=<��+~��(���(�|��l�Tb�O�9F@���(:���!ƿ3W�ϋ������A��8iX<^���H��[9j�<Y�Mԉ���)�'��i���V�,
���Q����Ó�LT��5��]�z�P����e�|η��0�Ӳ��f����j�v�n��&��ؗ0[��ڄ#aO$�U�]�tYk��\$���<
]8}�?K��)�*#�'�/ٻ�/c���|�?�H�o�L�k6	"�ݷd�Zҁ��~��a2}��q���1Ю6���9#��H������w�ɏ΁W4�x��M���%*`%�FBud'�����WJ2���c'��.R���1���K2d��5H0IF�u~�	�6>�@�<d�z�T["0�v�R�]\������gW�w*�T�v��b����V�M�
FmJ��AuV�9ݒs%jV�����A4�\��8q��ܫ	:r_�7��B��5���WQ�?�)��f;IN���4�5d ^n�`=�]�����5B�!����d�hCd��5������@�,O5a"��](4;z��aR7R^����t#H�pz�������,����ds1��:�����9a&[Դ�t{�I�����?�*������tB�1߾�W�R�?q��li�����;<DIͅ����,����𞼉*Sݺ;	�B[I���i�c���g)n���k�q�1 �Qf��������b���ٶ��{|w{[�n��!��=��8�F��4��_�_�G� ��T>ٮ���f��b�@�UC�Uko�|��S�F�b��:�7>�Y�Eac�Zv�-�z�o�ر���#���Gi,���9��aK:�;�W�Y�(��� 8����B�ul�|ޕk���4����8����s;s�њw@ �
�b�\P)��m⒂"�1^[>K��/o���0���k�q)����(�#n&���1���[VK���?i�`[�哠e<u=������j8y%�SO�g}u%ro�{|���R��CK�{r���~B�m��ֿ��$��z�|���3��vޥgSn'_�����X`�%�]�r��yo=2�(��)�*�u�� �S:���,�4���y��C�����0�E�_��� >��6�kh�"���8�	ٯŧ�M��l̈� &��l �	�殃��.Xyg�@$l�N�/ֿ,��<�?zF�n~e48��%ua�3;��bt��n��R���(��al_���.*��o8��\{�@�?�;� �8(��Py �eh�c�+>��o#Sш~�'�u�������z�=�����3ZI�E���Y��V&�J��~8�nE�V�Ėҳp���E.n���uu�~�X��v���>f�6z9P��R�̔�=��L� ��*��`�5�*���a�o vMD=T.�1O�V��:�G�#�Ť�<)��)�_�\	�Y��^�� �:��m:]ƍ���<%I��k���o���ƨJ9��,��ތͬG�b�yB� <�E������H��&�&}��(W١�'�){-���m�eH0\�o~��L��]9}�p��P��'G���">J�-���Q��tw�D�#:�vׯj��!�;Q�Q���-��Gٺn	�k�r�&]�xO�,�lw���́�>��i��b�Xz-5`:��y��T�f�S�C)>w*��u�Ն\�w%s��:�?
��/��6�#uԪ8�_��|D4SA��7�Du@:�/�@Ϙ�2m'�5�A���p��x%�AP��h�N�C���i�����=\u�q"�B��2r��K�wd|$��H��{����T�P3�1����u(���|�K������q�6F�������bچ#�܍�M�_�=P��R�~M��%&,QYWc9�PԸ�ت��O�`S�_*�R��&�q��̩�ު��8��HM�"&��,�9~��J���3��Q%���5H�<	K�햿~�q��u�Z�-`��fT������R�+��G1"���x@	��*�MW��N�w��������������w��>����A�v�}���Ȧ	������h���5�ĸ^9,����P�}u�&}����V|y�)�Q�f���+Z3F��Ճ0HјN��Q�ٳ�=��l;ır℥l#�H��� ���Gb,��l!������Y����s����um/�y�(H`���$D\�+���;$�$�J�#&��f�����Z�f\JA��|�%��gn�Z�����a.�>�iM�SҡZWй���*S{᫭]yFG�V:�+vvt����ː6�	�I�$o��f �f&��[G�z�A>&�'�V�����#�3�)1B��h�5����e�e
�gۗ-K�j�Yc��%M2���f,J��� �)�3i���/��_�����
�gހ�㨔�6/�b��sb��wV;/�,ZAg�X;�4��$�R��~%���jG�@�
m�f6�t	��G�J���i��f�]�N��#��SF�H�� ca�]M�f��t�w :������R(Dp�㕞7�L%�����g�(��|�\�K�U���E�j����gB
��W�1x|���ʛ���|����&-ʎ~�i	;ZB��BQDt;���ihvn��U�ԥ6��§jna�"�S]�z��MM��<�v���U򑎫H��y�$�+� ^~E,�����dF��F�����;xʮMM�,�)�)=�U�����2����$A>y������0FM�f�LcV�h�?���	��vz��ɑ7��?�L߲�WΨ.vgrF=
�����VV�(���دf*����`�]=_��
-���kk$����Ɗɼ�*��q��k#�鱿NěPd�)���b��(C�9�%(ה����6M�������ѷ����e��1�R��%���®!��<�;��%�7M��='^���h3��XW��ž�OD��ak@���SV�铮(d�f�`���ٞ�L�;��|��#�!�.��!d��M�=_�{���ƋJOB ���W�0S;�C��N�y��	�A&��5�s��R�;x�>,�=����%(���(��i0��҈�țyjhe=��$�Y���.c!����M5�l����%>3m�e��<+{�l�M_W}G1�
�}�(��J����h���W9š�l��~Х}*�[�H]4�'���&.|I�%�&զn`z�:V�v�2&u+\p�(n��ᮍ���K�s�I-��J*�SC1�b�C�I�&���B2�����<$�ikq���$����s������Nn�x;��ČD#I�l���U4�ip]R�����'朌�@���8�j/Q��D��h�ឍoM�	%oO5B%�@�q��o*��Yy6+�t��v+�4�)	 � -�!J��߂h�B����ѻp�4�,�rL�����e�����}�m}"�Q��)��Pt��eiX$5������k�zN׺�5��N�?
�"RV1x ����D�Йw?z��D��>�:��(_�=�8�m�3�D�S��FZ�Z�z������	ۗ߂�Q��t>��c�9��a$;mn��j��r}�>���B�J�Ζ3b��3�>eS>*ں�Ϳ�ܒ�yr/��B��q���E2��_�	��H��������4�+��h��<k��g|c��檖{��d6��Zֶ�G5��K�+��g��� ��>��WF�ZB8:� ��|F(�~H���;�M��� `���أ�jd���e)�����7A�-#%�����褤�*����ӫ3�X� y�.���M�ɬ}D�Er�ҙ9�9�;n�xFC>��[m����r�
�`9̱]>|��`)��L|[6h�Ix�Z��dpmC|2��V�4��hU�:ywX5g�c`\Wu���8s��sm>:h�iv���_��@�Ǡ�4�%����&�Џ��a�Fdz1��KDh��&�6��ZПu�� HK���%~�{�3O9�z�C��!A�銁��9�����7;U�ݘf�pPI���D�5i��	�"	xL~$�V��ѢUÁ�y�wf/ ��V�;����4�$��{���>��n�/a�0�Rn��kJ�z�s�η�\Y�����~v �J
kk�tuK��,�1R�
��?(��ݬr��\��z��ߺi�)JH� �8����ȿ4N8�11p"��Ԓ��1���o�1N-ŝV,~:���%��.����o��f�Q�
������['q.;���s�Y��]��x���;�'�.L籎��!,,�^y=,fr`�/�#Ϯܡ��5	bJQ��v���w$�>��%�QF�|�O�2:�ۯ��L>�������$_}yA?���ڳl8��Mk�j�/J��?���P��>h]_�7�T�:�
�	��^J��Cig+C�}]?k��"�e���"�d;۞,_�7FA��� )����i=��p�����Q�2y���(��,�_�*�W4�lO9k���/���l>G���$=H������ru�e� �����8��u�X����`�z��i�,�Ɉ�2���c�K.�m�d}��k�=�e��� �<+�6�ִ$�73���jg#�q�<J���.Hw�P��:r�!�ü{?E��1�� -e"����?�o�Ͱ5�m��s'�N<�NNy5���L��4�}�T�nHv���~�r�J��?�׽9�h+��@�X��O+O��������!� M�Q�_7���U�bȓ�K��mV,��ux@��ɪ[������ul�2���ԓP?�J��T &�2�!�" C�w�q�|�n[��ڲ8��.ߚ�d�W#��P�2?M�Q�(:!���-�B���8#�����'����y�i�kZ>`v9��*/���y�S�Qj���0��@�T,(}4l�ݕ�'�':�O��$|�@%�q���yJ����5(0��<Q7�k�8$�*����d��/7W����]���^d�6���]���r��I�1�0k�~�k�(i��*�epe��)Dtuk�Lu�&�ic��{�f��1����V�ey㙑_A��U���� I���7���\]Hq�����Yy�M��Xn1��A�p*��Y�&"�|��ɭDz���/\-[�b�j!�y\�{$���I��As=7�>2L�!]e��Џ|u�s\;�M�?j���[1���P>����k�vj�G@�F�{�����̿�֚�������F��Cm:5�o]�t���Z\�Z��p���vY�\�VR_I�8&No����8+T���Z���V��Q��[�,����y�?��h8���F�1���6��~xc��mU�f�F�K#	�UzՒ����>�|�3s��^�乳<�����.*�|ϖ�P��ā/�
j��0����&ׂ��>�£zN�3Ъą��������5
�򡪧��2V�l0r߮a�_�]��Z�q��*�|�U�<��&�H�T|y��'c���/<9#���DZ&FM {��oe"�}���Ή���5w��p�� &�ĜӰL4�h���?D�K_�$̉R霦��Թ��p�o"�����&Na�x�s���zF����^�8��yAr����(�"�o�I7���(��*�VqdV�C�O��ɟ�s�`�n|��6�4�윑5��>����I�0�:~g`w�z@*:nU���Ɩ���VQ�8Ĵ�3	�-Cf �&e���	x��$���@����h�e?I��=��P:]�pyr{�ʢ3�W�u�J�n���R�p�nw|�tՒ�/{��rGC�s#2�����fc�I��A�����!��4�k���ĵu��\+�ڻ~��Y�?�F1�(����H5:�Q�����&[��R����[���sk�.�5�]%���6�%T	�Fz�e�K����v�,��$��F~>�Б�u�U�)�_�B	�j����q#X˯�r�VW���ľ�k����I ?z)��X�ȖV1�Q(2�P,��xF#�Z�g��g6��>F�(gAqS��G@Z���l}�}e�[?�:Y�Icѻ`6I�%�����$�Yf���/۪]�����vC��l�.}�
װ�aב��h�ɪKF:jL���hD���ſѹ�6�`A�ơ�oK�]��:7�ׅ"
fx����32+�+��-�d�z�m�"b���<����¯������Ei�ET�]�	�E�� �P�����0Q,N"�*��}�� ���T�F���v!�.y'��X+����d
O�a�v5f���?��v$E{'ӱ���b���js(`V�g��MJI��I�j�}�3`�~�N�~l���Ж̐x�7�qo�t(0�:7o����,_2�'�R���V�"�f��$y(upM��{g8�Lܖ�q�pvn9���Ӌ�YB  �!DM�ʤɊH� PZ�mq#ٷ���ZC����N��XJ�@6�8�)��c�̖�?��¢T#>���[�G�4�Fa�[���z/�����k1�*�K-d�	�߹���z�&!�DzLy�-�ܓ�``Z)��NŶrd��WÑ!B�_����}5�Ơq6�����d(٧�85��s3��ODBLF�b���A]��?��`2 SATBu'���R*�j)�gGӛ@;���,z��g-�T�pK�j�� ���"f��П����H)sŰ/s��@?�y�R�de���.Cȯ�U�DS;�?��_`�*����W.	H�n�*��gMz\K{�+/V�c�(�q&3ڸ	d���6aYd��/���$�A\]�d&�a��ڐl[78D:A�?�o���nʘ��_Rm=z�F&��ɞ�3�X��,!�W�qdbyD]���.+��z#�GUm\�����P��gP�坈x�U��s�AT���E/73�sB��5��L��*�{"|F~h_M�x���LZ���ՊN���8<&U5!�8�i.C��$���D[`�7�})��l������nObj�ݩ�
�0�� .@�61�Z��ԇ �A�-"�Zw`�F8x�qY��9��.R#�GD�!���-�6����Q�װ�;2�\�|�Մ�8�p�510��1le�	e]�.?6S⛉౿�KO'����."�^
��`B��V;�~҅��/������\�I);����zf�#~[�V�}��p���t���;���������9Ȫ��U����1�d?�ᇴH�K�7�{;���h� E� ����9`z�Gn&����vy �uȷb*�����"�C��+ՈϨ�GZ_[���6��g��w��w]t9��	@��?l��8��G� �u�fE�l�D8�!�x�.�f0�7���1oǋ��o�D�6�����FC@t3��8����b�\nGj�`9��3T�*x"��|����i�R��D�T�u�9>���zN���a��:�F����z%c��5�o�a�77adϚ�%iE2��v�k��C�d���Y�P�bgs35�����`R}�T��HUX�Q���_.���v@ �q�[	5$s�ͽk��n�v�7���l<"�#9�S����X�s�E���*�Z@=KI�Z�[-���~�ؾbP`�hނ��D������C0��54�0���CA��Nnv��٣6n�P���҉����n�d���7�m ������ϲ�%@�89�:�t,���$JW5��s�`��1���������:@�ܱ�a�u�qo�F�bkc����_w�4�ci����fs-�T�O�I����Wm W~�d])�R���=E�W��r��,�1������xZ|"s hqM��,��)>���	 �l��z��8���,[���K������M����T��1��m�K��H8^��^���A�:�p�f`DRpX;��L�U�� f#W#<z�)�&O�F��� @���M��:,�3��JǇL��M�͸w�\[��Z��@�{�<��fMl�Fק,�i�U'��Jf���kQ�V�h1�ˈ�i�9�٧T1"wYT����G�ܱ��0U�?�MuIOy{8A�������#�ݙc�ˀ��Tʽ��5�C�d��v���wl�KT���~�����.wq�f�e8�:2�d����kT��t�q�뙍�H��A-z������1�" ��lq���v�A&��6f� і�{�]iNr�R���VT��!��`+�a��V� �g�\,�(�j�v�*��,)}��WM�Yӟ��0y�U��o�!���V����>�\�7�>���@�Lt�����[��Fl�$q[Q������Vߎ&dTIf����\ٿ���W��6�HPhr�K��_�ڈ�
��P�!]�4Ed2�y����2z�V�b[�B�ӎ|23lhݏ��J}2ZT�%F�&��R�C������п*w�g}������	l�؜d9{�Y�f�z#�V]�C�La�*
�;����?B�럇LdOY����P?�s���(.��T��f�&�p����^�]ohv7���~�� �PG��W$��TK�.���s-�
Y)����<������X��U�gA�Yj.u��M�K(6c�ܰ7��|I/G6;_�ߋ[uq��m����3��aձ�Ar����ڽ�Y/��k0'5�>�(�t���w�x�b\'�d"ŵP-d6��B��s�,��B�A[�+�6�����T���� ͈#1]����sE���g���<0�~7ۑt41WFPs<y���K��$�`�SK;��|zᵢ��0O��YGa�)��;a*bͦR�Y*�_2��q��٩�p� �Nw?z��$"͠c\hL�US�����U�)�ejd�j g�ޕn�Z��L8m�	TÇ�89�J3����E�os�ߝ�u7}�M���̧�)���8��,l�˯�f2�1l���҅( �>�=�
U�C���w%7�ň՝ h{|/��m�ᖕ��7��k��&��1s/<md��;�|�L�U{�&v�F��8�-�\���"��	A���ek���߳>����N��a�;f+,�����&��ޥ�q������InH�B��p�Є��0c��X��Й^���v�7�`:50k۾/mň�_6�ԣ�!��8j��n�+a0ô��	RJ%�$0i35�̢�� ��mĴ����lMJ�{��F�̫�����-���E�9C����c�c_���t��7�(��wq�´�)=���wQ�S�,���h�h�v,�Տ`d�[�����6�[Ջ��X%J�'G��R.Y���f��{�݇�K�R�X�utT��]<�P(�	��G=o���A\���Ub���[�$wTY���L�R�9+x���/�_�����>��Ze"���q;W�����E�c�[��<��$����z�W|��v67�:��/E��!����`�I�ӫ�%1Q3]�D[7I�a�[��b�Mt�S��v�5�y�V7؄��w���i��
ɞ����t�=����13`�Z�n���kĂ��}�oH`]��/���>��#>'�n����;-&�>��+�y����Ks2O��!�	r �&���J��C��&�ExvZ��x#�9���؋��%��Qv��kV63"#-8à�ߓ7p7`E�s����5���]��Q��M�����u���f���[@Hq�{�kg���q3�^�r�`���(���޾ # ��3���K�f%�%Ok�c���k��c8���MG@N�3�GN��&�E+����طu$����=*�L�NŐ��S��6V���FgfK����gM�� qob������a�6%���Yd!-�l��W���7m�U�k�=����Ꭾ���6Q���M�5G�X��/��)�04�n�0��%M�g�rn}bu�q�@ۦ�gaF���L�Q�1�K�]�����2��k���:�v2�P�*�V�A�M�T��Fi4�+ QZ����w���E�4��4���-�t�L��L������q0_ro��o="韮*b�"�/��)�#���1����uB� ��9�V�"�h0;���B�Ԗ�3�h_[�sp��>�r���x�U>�<�6׋'�ӊsC�OJ��:���M�ա����@fS��G��{c���&���r�qH��D���mG�C�����QBV=ˡ���C� ��g�$JĊ2��0?{�O�ߣ��T���12�L����»� H]���Y�G�v���ְ���5_����1\�N���4�'�Z��~��� �lA�َ�(�!�XP���uB·ݶ5r�Q����)i<(�S�"ͬ[9�ܦF��tM�d��c��˳zV��=��o�O;	����4%��ә]��.qqY%l�\����S���2����(��C��cSг���)�y�!�Y,a.N�?���UM��ʵi����^�#��C�?��ruU���Y���S1 ��|��_	j�a I�2z������)AE��=��t�)�*�,*�VY�q �\U�bM��J�گ7�0�̈́4��g��ex�4���$"$������3�fo�0p����Zӻ�^��t�5�FB#�|kӶ�B�2 i���y��I����6�o�B2�))R�gm���`��h!�R��EM���i��a�':]�o�iuU��ф�ۧS��������P��KCdد[B�Xo�����/P�Ž��ơ�H˹o��Y��b��� �DެmXI�F#�B	�[g8�����^8����hg�-���Xu�ײwB��޲����lY�<9#p�<�
��%p!��J����D[���r�����|�4um�+�b5�SWc�L��ә#+]�E&:�"���M� ������j`��Ye�S�����a'
DCy��.�gcZ�: ��ǜ%k��P�p59���9T��g����tdA���[���@j7�jVL`D4�^l56Q�?�و��-5�m?����N9W�}�rǀ�o�?���m3
; ����iˏ#CX�`&��1r%�#�t�Cj5\�07����vt�R���8�l#'3�)��* �^R&,kfK�D�9<�
J�#���Ȃma�m��XC�4h�<b�Θ��4�O�mI	�_�BWF�?�!���g�3�_ء��hY�O���̰q��]�z���tZ �QC�5�
n����=|S�;����\��`lam|N�-A�f���>����$' �Ե:RT;Rp�c\�J)G���+������ߪ$[������ҧ��D�s�+�j�GԴL�Nˬ��v��۱wB�>��B�ʌ$7�:��4����F$���̧�W�Q�uN�y�ty��M�5�R+S;�6~������?�a��x�ª�4�V�۸�L�� ��a�ݶI�K�Z��+��}܄����1AB=/�h�O�@����:�ǂ��7�#o�{K�yU����B�T=�R�B-s��e+��q-T�z>{-S%=�F����EfZn�b�sϭ~��U��1Ugc)O�N�L*	9�8��tV��_fq}gc���QN�f0A;Q_d~%��	<\�-�Z�=O�G\+]�,�h�p�b)�7م�G��U�%%�$Z��:�nA�a�U��]�CYV�~f�9�]8:��͒SC�g�jñK�4.��Qg�o^$�bHjF�l�uux?�V�~�&��T��_ryp��%
}�F��ol�S�d5�_xW�%=m�y���x|e3la�r��Ter�v��|�t=ݥ���2��2��\6�_�E�Jj������zL�]�H��L�:+��B8r��V���uَ6����)�Iư�M�d��,�Q�ʗ�I�Ҙ;*��ty�'q�2������y���}�Vs9�T9������帄Tƽ����&�zZ.��?�y�Ht�!�O���u���W�#[A�l)��A5{�Cq���K�\�S7z���8�����~9J�G�P�?�\C���¹��7���N��SD틥3�:>��~�M� ����e���$�f8Qv���K�� x����_�@��.��Q1�$F3p��p?��9w`�J��h��m���DD7�w��Um�|���E:�mjD�	oJ���t�Vד���@5t���"�Ʃy&|&�tQ��5%��
�C�T�Ԑs,0,@�G�M�vK3yi/�$m$?��^����z˺�x�ov�b��Q�0G����b�e�j�|,�i�5_�2��$t�v���Ҙj��Q�*�s޼�L����n�����G�拰-Yezt9[:aZ���p�S�&v|B�>	�
��|@	�K��R�`�} �H��	�?���ڥ�h"�kLi�3>|�O$�yPrd�S�d�b�)M�u]�B�A5��:�������x��k-�n=���w�ϸd�XYL�S�5��,� �@�~_�p���^�X�(�F$�(JU�='�G,W!���U4�3#������-��y�+�< �W����,�麕�Z�t��
�#�zE�ƈ�;����*�������V�&n~z�;A�P��`�TQj@7��.^HEڕ�3�Y&�7o�4~�l�0�#�B���Bf�Uܤ�-�� �!=�n��p���6mň)q�R��C�nU�)��w���0U
E�\�zm�%���$N�����t��@4*��05aB7���Px!i6-�����]�_�f1!�q��F��pܤA�҈m�c#���2��Z�n�.�'C/���r��<�=G�:�[�C�c��5��1eq��i} �]��My�!�=����[�Ƴ�DASjI���*SxP��YצgE����V�('F���|���^bŀG/<�e��6	>Hv�&�m6���)�U�>�-:[g�I �۲"%���������@�l�A࿒��[����%��#z"�#�t�2,��U�ϙz��g�F�DbV�$�)f���K��x?������.\#T�����\���ĭ��<Yl�8�]�����V�o�B��?`F,��{ �b�s5w&��3��o[��G/C��¢��S+�`����S�G�9���N���~�|��o��wii�����c��gg�&����i;~b�c�A�����$x�u;��=��˫�� ��)�@�poS�	<�5
V(!.'��x�Ȉ@��R�
�2µ�l�<��[��k�o��F��/���2�ck�_	��`��T2�"a=��M	kp�f�2�W�ǅ��!�	���&��_����'|
����W�������|�����/s��5�����n]y?]�7}ؠv�\}��'@��nX��N.~*�k�;tP�F����⅝��c)�0�������Q���LL5t���;��8(�e��B���
�z��c��Z�	��=Z��K�*^��-Ƀ�hT�����U�@&r�,��1;m�ޣ*��WQBB�#�&_���Kj|�,i/&�,�a���y	a�h:l�����$��t�B���F��QW��gG�T����Wy��Fw]�ܩ#}�Zzc�Җ_�#�N~�O���y��T�ek���p0Ќ�N'�SK�2�t��f �)�~|��� �a��i�zֶ��zNo��}
�.�F�~#8����b%hZO�o	<���X��VeC���UJ]v*�kVc��a	��\�^R]�����U�N��ɚ�h�6ne6@��mgi�k��I��}�	�h����Ne�F=40^^j�,���Ɖ�sX[�g(�7`��z��\�`�2�AOdO+�މcq�7��#�g?��#�\b� �Nd>-4������k_�|_���Sib����nNn���6��1mC����V�Շ�I|�u�.2N��m��ip�S3�ux���-�+�<��Ru�k�m�<[y����%ru��큗6��>�ӊu; ҩY!T$�v�ƨ���7�:6��D츂���1�x�j�I�T��f��j[�Z����]�/&����; �R��j[��1��Q��i��⦚���<d�u�<�#<�^#_����G��.�7�:�@�ab����d�_�z>��	U�Aչ�d�ϐ����F�5����5�M�������e_�����B�!O~~��;a�?P����ٴ�.^� ��c�O��ոB1�pS� �Y�f��G�rp��/m�A���e����>������ ���d0�~,>?�L��La��"���6�	?�cZ�P��Yt�E^�77��$���'�.���)�-���!�"�}\WI_���#��'�e�� H�@�w��V�bZĶ/ii[���'7�j�W�X��Ja+VxyH��84-��z�!��>�g@�/��ypz�:�+��Z!h8�v��s��#�wklj+D�>��7�W�#I�<-t���O�.��w%2�H|���]�֌��Ghy���3V�Nß���e-A��v��t�����
je�� 8�;#��+�NX�=��*K�c��bOv�#���O
�:��X1|P�����gC���H�\��xM �y��D��JH�?�&��Y	w��ҜY=��J��Sb������k�6M�:��3����nv�!����Oq���R�y�j}��z%�6@S'Ӣ�A�}60:1ُ�����W!����:q�\t�/[U����R-����S�sz�6=�|�����2E&�\yx���#uRr�?�!66�L����<��#�h~�����w1d ؛���	\��#jĂV��D�=}����D�S����\��T@��\e��ܑ��:�`W�82=8��W6����#<
�/\��Fu�$L K�k�T�6��]x'�-ElO��;��)�[%P�M�t�s�T�:]�=�9G�v]���&�1��_���1v�Z�7;h�i̽(�oīg1I��-������?�Q���&�y�I�/Ϻ�鳓��3I��T��8��sFq�Z��Hi��S`�"B��~�I�rj�ў�	n� ��Ѷq�l�Ѳu�2����1QSL�-�Ԧ=�_�f
6:/[�q����5�Zg5ՌYVA�����3�`lc_�dڈ>���i�����}	F��>��r�a.[� |��
��t�:���9�D7��Kⷅ��
JaUμB���`1@��n�y�O���FN�*�kT%�Z� ��&���\}'��=9:�����}�(�,���J\K��e�]��XjM|x���,�N?�nv�d�V�}��l������n�BM�jH�`��K��N
>A:=�9U�5֙;��)�h����|;J>�x��|�^�5�o���	�(f`���L��2�}�h���GQ�`n�`�m�c�.��)J.K�(�{����Q�����O�+]�qt������a*�e�&7�b�v�?a?�����P�	Z��~Fq+N�c�αP��`�u�A���*��f����F�r����.�JC�$�w� �y���D��|j,k+�ŻwfL`j����J�+�w���ۖ�᧫�� �L	��`�6$29�\)��:'U���Cx�M��fU��<Yپ۩I.��[oiw��o��;�?��¡�*������5�ڜ�b���Q�n�D��!�P��{ER�;���u�x7���di�&�~�B
.��	lz�w�oՇ� bxw�V�@I��;[�^�N?J�8�0d�$3�^�X��v0��rWV[Ћ�	<��#�i��Z1���]Y����y�����_���
($K�טJ���C$�z�Ws