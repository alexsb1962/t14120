��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�������*p�8�[�e��)S�Ab�C��%Ɏ��$��?�����.'��|۲�7��?f��O�������#�9�+[�[<��I^��3�c!�g���]��/�k�<p�5��D�ӆ�p��'���RD���mm��>�M�|�K��d��UT΃׿�!?�7|?� 2J��,;�
>؆b����u�!����Sk��,�	@�}������CME��w�������pb��ϳ-��x.�M �5�|������渷���O�ډ`�Z

%�#��^XR��*Z> v�)|q��y�bЅ<��i�x6�H�lCٕmΑ��,ԣ��i0~i?�H���3�f��H�aa^����+(�U�����AK7�Q��o���#��9bwj�	��f<0����|�K�����
� ��Q�w��q;p�$j�5�5�v��&!�N�K�NA���._m����(��.�Ws`"*|��8(vr���Mt���� ��sF%�)��b��uk�G7�����_w1_M��4�(%I/��{��G7wr����{�Tz�����B:�u�6��s��/�ZJ�^�/��E
�֒�r_���٣�O�p���O���|��BT��@R�+؀�@�;���Z>�������LSĴU/�T�:褊�MIt���-jd�$p��	�0D�	l���W�OFըi1z��)b37��]��&��>PZE�MkLz��Xmw��K�2�./ �_���j{��u'�3����EA��M2���٘H"���CV��Iu&��(a��R�t����#D����]Dd�6��Z�Te��C�wp�ڌ��^�	��%�D"_K��fBÆ@XT������
	�t��C�G�!k��m��~��8�[�#����U��,}�bF��e�k��>Dj!�؞H��	�bT�畣�m�2x��b��Jjj鰓�)�������YI� U-���$�4�n�����ȅ]}Sz�nl�f���b��B,���"%�$���Vnϡ�6ɶ3���Θ�N[�`l�`����!lJ剥U��>Nec��� w[��^(���DAN�)�� ��G(���T>��D��q�1���<�� g5������{����(XԽJ���{�j�MeP��Sw�C�|O�[C��?�$L���n�@qJ����4��j�.	�$��[wXz�T`�� ���dGE��ww��&?�l��%���qqx�i����.�x�D!S+�~;l�Bk�u������z��ǃR=I:����c�t��#���m���5�<�(
-��(�sܡ�����̌&�Yw��ߪ�&�����|L�d*߹��mp)UQ�{_gJ%��s�=��V��L���¸/��;����m��pVL���JR��J��s��Y<��a�p��a"A6z���`c����O�~��Vo�N�_L3f�FQ��5T�����2�R��>�50�IԀ*��9�ah���e"�9��ե$�l�y0��:�j+i��i_����d?�BW�ďe#�w9��\��LF^�˳��
9u�$��0�"����ó�^� ��D�lE.����̞��Ս��+BG-}D=Dm(�n>s���0P��,����$��K��&�\`�K��{�K�h�Jt�1�-lu�4��4���n�rH"��~,B�ΒGY��V�=����[#��cե<��� X�8�ˆe	��F��p�h�54�HfK먚ŭ5Q_��(R��G�����M3�\ ̷�ZE���4�����auE���aA��j�ĨY�"�o�!��xC�`1J=~���Ĺu�+����.(����)���W��4�y���_Aӝ�W0�"�����i$O5�B���P�R��Y*UD��[p��_T��J��0�6L�'m�3]"�6S���أ�0��M
��bT �&�;ք����a����Ս;��CcAu2���Dv����N�n���oJ�̛G&�*�I�O�ƀCu��(v>fR��~� p_�fo�W��C�KP�qH�}#ZP�
c�:+��.���f������m����,�Gs���L��cl�#��_�A���;V�~.%�O���V� ����3�f}�����q�v���f�p������$�B����Z���S�+��ގ�p4�y�a�
I��(���ն�ti��6���!���m��� �3�6��n�	�:}}�GE��c�Tnժİ{�¿..}����n��,�~B��y��]��=᥶�i��	���|BOGe2���;&Q)��?B㕘��	؇�4* �Fa��+�<������=�dg���]R��<b�8�$�X����
w����f���@]�n��q�r�/PkT%�*���d��ɽ�D��/���3M�^voYhBʞЗ�t0[3�1�#�8g5�Ǖv��6f�(+�x1\������"�\����A�a;�U#;y�}xэ�q�kX̢qO��5�u�M�i����g1��z�'w~�}n[�!�v}�9������1%9s�`Kv	�4N�aW4�(F[9Z6R�Tq��%��?S�_���H�yh����Z�;�+V�(�ۭC�f_�B�`�+���zv�ǚ$˝'�q�k�1��!�<i��Ҭ�K�xO�!>P8|^���S������4ȯ@*7����� ��B&>L��������}��.-�>�ܐ��x�`an �7�T����=l-x�Ȥ"5��D�z�v}J��J�t�lL��}�KZ�b���+s�����"��9F�9P��G��&7���|�XD�єʏ\r�Xh���;~��ZE� �b��-b�@��6}7�0�h>������j����Dy���H��PNg�t;C�IV'��P('�z�#$?§��S ��㕢ƅ ð�4�5���s��g�D[+IZ�T�H���<�c�_j����������с���<����	 �y�Rx[�����]��0,/����<�Q$����M1��zң�.�"u��eΝ�`M>IŁ��$��sMb�1��ێN���wG�?����&����C�@$�<'��Z=j$ �?sH���{VcM�<�S�K��P ���&�R|�=[��4ͤ��5�B@xD��O������Џ�pw�U���@r�8�OŪ�����F��x��|�P�:q�=Jy`OX�A�U��uj��'k�:}���K��㞇<_�3�7���q>��F�qJ�?U�7�c�=::&u�/�I;���S��5q��>wo��ز�G��&�a�p8HX��A��y�^�f]�6����^r�T�-o���5,T߽	�&��	��ITt`-��1�ά����l�����HǞ���J�_s�;�:�ap��X�j��m���
;02�<�����Z�c��>�!�Ln�H�T�N�y�F7���THB\^%�ALF$.*Q�hI8p�����+���als��Sq|���!�$g8{O1ĺ����ڌ���Vnx�tȅ� ��7�4���o%O��[_)!1�)۾�EH��LL^k�������yx3�����l�b�>�2��3����M0�@%X|�w�]���н��u,��K���zM�28�܍Ɩkk���P`ȉ¶�4��(P񬅪)����3)�x3�w��'&�V�m�W�ܸ��s�����x����U�=V}`eׇ��R���r��gKaķY�&Z��i^ވ��a�ҙ
��j���( �g�I��k��6�G��	�+-ݟM/P}��h�c��!L��-P2��Œ'��U־-�7c��2+�x�Oݻg�}ס4_���A�:�A]��� ��P�6�Y%ȝ�F�r��+%�r;Q~�j��&x��)�3bͷqAi���iL��5�Z�c�:Y�ZH!)ruu���7XL|���󨌅R�F�\��|�ֈC�E)�'d���
�q��T'�]����I-�;;=���εb�q��I�%�uXV�P�|���+A�^!�� ��9[�%-^�
9ŶP�>ݘ��|=�s)`�E$9�D����a{����7���\pڞ�s�H���`E�mm`�9lW�f��ș���/˰E�=�X棰5"'r�씼���!�)�FF:�/haOY����B�üu�K�k^������y J�}�ݲ�\�Y��x�R���� �uSU�2M#�P��Dl�F�Y�2y�[gc�A��'���b0�.MB|>:Æ
r�}+yS���L	л�C0��*|M�D�x�Dm2n�[�U���&��Ff� ���%ـ3>һ~8)��ջ�V��7J.���))�ɍ��7��_��Iw��w�y�/����2��
w~l��g���a��ײ*@E����}f"�4P|��_my��#<�֋�[����U�2g�o\��z�,ݎ(e��rh�6:Y�k�
9	��������.�1�
^�AI؟�/�\"�հ�%�#��F��kbH��|z�����\D�)�uR��
#G��'h�Ļ�F1ވ:�`������?D�O���l!t�Q!_Mp�"�8!�C9Q�v��E2_`sJP�Z�q��xPNjLn��e�u�z&�k)��b�3�e��H���&��@`&�k� *�~���h�`+�#T\
�TTӁ?I��Y�.�=�e�1H�8���H�u;��r���[�Μ��Zb�N�*�r��>�-&�2]�	���;OB��m'R�.Xm�zx#/8�[��̕��!_�[�O��1����T��hW�qK�����0��Oy�������i�uL�u��]�wٔڅ��w,\?fe��y�j���1a�����m8[�\�$޵KDZ��	:(�A�r���m��<'�iғH��� O�
i{&�h��`[V��ZஏW)UƱ�Ow�t�<5̠v��o/r��W�;�4������FFPRd��;p@�/��sa�о����N

�Mo�˒��.���q<@�n��^t*7,�˥O0���}��Is�g��zf6R������$87���y����(�ײOث��+ŏS�-Y�����>ez@��N�\��vm��3��?؂�^���Ӣi':�
aя���GL��y@�n�P���O��A�Q %)&1��,�(զ�aF�z&>�c�]7̟*���wE��Jw��/����|.ķB6W��D����>]u�C�d�rlRt��&�8Twe�)��$���|]������X�rV!�[�py�\�;�̜�x�Ӵ���uƮ��=��:�h��s��jF�^�~�:�e��U����h@��Sb��T�5_�.�����w�R=Rl���E<4�l(A�R ϔە`�K��Os�~|��'�,�N����U{���d׎ �l�hml�1�i�D�v�W��3�s�Je8f�m�=�W|�H[�`π����l��4���я�g�B7l�:�:ݷ�^MB� ��K�I�^/7Ðr�)�#Z��Rc�(�G\P�!!qn�����`�i=m��C�2���1� t�Y��*A{&r�q��O  
�8�#�l����Evdl^�x��Q`v|�U^:oG�fE�S��Pݜn��#��_u@G����ѕRZ/"J^pֶ��CR`W.<���f����2� �;���qFN�p@x�2Yq�
C����A������i�Q��P]�aAF�٬N2�"\�x��nꨂ��#�5&�"�M���Z��i�S���AP&�/��9T�)Il�dV�Oa��㝯�^h0�
�I�L�VE6����O�����ڬ;�gPb�kJ:�f�gT�dFUQzP'��I�] �u�=�Ɵ&v-(��&=���Љ��^�`��Y���
<�v)��n�С�U�3?��Y������O�Q�r�����7��ϫ�;ԑ�-'�%��yo�C��v]�VC�l%@�?,��	s��3����a��ȉ�
#����z4��P�%�v��[��յ��i��~"��q��Χ.|/%E�b���`mq<��j�s�(6#o�S:{�����L@�b��X�b��¸�pp��7�vZ���������h#2?i��"9+���F��]"�,�y�r��z�d�)����1�S	���y�.�;]�����ETp�3Ǧ�U�ӈ���OU��f���R1���d�'��Ӈ�ʭ������.ت9�����
��a����R�z|�lČ�c�S����
<�PHY!��F(�V�O[�M�Ӻm�7HBn6�P¦!���V��/�ϼZ-���!o�'�����$��b�d��}=�����ʝ'�\�|������՝�V�ji5�kv��$��pN(�]@9�(����Bq�uLu,���tP��Ya��J�*f��S�A��y���5p���'���uˈ��H/m�4��{��[��_�e����-�_G�).�Q;$��_�������}D�یe�[�L�Q���j�/��@���"�;�" Y��.(��܆Ѻ���e������[�ɀ�~�f��A�ޞ]���j��"ع�'�Z����c��4�D��H���7s����U/;�YgBc_�#�Cۜ�"��V�Iǲ�nf�>����WLm	�\Ü�/>=bÔ*�,�X3C�&p��"�ҭ�MH`���H�<E�n�j\�TǑ*�8:����E)Q�6��a�D�U]���׻A�.ޔ))��:��>;�p��剑<-�;�;WuL��`��9�Pn,��;!��ԑk~�"���ن*�s�u��*~�}�t�˻�+*�P~���'���e�K�s�0�ѳ�>{����?*�;�+�=u����=���ɃƇծO�A:����wBK��>~.�����g �d��ȗ�4_Ԥ�_��EP���Ǣu2��$��ZY����R����ƃu�o%xE�L�M�̇D#�CXZ��:�@RDw�)a�d��%"�z5T�X[X�ނ��^�sͿ�����2�Bצ4�+��"�,x����A�ARL1���4�
�Ptq�-K��_���V�L�����f{d;����Cp.pG#��e��]o�ڈ��H펡��'^T^�&�4�gǶ��+? 0:�=�Z��qk�^縯�ğ	��o�7�ݟ�뛖���MߪLa�6+��礼��&�>�����DB��� w��e�ۡ�	�2��d��	��)�����.gA/R��^��8�f_�,de�"���'�������{�Z鱀��"ch �o�k }[�}O݆s��0��Ḅ��C�W�������]����o��aT�{�#�+M� Ε�VG!��n^T�>=��q���_�,� zR�m2�Ȣg�����0/���#Ԩ����7��_��@�Χ����?�uvk�2��ä����wW�Ǭ''���	�gK�^bj��|霤n���ҟLU,�cv�jZ�r��n6"���3{�pC�a]��p��x�-�"l<�Z5�~�߸�&f�vٙ\�O.*t$84�I6�ޫ��C��MD��.����J�7e�/��iM�>W�O>z&̍����=^�ebѤ���W�hUqX��5ZPd	�)���⽄kY��6lD��L���#1Q�$o���U[��� �O�gcs�.����)�;����	��p�O�	WHC%%](�(���8E��9#m�V#�7��n]���1�|8L|$)���ؐ<�^R6Zy�#\6�c ]5F �5E�qt��O����KH7��0���+V}�Sp6�;\�n~��(ӻAB���Y���6;�f;m�6��g���G�2���HLoԊ�=���_ ������-��!�H'Vݡ:|s/�	�j���Ε���pJ�|ݝ:��'���-g�<�Py�E��`�c���yQ�H��!ףG{R��e�%ɚG��R\��&���ثGS>�W/��֠�-�ֶ����"���,�ty�A��&���_g{�BC�����H�Fh�L��Jя:kc>�]e$�k��M�J����҅�A�+`(�h�J+ �^�
t�ݢg��<w��8��4�H�s�W����b:��,r��)id_x^�lzx�I���3�Uy����ijq�|�ì�1�v����ݑ�}1ޜO�O^۳.|�\t����vǉ����yW;�!�qbѬi�����FF@�]��'Q�&��=�>�'�|��aL��Z!���t�Q����%Qwh�oe$�7��5esB��GͿ�T�N�E5ޙݞ�����������+�<�U���	�Ago�v��A��x|am������xhwg<��$�h\V_)&��E��]̣z �̹�?�b�qh�>��� U�p�.nC��מIi��uo�:~W�+��c_����|�i�B�:�vxOT3R��(�N>���P�g�NR�wM��ח۲Q�麘�J�%`o{ӥ�U����G�DI�- �}���J��$��Pm��v63�n�Q5ϧ���.!��9��s�u i��u��vG�-U(vճZ���p��k���@�.�
5K�"��g+n���T��q/�gUqޯX�����Z%�]EJ�I�1�x��Ļ�af"!��<sbЋ��t�Jx~��C�4'CW���Э��t]̹0)R)��5�CTz ���0� ��itz�V�R51�N��R޶��+�[�SnᪧM�O�����\��ѿ��L����y�a��ѭ	�B�^_>�A����ހ�~��ι��~-�\���G�t�����
�Zv�3�&>���.�qi����}d����θ����*�
��',�3��B�w�cH�Y�kg�տ�7m��L�!$gC�B���k����o��M�X� �-4�~��t��v�C
�$酉zړ(�_�i�˧#MbpT-�;o�&w��}�F�q�If5qi�����*�	��rL�I��A�c�(�3)��"��D��Q�W�H���y1%]<6}\�#�jj�����/�;A(*���"�M6o��8����4^t����}��Y�kN��4??�4�U�:�v=�)�z]P�v��cfh`-����T��x��JC8�oL�T��}h��x��;"K��N��/#��4UER������ѕ��<YAȿ�`U^�Xl-))�Lq�^��Ә8�.�N�
::�37%{`�NM\��f�K;X0��紏(xNmQ_���'�K���r
���:�k�g���0ƿ��M���n��b�����Kst���8�������Z�CƣB��'��ҿU�'�����f^��Fs�]���j����D���\U��霏мZ}+jc]��D��3���M��9�4�7�����G��٪5�]2\ʟW\�z�=����S����#�011K�	�=��:�8�~,�xz|��� L�(�����A������2��Q\�f�L����U����i�>��0�4j?�pz���u�8<�ES�Z6��Q ��b�]�8d����B��=�R�F�O�.�� 2�?sH���D�Q(ch�t���g�w�P�.�9.�=$0y���N�F҇CJ��Cw�GRȉTDUO7�}��h�e��������)L�d���e��\ ��nK8CV#7�q�ŋ��.��k=�A1�Hc�\[%��P�^��|9���c��3!��dNF�Vk$�5}ыm��b�;�E�<a���ʈ�}�//-���k/`�e�mj<����9G�#�1VK����ln�Lz�C����s8��/\�=�c���sR�~*K�߀����*�ǽI?�G|�ȕ����Q�S�s��zݟ�4 �� ���l���vX�A_0[���(��=�����#���χ勫�8��v��/H+| �a������~�e�_M�w]1-�� �^D�֛οiw��+�A���o�@��pG��dM˂@���(	XPI{n%�:�_ݳ�9��k�mmGZ�?���W*v��ۛxAyj���x��ne��d}��"oSt)��WP;z�
ZI_g�
(�'3��t����P�X����֖k8�a�71��B&�~��U�]/��ͧ�7�b�e��r2��X^Բ�!~���&�(w<�gҋ`�MCK�f���p����Y������MO��KS����h1�7�Ф?yjvB�H�t�sY���A�6L ���74����ס�Wi�����]%Ymx=���N�_��T����r�������c����+l�@g���~��ˡC���ֻ�;U�,_��,�
>�E �!h��k�#<c��~.9��u�D�������[�1�䷍�_���W,�Sv��,���i�Zz6���3�`����fD�<����׉�Ҋ(ct�ڡ�WB<=���������;i(��2��0�%�1��n^�"!�O���i�#�J,Baj�{�47o�&w7��|�Q�?������P)�ރ�%m7_v��U�C�${#��XQ���H$;��y(�?f�1%�|�sq/7����~�q���f����5qP�}��1�$TV����D�q��ν��4�/(����4C`@v���7�i�`F-�����bm��%��cN�%�{�V��lx%����Ȓ4�9x�|�V=�$�����
c��nS���ʩ�C�}�s�s���+S��kS��uy9un3M������5��:u��]'.��*J8G�=�h}o��I�����\Lw1�L���q;	���`K���)�ON�����&����J�#oV�DX�L�)�m\�#Dr���-܂7k���6�.E�aJ�.�9�ˉ# ��H���ҀB&��)���FL�15[4������%���Z-3d�m ��Q�.�'�!�}��[L�a�������]*�w�����O�a����k�D�g4��%�+�{�/%ǺL.�*��� r�_��S��]������q)�U,�����?.�� 
]��A�+7�k�Z�lֳeB��7X̄���w��{��_�]�sa2]��-I�q�t��d��u��>��'��d c���Kfy�cg��Y��+-�x$�`ח 	�k��Ġ�����֥N�;�N���I�Sr�k��{Sk��V����
��"�<A�`Z�K���G@7Q�A�f�R��Ed~1�8�ܟ�t�9��Ị@�1��Rû��������@D�mo��Ѭ���nH�N�����W�ANI����O�f�bY7��.	B��y�o�F +\����=��$��sYb@��jq^2������cq~'�huU���{�b��#��^�R�OѦmPI���T�*0����0sN�:��leC�W?�^Y|0�&)��׺�|�yś4��62��@'�]XڔWs�kؒ��k�ˊk��|i���{��_V�˦��T[v�jk���
4d0�=�/ 涠�xR�PA�ўP��uΠ}KA���qO�&c�$Pr�5�&1���l��5����S�2/$���^�$�mM��)�R�������5׭5�SՁ1��(d���R��s���(����s6±5�(��|���=��Tt��E���E�����řeO�d�9����H�5	$�L������#@�`�	�T��D�3HPu�Yi�To�M�0�ॗ���UiΫ5T>��C1�- ga�|�ڥ�W��$�ɝ��̴n"̛�u�>��,i�E���~�m~p�i�@�"�g��`�����!y���VBv�M�-���W��b�?��:�!ot୹9O_o�M��t"�hq�l�2y"	����e=7v�9���w�{E_���ˏXg�esLP�m�w4������NugS�I������H��2���m�qzt��dOq�?�j��l��5�x2�p6�Ҁ��^\�d�8�H���D'Z	�+�k�8��z�T�?�`���\�Â2��`H�̛�+��c̦>.rެ�l��ɧ�#�K1���>5����A�N����8�K������p<��#�YR
�.��:*�$.^K�޸�w��}�T��{\bMh�k{�a��3Ӭ���4�4�)�>_3ǝ�_�4�rCs�:SE�qk{�
�Eu-ce¢��bD�2� ν����˳CF��v�+��m��Ѳ�O�-�F񾵮�Gz[h~���\�U����L�Bg�Vo;�ޮ��%�����r1°ayvP�ߜ��І��21؈��>_:�4�� �H���չ���O^��Ǌ�~}���>yx��^ѕ�؅��"~xmLX���0�:�%,B��G�K-�/���j2�<��ұ,"�ޫ!��n��5�M ������wM����Z�o��� g�2�������JfϷ����x?�TdOn[,���<N���T�p3�FzK	A!MKs���?�YkH��4`�|�*��L�^|��QV�:E*�Q��k� H���ܹzX�#�ʹ��c��f�-� ^v�9\���M�p�{�^�� �=�֎]zt�X�U�p8�������	MBu^���M�0�) /�;�x��J�N�?�9I��f���`}j�F�t�}�jk��'��L������O���;��Sb�+r@82���а�}�@˧�_y88p�,��`r����NqfNX�>,�;��g�]�� �^��Y+�˨?'&R�-xAO�����O���M.�	!Ph�"� l;�B�������'�������b������t�->�c��,V������,�ѻa����+�#��LG]ʈ2 3� �U��+M�NxO*ni���*�SZ�j�Xte`?�#(��2d��Ƒ��	<0��Ec�i�I���c���iC`9�.æ4X.�[���bͶ{(Q�Y��L���k2�g:%v����Ξ �˚�>z����B}��Cg�J>��BBe|�$`F�r�~���h�e#��Gmt��6�6Ǯ�N*����QQ���wQW��%�f����`\�C���]�� /���6-�5���{\w�m����>��p�jT�~�tt�/p�{���bv3#c����{��5FP�L(8P�*{��C�d[�y���"^UP�����D0�Xv��P����i�QTr�O"�G����~kg!��x��!��5s���u�`[cF�F��Ѥ_�d\i5�D5���¨V&;w�;�k�y
�73��K��C�JH�����[�Rڕ�Y�|�Sr�7o�U���yFE$ss�q�'[�<�.�8��+%׊̸.�Y�#ly�v��pϞ��B�����o#Jt��x�J�_�wxλu=Z�Z"C����<�Hu���1�����Տ��)�3Z����0�##��Nh�,!B�w��!�v7.A|�8r�E�L�F�6UI���DyJ�+��XP�K����:�;�<�1�A/���_XCKC%7Vw]"g���юj���F3QP�?�Kr��Ec�V�5'��t��JRۇ\�QK)�ծ�Ӧ�
�'���K��t�:�� �x�>�G�\�������r2��`G�W�(��ο�>R�}��k�nhIL��VtL+@>��kc�dI�
i�>2)�g��Æй�&P�O఺;��G�ۀ���G�^��pS��H=Wz>��i�o����"��c����B��sǘY$�����%pbJ�	Yͣ���l�;W�}��1ԥ.���Ze�z��V!
2gȕ�.+��hJAj�)����*}c�0�9�� 
����T���Ƴ�DK�gօ%��bZ%��p��榹��ڀ�Ꭼ���-��AO_�`><)73��2JՔ�Qm�2���ӵ
�SD���[�q}�j���f����W��!�#]vû�v����ư����-7�8	�i�H*%�]]�d�rϚ��2���jE7%��a崇C=�}�n���^�2{�:U�2����y�H?���(̶,�)���lL'_�K�M[��!�Nz�Ŵ�R?Ë�?�4�L7YZ�O*a?��,�cx�M�HC�K� �j��<]�A�Z��������>ܺ����	�$�Ա{�ҙ�<�
b��u�4
 ��V9�@=%0U
�34�4�I^�lD�\���S	^.P���,K�@S*�/V[��4m~b�w;�߹��fԷ�3
�rfFZ_�� �O
]=m�~�\�C,l�q�2����3���=ߝ#��d��(N���eֈx�l9��^G�~�b��[l��P�`�:�q�j/I�nޘ�J��.`q|��D'�Ѐk��S����fGϛ|��ǹ~��9����构P�
���We�c���!4	�M2������5�L9� ��/D zg]-1\mS^h�5��ǡ���D���g%�c�������Y���A�~(�5q�t��	&�����?_��5�Ah�mk���K��Gdf�ur&Q��ı�(�LH��c��	~`�������H��)g�Ð�P����5�~��V��Ԙ��>�l�1&�1Q�ӰΟ���U���a��8c�}D˼��"�p�ޫʚl�(L��,�r��p��gJ�1���,�.j,��e�:jpvU ��KVx�9n�!���Y���-��w5L�y��NYȼo�������r�(�1�cjd����.%2�i�>c�o-��ga�����gboA��큏��pK"�Mg��xVd_)��F��a$�QW[��"eD�7'ۈ�������4v���8�HJ]�����;L4��b��sr�N�ō�$����'���x���	'{�`W�X��b�E�ҽӢ�X�a٦഻E���qvj�N��x\D�gRq֩�|��_��)#,Q�=.������i,ݬ�rq��&;��#�].�h�E[��b����0��M�?BxRH����¨��+߷�s���i�*�.y���l &���3�>��0+��`B����>~��foa� �j��FW��e��`��e�����MU0f�{����!SP3Wz����ʼ�E�C���e�/�D�U`n���M*<� 5n:��a-!���#D����V���7��n�>^�5��n7sl��7�C����xnU��e+������w���>�5�k����ƻT�2?��.�Yvc5VH`�0��䇺��ct 22o��)f��ѥe��6Ī%	*��sݗѝm�%2��1]h�y���ʙ�3�@��j�I���#�Kj#�`.�[�&�#1�����/7�L����F�I�GF8<ˮ�������9�)4����F��"��4JA�~hKn�0���^.��
8V<̷�(��o��)��8��zV faE�z��G�� �pI)\�D��}���2r21�[WǴ.ty^��q�z>P��M�{��5�.��i����e���<�냸:��Ĉ�L���C�H�)P�F�
Wu��P6�"�5p�rc�x=�%��te��������I�.rެ�"�B��ELx��Hd(�2�\���OuU��;Z! ˌh-CzVk��Z�EM��יsn:��w�����д��K�J\T��e/�O|�ck�$�0E�W��AM�j�崱��4�ց�@4��HY+�3���D�9�D�x�'������Kϊ��w��?83�R��\M�KZ��L_��)h���֓~�r�A6T���#d�D%,�V�Z׫�E�-�	��E���CY�z���O.�V2�pl-ck=��n��D6���x�~�v�l*� �(����~��-:h�f��GCѽ&�BM�����]���UFpF#�Mi��'��3DL���u�C6��ڢ581_�-Yj鯂���0��U�H5�l̚�	;�)��4�{�ǁ��6s}� �AF: ͡� �V�8�|�Ў]H�P���$2_�.v���fT��1��ª�����fy�6����:�f�8�^�g��������=U:��7Ph��5���e���m���\�mN�~�l��߾�5,�T+��y�1ÃckP�-T#������T�m�+���~#���4|/��2r�������6:�/\�M\�9 �x��@E���h�� e�Ǎ��p��'�	�Q=o�k�O��h�A��B�����#ۮ�МY޼^Z��G���E�|w�	gβf����	�6=QPj[#9�τ��'���<mB�6�͕Ր.A��p����Zܓ��h��l�o���f����NNB�`�]�G�[o��D�n/q҆M�] F8��&eᢒ�JwK�|����<cv��'mv�X�Jk
q"�=[��+��cEEI��ve��t8���h����ƾoU<��7��
і����aa���E��'�33U��/��-�g�f8��pFbe�t��/Ս��5���E��
vz9�Sl�:���m7fZ���$# �b&��)S�q������-`r	C���;r��,�^��KiY������=W�̳!+1"�@�:
�zex^}����XB��r�7���9���?&�c�b%/�m>k��~� W�	k��aU,�ٓ\�.ewj��!&$!�6�!)�l��������w(��Ƶ���O�Ir�{��y�3� �9�Jk��(K�O����S���ȋ^�P+�{�e�t��i��ȆB�F���J�;7�2�c���/ώ��_�lmZ�KKɩ�B��$��Du�~�QJ�еJ����S�q��I�i����K{_�5f~�L�D׋!�R��^�Z �ׅpR��������vM�sf}6�[�)+ec�h��4�afȮ�q�S%�<��
u%��\�{Ofb���g����U�l'NY4�Z�t��7	ȱ�(.�DCY�!�./!�N�s8PE������{��p����e�A`��.=��| ������u=��G]�`���B�'6�݂�����F��<��[	�ͷۄ�p�HR�����(ߺҊ��ڬ��I.}�>���tPy���o��i"����dw�=�
��Ӫ���7A$�HG{)v!���~,�wI��i��T�.��R):f;,�	� �.���X��s-������7D���hVl)��R}�%����9A�&�,�&������3�6�U�>h��}��i�_Y[��"C���t �j��OJa�^�2�O�/�O�/a2��~Ig>�D�l���g�T�K��-fo,&��|*(��E\^�35�n�G�m�k�W{}�뢌X� �z\Kǈdl���i����s*dEr�r�����I7_8���ݚ� ���)�)�R´!��:�h�0�In�
�|���iEA�a�Ȃ�����gd%~�7��[�@ o�:�Vh�z�g^�H��f13�.L��R,�4a������yn9:� ��@aT=��j����	�:�LTS��Z�?�3��U�p���&)����� �z���Bh�g��;b.�:�<���.�q\�ƥ�e�܄�y�M.����w����ݿ�_;�osjwY�����^>�6����T�l�M�i\���^eE����&B�{��`�n�͙�n�9�̻������ǆ��%&D��A��o�'�Yx��M�zAHT�cE��)�-�g�k��H��qƳ��r]��e�zނ���[N�nl��V7�8�V}j�i���~��}�.�|ys䞰<�`�"�����)��)��՟sa4u̼�a��^��Z!�;F� [(��c߼ʧ�ܷn!o�@f#�g��M*���-	{::b{͐��ѡ����Lv�3c>7<�s�P�����I�(4�qS����|�E�}1���I�LȐ�Xۓ�͏��R����{�4�!.C>S<��C`|/U��{���}qCmZS�-p���L*���X�7��T�i.{��~�i��TK�8�g�;y����W�_.��s��u�*��f���d?7ʫ�&�+�,�G�:��z5_\����p�G�W���򎡥<����$N��6�����k��qa��v���ȿ����ݑ���0��0�H\�?.H|c�Xv��A/p�,���
p�[�|+s�y�&^���"�1��&J,/�3�PQ����ð6/�
�C�a���,�.M"�ԟ�w�dGc��xq�9i����]\�����;QA�r�����:�η�f�h�u��o�&���-�#��uK ��T�\϶��N-J���_g�C�V������U��a��\��p��}�Mi�&!��~@4��\��. �;
*���z�3�rk��};��X��a#��lR�`�A�r�YX+}ݰ^;/#��TN#C�G�Y��ȁ �4+xBBa�j|K��ʁ`��
dO�!���ݫ�Gr	l�-��f���쏰���,(��ճ'�J�=``j0�f�U��"��������F�ӭ��J>��3�M��r��H�)���x���]�q4�1d��u�2q��1����g�.1Q��ȷ�D��m����ˮt�"٤e�d�g���DA5����k��0jl���'�hHڟ
}�Ǌ7:���,P?��Ѝ�ԮZ�T�k�V��l9-H����C��:j��X*�0bG�˗�\�c���d�H[mPel�(?J�y`I�Rå��K�7�l�r��1�1 ��-	N���x���N��3{�W)�p(�Ql�����
�޴�PS����HV�L�P#.l����rc���?����C��/�.����M뵭Ɏ�G c�)@gKv^�^z�t�h$k���צ�]���j>#�˞B]͜�|��C�q��Q).I[2�a���U͐�!O�<�'���W��i�7���
�e��� �C�6#����ƨn�J����x�u{mn���K�G=�oI>F��AD� W}�u�j{f��鹕�㯼	�,b��&���a�3w[dNw<��f�Y��g*���ʫm�W���R-��P:F�w\��p�2P������R�Q��Q�&M6��G;�M_3/aoP�gx�|h'�x}��Y�w5��1�O[�_�&)�.<� "%��7�gX,���mf{t�� OsEG�;���2��^�'/FP�T4�lT��V��۱�Q�]�q��I��g$1ݢ'�"����:B�=?T�H��-�"4��1<"md��^���{�*�����$�J"�B7��o�5׼��9U�؃K_�F��Ɯ�F��/�$;e79E�'��3�I�#�[�u@(�Y�$DGjt�f��6s� ��6��aH	I����P?D�0a����ӏv�1'�$:t&cp)���h��>�>r�n���?����v�t�����8�L$$��[!�����j�ћ4�n	�i�����y�[��4o�6c�d���O|�H���n��L��.奦��Ҿo*�덼)"�I?��̢�Ju�s�˪@b�Y�u$^��2��-��@d�4=0�*�ʀ(!�B۷�1�W�&��bb�X�V l�Y[(p��� ��Z��>V��w�2G� (+T���V;��dkw�9�xU����S�L�i&��-���R��'�a�T�c�V�#4aVR��!�oOߐzKɑ︗A��ë�\������ֽ��u�9,"�raa��Gt���߬l3����z�+a�U�����Go�䓟�q���7m�!��i݉0���.y�2���ج�K�q��S�y{Yò�w��'�2��f=�;C���W�M;�L����K'dh����3��@��^3*<��O0���h劋�p>^4�vC��|��o��\�%+LK \�#}��MUѐ_����P���٣9"�t���9�Gmn��b
�e���܃f��s&�TDM��nݔۉ-�p+v���1��9�u�t�*H������Ah6�J�X�!_#���o���bs��C=)m���-�}a<�ן�)��kM�J��w�j�`�呇B��lN<b��=v�\�S�� �y��7�~V+Oub{e��BR�s���o�ԔA "A�j��\�+w��=��H;�P�4 �F0�I�DApc^t\A�3�1^-*m4�J�aȨp��	T��pb�c {v�V�=Ow��E��3��=ݚZ�2��ܹ��v��6��
$��5�6Ĝ=Gs9*�X��/ݩ�*wq��������(��'2�Z8(�]��U9����*L�g:4�g��'��8�\/�)��Az���x88�)�ᢑ�`!mU	��6@��kaM�bl&vOvH��䮐G
R���$�q����v⚿L�b�qx�eN]h�\�Ol�pJ�BbT����>��������EZ�.ֱ��[��JG�� ̈˟}�S�<�P�~��9���^~��!@SU��2��~(;Fܦ�j;�b�)���zh�
��O"	R���`�j���h�$�X�`���&�fAF��
�
���'r���q�h+am�3�&Q��W��/VF���3�jFBR�vk������Ab2'�8���v��ن�Qk��g�r� ��X� '�M��4;+#�k� �Vm�z�I�fp�(6��&�	 ��պz'� j$+s�v ���c)������i�-y@O?��'��/'Λ.I'b��z��͋%��>a\D���R��A��>|v/1�Qw�P\y�8o���ЊX��P�zqo��t��1���_owYbo
p4����"W�xw_�R�(�F�m`4���Z��P�T��{W�n���u�#R�V��ye�v�@��S��a������瘤P�>f�[�]2�x�r�$�2FL�$���Y�Ƴ`?�<T��@>$���
Qš˧ơz��d�^m
b�ۙȻ.C���aO-/�@v� dGw!���ٻ�K����xw�BB��?՛<&ĺ2)d�?�iKڍ�Z���(�����D���(�v����ż�&4
H�D�<~Z�n��R�K��XO!�&P 58��n4�����x��%N)E4� �s����a����R�i�#r,�4�<��p�nP�H�y�� ���iY,	�{���
L�ܧ��P�*�b�[P��`Yٛ4o���0���x��T3d��a�g��� �mm!���)�"�|��c?�(�F����ZE�Y��ƾr6d���hp��:�J�-{yd�[�u�%TK."ݣ���;�=���/���S�h�k��VV��猦̯������{�m�ѱ����y%����S�Dv�ʙH�;;�xe��-�������yN�=ۓ���'m}��{��l�h(p�^ш�-T�[�wHY�N)D�Y�~�Ϩrv{+�'�f&����B��S�uVZkv�='�8��wW֩ ���W�my��RIS�P�w��.�U�\n0�@)^D�-1ЍnJ���C�Ì�С��/��0r�JաHMƁ���DM;�b��`db�ƨ��1�NwG�'�sX��H�u�K(h��؛<m	�8 �qD����<Zbv}~���3ߓ?�� J-��VfB�һ�T)(����d;�qh�����>���}ⶑz���*[F��2�?g��������)�=�(/	60(5��ר�?=�J�!���7�|�{ć�!-8�����^�1�Ċ��S�)�=0��q����e��V�CDF�K�?:�~�?�,��l���P��sx�:G�n`�H~��<*�2q��0w�avP໎i��y��"d��1F����/� ����6�����x���2C���(Q���If�{k�>wH}F���v5Fj��~�h����TDܕ�v'�S�1�J�*���CGC���I��y�aCޠ����n��� ��Ƽ�..=���?d� ���Ù���	��]}���f��0�D�7�t&�7/�;�d��(����W!��<�j��$*�l�#;�����U���B��΍�b��Ac�Ã+�>+�� �N�"t��1���Hl?	g�ݪZb%sA.�R�W-#(�r��a*J�k���!{ߌ�T����q�RћJ�e�`6����;t�C�~!���}l �W7B.��i�P��F(�ϝ�_q)KVo)*�#+(i�VA�_�<6P/k7��>|x �<�>���S�*&֞�(%����*�Q�R��#�cwK�jp�xZi�8�6����R���
ub;O�^��6�M��G�j<~�� .�@���i]��~vS�qo�ɶ��v:�u�s�*6W��v��U�� G!آ��C91� �J̮��#�A>���_�cz�3Ty�����#��T�!�m(�r?�*��4Z�?M���,������lQ,V599���T���?:��2I+�Yڄ��K3�>����.^lU���¥2rC�7��e9�QY��WToXE�{R�rƹK��Мɧ��}�ĿDg�����S*Bk�x�Q�V���o�g�qQY����q�׫�k�e*%J���@�"�%"|O�|Y)�Wf>@�U&=��t"O!-�o��|�[L������i*����Q�������ـw�/%�
�E)�[d/d~X*�ջ.M�b����Z^i�	��C �F9����a�V8 ��.��1xg]��snzđ��C/�U*�w���-!���Q��B�lAKf{�+i��'/ޘO�J��
��V�w[z7�䄘#+D��o	����|1��O�;7Jxuhpl����CMG��n�nC���H	2@�ǆ��u_e��'=_���d���6���F�5y�!�~ �~��J��bzYn�%L�,����9�G=�w�XR&���%U�n&X���S�7{j���x|��U�F�!���ra�����D�X��s�滖z5����v:��]t��G^M��+˚TqƊ�r'\� YI���I��7و�=���V�Н��9�q`,G.TH�JG�Y�)������Q	�uO�+Ѐ�W�0�[���-@���?�V�aԉqE�?��^��*Z�������%e$[<�{��`�n�1^�M_�����L�UI~Ҷ�+NM�*��k!�i�\�d��=vn��7����ؖ�Q,@�c�Ưǂu�zez}S&�q>/�l\��FŞ�,A�E�!]>]^����叭*����d>�ӟg���rn�خ��,4�]��$�P���^z��gom��68{��R՛�t�.*��1��{����Q#�)~�5_P�GɌ���#�F������]�c}@P�V�Ќ�2��(��ߜ���|{��3�o�bV��4�tqq�;'�;��0"+�jj��������@m�׫E_|�?#� ,�+GB��m��Q�>�xf�U#������Q�x<S_%bi�RЪ�oC���yYDhڵ=�'���������J��[��G �0Ɗ�����,�>m���_�$"{�2y%a�M�z�������C�
`������2�ͣ���=uiv��1�������+pe�HF4;巳�����Eb�`p�$�o
���������I�gㆯ���U���;BAAQ��D�9�������`�����=�![#�H"S����MM�2߹Gde�k��4�6�\��V�o��*���т-��2NP�~�?���f�0jrG�-`}���Gm�ԎZdR,��(a�����Ҕ	Su ���r�pY�X�S=�x3y�4%�$�6�U�!7�S@k���IT7B��Hw�K;�8�Tɳ4���bc��L>�s����	^Y�h�j��?��6��"HƱ�z�F���+@���Q��\�K'
��(em��~���a�)����׌�3����V#���Q�Qh?�c�[*l	�����[��`��w2�? <xE�k:��-��9jv��dEg%?��}��"��K�o^5�Onz����n��C�X@"Qoe���lɣ�[K�.�sY4gVhP!>]1?P3ƅ�WTZPd:�"$+?���>hM�fHcMܖ@��B
�ޓ���x�P=�̑��{�'	j�9!Μ���(��3��
��o���J[G����k3ZaK_�Nƽ�UieS>��F5�TlI��?0���2θ��	�2��t������2#���wB�ӼXp��\��,��N-[�[���:i��A(��GC���¶FOb��_�t�lǏ
Sl]�v�Ӕ=.�O���x�~XM�1k�;B���$;���D���k
a\�)غV&���Ē�.t��a �d\��y�ԿDZ�1�^�d�%K��L�J`�H��S�5�N���rΗ6����j�|�a����tG�����Kۢ(�|��,.���JRB��e�z4���5Ә�s����Q�*	������IW�p�<�۵B���&A��M��Z���ô�Rx��ڜ�c�?��1�;)�PW�ڔ�p��ݽ����_�l��6�('1�鲭�ЦS�Vܵ�>R�*Y���خ!̓���7+�
9@+��&�߭�S�_��_��-���'`��[ŷ!���C{�kh@~���N�V3n5-�9YGc5ҳ��K�9�|$З�BW �Ư����������}�D�\��a}�4
s��r��R�z��R�0���aӏʋ�6�}�>�^la�d�p�W����C��=��v�L��6cu��8ڸ����MZ�.�C�A�Μ��[�/�#��a�Ǹ*��;�"&����&�x�*��Z;�4A�|M�7�s�O�
��q܋��k������@��$_Ms�ܪ"�r�����6����v��]e��`1�!�L�p~��{�
C���D�@���>]4Rz}�O��g�
{i"��A͇{��<e���L�.b�M�c�Ǻ�!�F1�7V���/�r�Cɒ|�4��7�	!bC���U-.`��C=�{.��X�W�B�`����#Ĥ���\��!���b=�y��\�,�\�d2��WAd��:z�M��ɢќW	.Ѓj�\�|U\0�������-[fG2w�t�c����m-�/m�����h�֏c=�_�r�M� 7���n���%�0�;$	
(������-�!�D�!0�K�5l�Ef�PP{�A?W���$6����2*�＀�s��p3hz�����7�ظ�v>������+�Uyߐ��&���L!�x��d�Ъ�Yr�V!ދ��9��쫨0J��P�� *$3ۅlu|+�Іv����,��"��*E�W �q�|�n��2�u40ٕ�un�ji�I�E�+Q��S��վ~������hߩ�����P�m��8�<�P�cMiڀ sUG�^�EO�lBM����J0_=c�v5�N^ꑶF��\	�ɶ+^��!l�����<�sr^�,��Gk5���n*@"׾�����]iope�݌�{!w�N��a��eߓ=�;ȣ�p@OϷpk#R����]���X��$j�"�O�� ՞2z\��TY�3w��%.i)�|�2p�j7�Rc��!m����`�mqU
v�H�ܣ���]	%?�aj�2uZ��{!�Fn�)��3�un$>Џq�
)��&�x|_&��.�PY����A�nf��0����>�
�*��C�����i�5�����6�\�Ȩ�C�H1˳�L⳵���bc�z�̪�G�#~��8�Ú�`H��	�٨k��@�۳]�P�k
�T�9�V�`�3��n�Wi^r��>��o���0�IY�`2��j��;NI{UN��XK�[�!'T�D� ���I,-./&�K�7���=���%�G�d"�k��/� s0�sZSFt� GsM1�0��/
oxA��x�'�"L�ߑ���.�]�k3��ˆwfȁ�-!w�����u�(i����I 0��d�����kX��T��+h7̫Z�P6Y��a���ΚX���Ag��'��N�@M�F"rR\���~P���[֠/B��vB-��i�8"����u:�_�O2�R���!=H=Nq�,�2��uT����/��#�����]�>]�K]K��eָ[ſ+|� �cN��&�����q�-�gk\�j�}���#�z�����,���<�o��^C���ZE=3=�G��Lώ�z���z�,<��ܙa����"��!Xn"&>����?�o��}s�ᭈl�X?QTG�&+-O��+?��w�@S#�1�N�{�r_ޝ���H�(owma	�����2���s�LO1C�E�>�$���`����}x|:C��]^~o����,ktu+��N=҉HM����L4d��a�/<fW�%I8^ˢ��mlM�ԧ��[N�q�!�C�\���2r�����].����I��~���\!ƭc��>1�p.�5��c��G�ҁ���|]��Y�EE�?�9ÑW�`�h���W�^%c&c^/#|1�'�l-/Pz���W�ۜuYh��^�dy����HWr���`ś�;�}��	����)�Rr�$���R�U��vK�}��+pME���(O�)��lB��%~�Dg�����&�.�[9d2_RZ:���M��c!��B0����it�)�4	s����B�@��$�����z�� ]z]@W������?@�:'�-S�IGzi�����D������D����jh�I�ZX�O��A~�":����snΔ���-���(�Dju�? W<S� �_/YuQ~)��T,��
���-" �3�G�i�v��?�C biV��Z�|�e�{�y���ba�~�F3�e�)�j����V�_������	�K3� \�����c��k���Z�5O��nJ�K���t�wR�6����+䔦��' �?�iɥNB�O�ͳZ��P���A\����0����E5�}�V�6T4���fs�
5F��
�q��_Ϟ��/��v��:���5�Ti0N�1�W�l��*�$+�����n9vtrAmX��3P�A#��o_HMa;)%O� �ae�>�o�҂�&�����u>�3��*�����Pae%�ݢ�2���ɱz��g����5�Q�#�Ey�;���:.<V�c�E<�]��FG���v�B����W~�	�[�E:��\�ij ����6�$={S�K�m�V%We̢����n��.���Yv�xJ5�����8�9�~�E��qB/���� �=oƁ�Û_�yU�.���~f�r*ɥ.�f��^^�rr��42֝(�1����x�c�:㎍U\��~��Y��-Y%4�&/�~֖�a�K
�P �K.x�i:O$�aS�%k��48$�8����"4���q�|Ix���z�+0�Yr��PҌ�Q�wzX���0������C^i�Է,�n�Jb��ɏ�?h�w�O.��n�D|�8+�;��N��<��@��%u�C��lx*�ћ&��~�A���2z���\�8�G��)B&3`�9"��Jv�LI,3��T�e9ۥª�������g[��.�,�ĵu�v4A󄍍����h�u���0ES��������O��pg�+�7�y����^��Ȯ��"�"��������F-���qqѤ��9	I�� ��]���U��m;AHepfc���
�`�eY�/&������R��ؼ�bnf�P��{��d�Ա�����t��7���pSؕ=a�'Q�f³?v��1K'ZdHB{B��	NF�V�oW?�<w��&������$&nM�h�����|#�vo&��B�E O�ш����>L���^�+W+��<�Ar�����Of^�#��{9��˕�u���:I�w����?Y��T��/�<&�,�G�#���&N�J&��E�Ӟء\��~����M���R���C<FP��	�B!�[����=�6PZ�x<��JnX:������&�~l�]y���!%��Awrq,F�q���>�bO��^c��vJ�/X��۷�E��0'�>�<��y���2:��$���\���K��/�g1�g/ҹ���ۡ�=ɺ̏�����l�+�������#� J���7��������(p����'A.�f��Y��� %�RZ�c�&����X����(���s�46�k�J�2R7�ү��|��z�9�N�R[ܵ���e���S���;v��Ǭk0�����nbX ��L��'�u�vӒ�t����fo�U������9�&��ؼ�x���8O��%H�N�n	��8�?�ui-4��%��ݬn^���E?���� W�&�éc�g{�p�v�"v�:N;WW �5��}M<U�A[��>i\�8*z�+w.~)�����q��-i�9
� �$M�Jp����j_s��8#����y���E٢�OV_���4:D��Tbɼ�=FIț�6�v�tU��}H.���7K�aC?v�g;|�`s��n���Kj��M�xSo`�\�g��M~��v򨸷GH�ښ?�|E��U�"K�A����^��*��������$���I��I����)}���L�_>Kܕ%1ݐ��Q����l�Vu$�>������[C�Lw"�GV�zX�1i6C��ȖM��a9dCp��a2Eu	��Û,�z�~Y�pzmD�C|�s���'g8k\�l$����F���砢^I���Ԃ��Eb�fW���&Y%�"<0�]��X[#c��Ip��O�����[\z�Σ�R���]`�<��tbf�L3�e���Lb��uhU�hк_�ꭘ�pc�DG�Ƌ�!�K4��I�6��Hʕ�}.�h�:����I�V�>l��a��<ΤET�2�c���V���߀��&���c$�:���=�A^g�1�w��FX�M��n� r�[o�UD�X��FXߕ�9b�>J/��XIZ�	�&��)���l����b��m���` !��������p�j�能�������?���:=[�ב�S�-�wܐ�!G�	�N��٪�!�ZF��:{y����D��8��}�\�o����Sqw�����}�qWj]���Y}��?Yz_�=6�q��WF���F�'s\�z��ʁ���W�� �/ѣQ�[���S����y��;$CR�Ȑ��C�A�Vl�Kں���uIb7얆��9�����)�nb�G���� ��^Ooa>zY����ţ1P��v��:h"nB�
ö�����=�`0��a���LB�t;�I�����������\~��%�"}����r�[�Rp�g�v����m�'����D*\������1~z���)�C[m��e�X��E�a�Pq�4��6�+
=B��c����N/}���K�6�q�ց��]OD�J�k� rJ�e�i����_,��f�0"6�J�F��Ǝ�;n�^6r�-�j�
�ZPQ;wc�[~����d~�/�Tz�v��1�>X⬮�G�JmV��@�O|�2�����j��?�?����Í'�I�������"��/ո�Δ�7'�]�\�v8B�5F��ǔ4c����������{���2�L�t���R��ml��ӵ��{~I�]�Yl.wl��*�/fұ�ND��1����Rbm|��`� 	L2B�#��`��{pw�pzY���ɿ���[����9���V�o_q�O�$�|S^��C1}�~ؕȋ�x��	J�P���|H�\�O:H����U�R�l�ڟ�q�S��9Z��X���gJ�Jk��	5���+7>�=|@�u)XR��j&Ws}O��)�)�i	���S��ZS�d�G�2M�!hB_����P�F�ɱD�>0���zbi��lF�'�˅^��$���RZ���pr��R�>B���t��GL���h=���:��H<%�����$�(�y�u�I4�~:u� �} 3[��9�C۫RD��%%��3Y����X��/Kwж��U�ֺ���N�bFf�tz�zG9c�+W��]�\�flȠ<�4�q��Xt���5D�p�s�ըO#��FIP��Z6$�q��|P�2B�䷈��x�e0��]�?���y��#Oc��X�c� ��u���
���Rm����]`�������zy[Ŭ�1��K�!���b��vޕ���PD$������ϸ�՛���(~�G��@h��R��*sNJ��M0s&�[���T<�l�h�%A���ۨ�,r"g_�;���ݥ��f���C�>��<ɯPЌ?��c�!�BzV��_!���7�G���.%��Պ�c�6�q&&�����xfej�,KQ.L �NΪav��l��K�B���}By>����F��	�����d0@1�C�M����Rh�~}�f?���g����Q�Z�
��5�gdx\e�d��4R9��I���gJ�����B>�I��� ��i�]c�Dw��?Ba���%�p�6���u�5	q��n`D-�ε���z����v��I5�C+@b��U�\�à�&���r?�@�[x�N�%�������؄�%�%:R^�g�/Fl�;un����#�,
 ��^���^��� �$V�x�g�B�:�J�CSC�Z͒٪as�����z���H���D�����F��.�Q�{������Tvw�򶅩L<�������,G�U��᳙@}j1��Lr���Yӡ-�c�o2#����$�� �wX����Hf�	�Z�LO��P�8%�|� �[��}�`��;5��f����;��_	w�zi����T@.L�1;�?]�XOF�߲Ǧ��eNV�!����H�m[[I����3rG͗j���H�=�c�=����k�WSYM����7O�o#;�xV��s+��~�hqbsr�;��G����d�tե�<<2{�2Dm�3�y�%M���,v���lzHCd��>p��yr~�b
�P4��w����vܲ����T=�!2V�����s�h��tr�Ƭ��3n|�3�~<�|i�2 ǉ��*)�:��7������}�k�#�eD���Bj���K��|��7j���|��K*�M&����ԑB��V?�������s#�v�I�=7%Q���?T7A���(�F�D���b����.�_�IP䣱��U�۪K3R��d3H�~�iH���_�~�_�"!��5�fׁU2̔-�̽ׇVd���հ�G8M�'-(�'M�?��`��5�i�H)�k齩�u/�xW��?�񘚔�4ӂJ#S'�C�c6X�CG#�۪�*�}�z����P���G'�Q`�jwY����ְ���}�����ص��b�w-��{��>0����d7#�#�l%i����46�F�:`W��[��p >{))�՝��K�x�K;���i�V}3v���$��D�>@_���I+$��t�f�c���;�N��g��s�Ǯ=�>Q!����i��x9�X{Qa?R�����k��oT�ٷ�2��]��t��8kB�6��s�}�7��?p�T�3�B�j�� ����I5o��&��2���>�W�x�A��[M�	��\��R�#��~��G�������	�F�^��ca�È�j%��\�qa�'?�n�Z=r��8ok� A0�ݰ�a�nj�]���U��J��s:ڹ�J/�Ԝ�z�� �nz&��`#�Zȿ<�VG��e�9��urC�ܖx��0��W�T���{�te}�}Mt�ӧ��g�f�7פbr,�r�:�,�C_y�L�[�m�׌	w��o�Ͼ�0k1��r���,�Y�Q��]�T��A�7䞬h���8J�%�K��)ޠN	�Si�	��H_��ȿb�c�\����\���~>�]P���%`�{����絽7���)�c1���Wd�UG⥵�M	�HƂ�"|<�g+=Y�_b�1�܌m}��E0�Î���N2mZ��{@��\�?��9�c7x�nr�i͑>=�a���Tw���U���F1+C�VF�B�AI�z�2��X�����.�U�3cd�  ��`�R���� �2�"�$�y��E",��?I��s�DIS���j�`ا��,��7%���L	�~�B�OrN^`\��a~RZMs�*�$�D��>��;{��ӝ)�?��g9V&���8�L-��ˏ����Q.]O�s=Q1��Ҋ\s��?F����
 dwl�3w���5���{�?��<��45=��)^^0�Chb�)���q�^g�H��p�l0�5rpu��E���0�!W�Թ-f�W��(��g���� ��n�9�U���7�y��w%�t�S��FP��*A�X��R��@���sC�V�������{�a�i��w�����Q;`����B;�,B�j��Tx���'x������"�{=�!����,�|��kq�ڵ�
�\��)b�'%�Hc�
qpL�9X���UW3����,�T6Q��K�i�a�A��\���rP��
���y�ؚ{ȡ��v_���M�����8�#Ꝍ�d����7k�j�`����H��Am�v��T@��C����?$�у_�,���:�u|�BL�$�[�j� �����7s'VJ5�3b2��zo��,�f�`;��q��$���Y��h�`_��P��<����+T�N�e���u��_��P���MoߍN%L������2�&�SWR<v��FLS8/��5��	�z��6	���=Vq��z�?}֓�2BE뼒ܷa���,��z��a%������呒��
�[�a������854v3��ٮ�k���*��&Stv!$����}�n�;"���S!u������+͔n�gk�z1TSƴ�P�Qý}��,�8�F(��ro���ĸ��
�X��ѷ��C���v)2��]�������u���Ύ@�d�NHljσ:
5Lǵ7/X|�5eu���bt	����-]�"�ҕ�)��'�4��ڣ���۟;���vx��*�"��$�ލ�~�Z�T|�>}u7���T����S|��r�1Ih����3�m˝����JV�<$����%S�7�w�[%����%��PQ����C5\kB詢h(�H�
�*H����#}��B!��Y�`�$�R�-��o��[˱�%��=�r��^��ZgpLҶ���0��M�W���T�t�����B���R�*y!j�y[ϊE^y�4`{��@ţ��/u����S\�Qg���&��.+��r�*��s�L��3BrYC#���NX�o���o�"��u;��f��UH�ʽ׺�Y��p`�O���=���FG��O&�`����NQ�P�$w�q%��:Y�eH_v�oɵ�6��&���Ÿ�	�%���ZMHV�%��@c���l-��������??�u��ܔ� ��d{�BM�����a!ݥT�#gD�!�=���5��h�@�[F1��RǮ��	�X�]l���k��cO����26��~Ω&���Q��Y�����#�y�d\gW�w���?t[����&ڸ��I�ET|�?�@�͖����m�TP9`¸��c�Ю���Z��,�c�Z�yS!B��hKT{?E���ꄗ�0	��3�G�p�}�`��C�k�1��\@��uSmz[n�cl
&E�N4ݏ1Z��Y_IrgGm�55��y�w�q�#�oc�Z�"�_��S+�aS�^b>��m�X����!Zq,R�MgVC &�
�Ɨc�0fS�u��>���1�ml�m����/LО#��|���$������/� 6��\���1ְS���0J�уz�PW%��0�A��d��*��g�?N�#A8 !(��Hm#�>�.�;�ӌ��:c�� �l^�M6�4�=�X��ǒ�#įI��u��X��q�}�c�Z��k,��͇9Z�YV�%��<�P�&W�խd50����/O]������F*���7%%U��g��\��Yc� �\~�>!�s�7x��c�,��jH��sPg�Fik���X�������uk�!k����l��N�yL�,�n��? ����|qҪ��x��bW�PIMy�J+�6�	�z"�ڗ�Mh/�=:�3�W�~���	+v|�A���m���O��;/�eْ�UU��ɷ01�$��%����:�)(ɢGI��n'.I�D�}�g��ʆ�G�s-O@s���0��F�jLe�u,��#���|U�B��SL>�h���Iq�0�4GyT�������۶&��B�ɍ�"�lF1�z�NOs}_^�XDB�̅<�Vd	��"���@�!}a��z\E\�ҵs�_Wa�V�u��):~���h5�cE@���ַ�B��ʲ��z_�_F.fa�2epJъ��Юؤ���{$�E�M�YQ�~d�����p`4w�Iǒn�x7VP�`� F��C+m1��B�WQ�����e�F�/����S\-�@_�+�K!8Ǎ�=zҐb�XK�h}~�7�)m[�=TU7����)@�Ȳ<�ؠ���{�v^��ϭ�?����re�܊�ػ�?�VbI����v\BMU�����81)��}YCWFӔh�!�3]�`�t�wJ�~U�_�ٍ��;z��_)�������~�w|�՜�lZ���s<��iA)}�fUDd��#��;�����g��>
��{����'5گ?�8)p�=o�Ky]��|6��L}J!#�neTi�܎֘���J7��B2'h���*Σ���g��6՚����[��%��C;�� �(���f�c����/���b
v�Na]fv�	�cB�B�j�0����[��o%A�M�-ɰ`GtXm�������Z(@ etJ�$�eǟu��K��j/]V݈�N���;�MqZ�y�թ�*y��S�%֠�8��ؽPjv�"K3�Uck�b�陋�����1�;�UV�<�ع�¼���H>�����yߩ������Ȋf�S�����|�Pr˦��bʀ�UYo�Xď���N��W��w9�?x�M�ty<���vE�� mݦR���z��u�Jt��m!�S�0�yXL�2��s+UIa:�ǘ��S����0��`�&r�9(�r!��#�l+�ƿL�?��$�t˰�I��YB��}6������W�K�N~�C��{+y��j��n�N��������
w=몏s-F� C���26�Uh�� �)k��A�` ���<qp	�=��>ѐR|�݂zЃ��5m��m}ޯm��X0l$e}��h[�<H{��ݰ��,H��s�$����>t�()������ˣCn|����lw_K�7���|��;K��1�,Պǽ���</	��0����D�
��TxUIHQ�SbKf�~�N=��^e��y�iJ���b�$D����C�ʚ��Kxq�:�渄�����b۽	q�3��e�KYZ�$��2�M�/oP����C��Y3�gHʹm�U$ƛcC.z�s	&���f�4�ɣ5B��]�t��8U���}�k�Ã�8]���r0��]J�_�hX�6o8̮t�i<@�\�oNV>�e~��f!�ﺭʁHV��?�cj�b,szc�/A�Q�.Ȟu�e��GC�&T����^Wɏ
��`r���̺����r��h�E�r!QGz_�g�ZF���uO�4 �Cz�E���r_SS�Gs�q0��9Ӫ����-
4(����?˳�F�rPX��eɢ��k��{K9�
�F��s*@9u��f>����f���'��A-{��>D/$�؍��98`�xwPQ<2�Ҟ��{�����7Nst�]��Xg�"�	!�d�`�����49�!�.��oqb���+x3��7��������M�~�5�}1dm)�'��6yjAۘE'[ڜY/qq�m����V������]٩v�1|f����#��˗����=t(��;~�80l�*�QF��#/����7*�Æc��L�m��~m�̸�	�����Ԙ����N\���?2�
Wǖu�եÛu�j��\m{D�͠�V+�0�f���:ND�F��cI��T٠�G��'�
����N{�q[D)&B����^eO��hHD`mpU�5��zG.����F��y#!q1�B����h���D-T��9�D����8�ݒ�.;#.���z0�;�#	�`1��'�E�G��K�®ښ�%���T�ˠr<�'cgISC����TL�zP������i�B��Q"��ݠ�$�Z� �/��c�Ъ���Օ�`��S�)��M�$��S��Θw����_o<	��h����	ln'm�f�Z5;���s���T�z(F},Q�g9D�'.�Fc$@:^dun3�����9����Aj1A��QQ�͘p�۫���� �/�G]�����A^2T�a����(�(��=��h|ex4�Pч��Vi�˃ܴKR�7�B��"wj训����2�t�M6�?��座���Z�n�}�G�{�;6a�a�a�s�&��Й]�r�{��Rc/�W�r�R�d�?��L><�7CuܑîD`����an��#����C�N]�����E��!J�(���&7t(�8�1T"��Ma�bb�H���:��~Ȕ��N֝���j�ߺ/[b'N���t?�����8鑩��qC���;�f4��J��w����A6�/y�U�ׁ��uBJE��=�gl�	�^���qJ����\�g ;%<e��x��Z"'�V	�;ang��)wE7�-&���\e�C��|�?�ɟS䥿�.���-�'�HP�C@N�5���Û����Kk�n�$��m��B�V�12� �(l^<�L ^�{=�Rs�X8�wn07j��X�HS �7c�$ֱп��Aak���{(��QI!U2�ϣ@�O)q� IY��*��z/�k%Öf�^����C�1؂��M��E��)CǣЪ"��^L�
�_�=��5w@C9Y�ZU�%�Y�W&4<�.u��]���㩏�䐵�Xy��b����,<8���G����]XR�>���[z�ĕ��9����$~g��Ҕ�G��h'�Iy;x,XǪ(o��b�)��3�&��Y�B�mar%&����s�p��^h�w���qJ���"�%�w��E�|P��3��ɕ�ٲ�;[;7��PC�-��g����LB�J&y�E�b�������Ӊ�]7�Eƒ��(q�6�#rw6�5,���h��@6��J�v-�`�m^����}PR��gP��"��5r��U2HJ�gôqK�S��/|b\�D\2><1��^Ƙ�?!U�zr�S��&2��L��%����{�W��ρ��#�Z;$�T�c��p��GϙeK4�\Zw8������FBg��S�%�%�v�W����o�?�T�̅�}+�W��]w��i�:U3b��!p�ÛG��6�Og�j�X_lLK�n�����w��]�vtz-��X�Ēs}����7���������m��ݖ-�C�RU����)��PI��eF�<�^�*�&�����!�>�����,� ��<���<���ȿ�k��E�q��u�ZR@h�d��ڴ��qy�,�2�ד��"�݃��T`�J�XVǕ��I�mT�됮����y�8 ���| ~�GKX�W�)f�a��{��$+��vH����B0��)�M��ho|��|f�`�%�6�6;�����kߠ@�%M��y�Q�/��(���?4
���D��)y@�9���I��7oѭAڊ�o��`���M�}�o�=O$����"U���&�����5�?A�����c���(���d�*����iR�Y&+�T���^j ���X�!�R�ˈxϟ�$)�l�Q�}j�VV���
!��҂�e����n��|z�$~�E�[A���䟯HSڱ�=���k)�O�������<I�����݌��_��� !"	��ߋ�Ģ��!V�^�I}J��-كx�V��ɡ���^�R�Y��