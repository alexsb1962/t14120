��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[����%��B�P�O� ʁtA�B(f,�yk�0�l��ؙ��'�|�я��vsZw�%���9wU �����9��v!;>i�������,��PY�C�j��\�w� �
_��]w{����ӻ����B>;�Ϡl[�޽�<Bu��F�6��[�E`蒱����!/F�r�\�6:��9�+'�t�x��4)D^v?N��	�yL�����B�A�f{��HC�12��+�.�S����l�>���uT6,�6F���b�YB��h0W����]��7;�2
�{R�@<l�1MAC%����m�҃�Sv�v��,��}>Z���Ay#��Ȧy���J�E��C6w�I+�y6�U8�,�f'y6z;�/���0�Ht~;@����!���<�A���M��׌�zp�4�$�c)�H8�tɻ�T�1�Pli!w;EF'�v�曯�Z���޵��0_�4
h[��N7�O�x��캧rE[�i��טu�N��Ĵ��P����?&1!�($T�#���[e)�����kl��[C~��0���+�ET�m�3�Rg�x1I���NV�ȥ>t �sz�ŗ7�P>i��J�	�V>�%m7K�|��8&���.����I�m"H�s_B�ύ����W�	4��u	6��!	�ƶ�A��7Y�]�����n�3������3�m�d�.�FρA�p�#���9J��.������]%���
u���6gފWw��E�4/;�'�%_&e��m���A���mL`8�O����n!H���y�5\�pA�8O59#��
����� ��e�fs�E�^��
�$Ǘ R� �8�4��b�8���H�����P��F*����I�yD3���@0��ӌ�ߛ�Pk�Kb��z5N̦6�=�`�&7ٹ%O5����czc������vt��٤���;��X�]�ZL�FNGо8H����?��;�D=��r�;�D��"���v�=����!���c���ʏ̆��2j-����e�FaU��B�mح�5y�q36���q�4=�M��)\�r�m�T�qh�*�� ����CƵ"q��U=Yقb�y�K���J����Iy�b޽��h�H7������[��Q��s_ .�ڃ�rX���G��	�f�Z0���j�?��U�JT�"���UF��Z�+a�_���0�^- �٣��#1݈=@̏��w���0��F35'l�\�]	��GV�8��wPS�w��=[k�'6ITFX��
�}��t3}��+
V."�7噣A�HLplq�-��Z<�R�Z��5剿#�?��cZY��ыOj�S1��G�yKSt�^��z��d~��É�s�\��DP9�]���[����b�ǂ���3�/#�o[;H�-�
Ya� ��~șp�"�R�z>�J�'k���\��C���G�5{C��z�<�\FVXt���qU��=�Xdˀ�i�C&�q�뺋��� �y��� �����cj�ǈ�ܸ��WAԇ�|���O�x&w�Z��!.]ooY+4�nZ|M77���G�뜆A����)ϛ	�@D����ϼ��5R�iRϊ�Igj(kZ+r��v}?Iu��4�7�Y��X�E*!�l--$�坄���]J�8�b�_�p��^����;o��M˟���}"��=֘`7��6d�]}��fl�0�:��/�NHUQF �H �k�\��UܥR��AZ)�,�4/����c3��1ҊL�ҏl��=?>Y:.f�ʆSHx��<��Rp<��Am����=[h�fm[�3 ��M|���m�OG��-R��
�L5�m��R�ji4$H�?��-�����ZFt@@x�Гg8�A7(�!6󝾟�!�f�k�Y=+}u)
op�M��w��%8%,Ҍ�~'=`�c�D˲p`�yѯi=Á9s��^���K�Կx]�Nb�s�Rm;��uM*ä�don�����h�8vK6'Tf�]ʦ�PS��5
m�c��*q�|ڪ@Ã����n�� ���C�����TfeÝl�d<���
Nx�9L,�7O}��9ʋt5u��O�L
yvg��䔫W�~�z�ie`Y�Vms��9�G'}oK���x�:4�|������AM>�4بQ����wh�~��K���&�n���K~%�q{[A�2\�b�Q��ܝn2+�f������4���m��9^2��������A�{j}��rRf\����+ �G$6�:d5}z�p��
U�@��hp{@B6�拹���W6�E+K��{;��>��.}k��J��L�8����5|��`pz,��d�+��z]3�����PuUq��&!�Ls������������:��!�/Y�7�a{2u=�2Q���㑿j 1#��p)��9]]Y��F&<�mQq4ӵ�^��S�^m�5���_(F��;��Bޯů����\V���OaIk"��h����;��zy�qء�2��;(/�"<0�諵�8�:<r[QB��|�TϹ�����sz��<���/� ���ir�B#����_�RyEŢ騙����9��`{�\���O� `l���ޛq��vE����Ǐ�#�%��}�Ki>�g���u0�^.�I�W�<ή>����~,Ck�yaA>MIϲeT:�n��uӿk,SP�8�k"��Is��f+Z�gUbb/��-�m�t73rKf�o�X�2RU���7KjC�0�\� Du��? Z�и.�΍��ld���-A}�ܧ&!���w��Ԕ�x|yk��8x�D���R�~�U��a6q=�1�	/T��G�����5� ��g)ʣR��'J��y/�A&7yH;�BY5�ؠ�����4�\��t���]L�Z�i��ɣ�^�ig�A�̬&7i��&���(/����|�y������^G�"�"�B���m`�֞��<�h���e�����Cer�F,��V�l��@_�6�H� ����#���5o:9l�W�A�����>a鉎����9pS���jw+-m����I~:՞�Z��N��8��Ȭ�ռ�fM��q!���*��
3(3�����p��Uv������24�S�_~*��GN�>��;��'T�ѱ��Q���s����qoW�f< �e�Ժ�A��,�ntH@]�W:7�Γ�ܜ�����ct��C-�A>6�_�\Ǿ/RM�X��'��@�0�uDk�o��l':�x��k^�+�π��4z��hqQjc@��CIJT) k��wӔ���fr�I�Zߕvm��&�y�Gg�
2���
����\����W��$]�3=��Q>�=��@��]ԗ7�����Yv�����k�i�N&;�=��}�0h�Ϭ��])�^���j0�&;�֊nJ���^d5}Nb����_�z�l�g���jPϳ��n��v:M�\I�f�8����-{�iW��|�4��q5����I/�#N��<,�ģ�i�ȃ�����{H8@ͧ�g�㞯v�B�����F욟+C����	T��>t����|�։�贕�c�J�?��\��G��8N��0������{#A�/��ˉxQ�,!�l�4��Ymu�G�ǁ���$-�w �B��9V" VQ*.�o5(@�eV4��2��WK�o~�,������֏��x�����^w,����V�!7	�WԬ�����P}����@�@$�;uK��_u� c��
.��\�f��dc�&�vt�#���z�\�7�����?��w1��C'K������E��J`-�Z���������׃<9܀�}7���uB"ʭ\� ����m|ZR������d�9���x+�G��vEP��DbC��ɧ���G~!m��Ga�&���ZƏ��>�]h`.2��|��3�Yx�]�[�E�fĤ�g�=�C1Q>���"��݄~�A�VTX�F��GRB�U��Y W���.#V�Rƽ� ԓ��0�0B9g��;7fd`F�� ��ʰH��|E��h��
�	������ݴ��]��A"M���!Su^Y�?�{k06d%��_̤�](������������m�a$����C!�8�����1��Mvug/�"%�Z�'�{�#��Wh(LW�.d��
9�Tz�8�E�.6F���|gI<�����?��[-����;G:O,4�M���ʂiˏ��K��X<�+#��Q�pV������lQ�%6I��江��P���{��]�`A�����8�ԋkO�a����JG3 t���� ۋ�h�qf7��]7�uH
���ἦ��
s��@.5 �J��)2�_�V�Zg:����3Cli@���P�UlU9E���y��@�� $�l�&>�;G���<��� �%ʊ.���:�%X���s��k깟ţ���?���E5���<����
��$�e�*�����FZ��m��/�$�r��g{�h����&[Y�+BY$R}���i(�T����?J�� ��_�!�+Jw>��tM~B��O��A�&�����Q�s�*�=��'�B�`�K�"TRa-��έ�W��厈�'M�#[�$���y�u5�d5X�������X�xT�l;����R%C�<����vޕ�W�K�C&���[J�WzO�,�?%����f7�v�I{R�'ve����1�e���9�h��乴0�	^�ٳ�b�Ɯ����)"�����2�.g��^�Lo��$�L�U��K�� � �����eS$$C=>�6�g��M������g܅xNj��[����:�ۤ����Rઠ����fM	�� �G��5΀o�.V��I;��E�4�
��B�&T�K�W��(L�h/%Bx�X��Y�� ��_-)t�ÇZ�g��l݈��d��^���ݦo����������#�I��������ըPۮ�3k���Je�V齩��&�/|���- �=�>���l�w2S��3�--�>R!#���t꡴�:�@��bP�
�U[�E��q�`c���42��Y��ܱ�,�l2�m�/�9�Ă<�@sT��.5�D��z1���/�?�,�nvߗ9烬�7���ā�؎�ǁǻ�dW�k6�ޝI��4�NQ2��	�U�&ь�xOvVO�(�wHF񅋝�E�Y�I#mꌖ�1)!�� d��y}�������i;���S��~��>�
�ee��l"�Q�V��7��Z�h�]������|/j`�]N��T9=��B9���޵�.*�K�\,�A:(�sKh��mq�h%eY1�,��B���E�>X�;����/㟧�z���6���#��������tmj5�/��6����3s�7ߒ�Ծ<[7�&�fL����rW��~���'l��e[97���I{]iֹ��tn�OF�cWy�agy�v%ig��s�SPw��ۦH��0��J����Xϋ��U����Cv\�ŋ��4}�h�
�f C��\4�q8/�Y߆��ґml��O�ǐ"L%�%�!@��p��Bс`����������X���׶ѿ��)������	&Ԉ�W����"�(�_�+~�еo�΄��[~�ru�
�ce�j��ɚ6y��6(\���Nq������/@��驪!q�����º��u�(�
���k�����_`X|�9�k�8��(�d�b|��&�[OШ�%&'������]-p 9O�@A��_-΄m�(��g�Ϊ\�JY�>vV�;}�j`{�R�$�������!�e"m&Ηo�_p��T^i�&����çG�uc�vφ��a��ǈ>�u�$�f+�;v��B+;I��<���̿ݪ�fI;B�N(��e�޺-D��/�?��!gTk:�=Nk]�ɖ�(u��ֽ�Ƶ�)��8_��u�hȧ�^���&��B* ;���˒�"?]L�7�q�ו~�Á,������8xא�����o#��']q]Zn6��^=� 	u	tՆ_��K���	���֔}���D�4��a(�NѤ�Hl����S?�?������ے�~��ɽ��t ��Y���Z}���N���u� xX�FLHG��<��W0�R�f��!ѥ�tO�z��a�rݽ���������bY|���Kn�e��܂~��.[6��_<��j%%Ғ���Q;���e�!�s�M�5/?��O��ᡛ���d�m|g\I;V���ƞu�q6I�A���w�t�����׌?�X�Ecf7���~�d�B8����?K�]	Sfm�59����yn��4�/�4����D��Tf�D�뛰_3���5�I�F���D5�kܭ��N~Bѝ��!_�2���Ms�S��rM�[* ��E��@[��!`��gD��*�3�.��:�����}���49ɲ}TZ�\�?�гb�g���[���ieI�_A�w�T��� .�H^�Nў0T��K��������j��U��ި�Je��bP[�mh�L�3[�q��$w�������@NV �_9d��h�R���|�/EW}6�(�-����ױ����%�.��mbX������K�GqU�`��gu_��"p$�Y
����)����������"z��\L���ݥ�6���\IP����.ɜM��R"���A_#fqS���]?�yv���A��W�v�`S|�f��竍�_�p���,��$v6$	��8I:��ت�ɸɿB5v
.%x&+��@wb9��iک.ezQدߑ�ʁv�ko�g�:d����a�Dzie�Ȉ^�
۟Yʈ��e�\�nQM(�E�'8�� %�$JYw���ZX�Q��Rde��Y9�OE[�ua
�-]�Z^,�1le�k���٧����+���|%�D���3ݐ0;��]�lÔlJ�ӗ��V�Ӯ�h�[�����ͪ����O���j���-�m�[:�t�FN��	l&U�X{��jb&c�%׈��c�㭅!�;J��f+�^�,� �5�n+��"h�#��$�_Nەٮ^
�#���(����NR�Zʰ.�oVO��Fs�
GX�&|cQ��s���N����̹��0�,�i��#�a��y!h��+�%���1��:Y�@#�,�਴����n�$���5@�%7)gj(�Dd`����g0���|������a��Y�p��|�cbos�a;�mo�T'S��Lfzw=��zA(ݎ�ǲ�`릎������/,��ʙ;�X�swܳ���[��NP�m���4&ٍ�}��A���%���	b��u��r�bg䢨� b��5�0�����M�չW��\J�����:Iк��Q�����=�6���qŽI�NH�O��IB'�q���(�`׺�L�H���~���Ɏno�CU�M֝���
-ၮ�`���G��Z��I�o
��@7{�t\\��2���
xW��hYj����%+@�|v�%�I�v<��0h> #�3��B���aN�+�g�)����g��l�b�y��b����U�d * �����٫�xɁ����2	�zw�C�����T|"/%1��;�8..��Y�e�ٺ6��g��s�xh�L�]��
�@�)�a5@�Ӏ}���z���a-���Q�b��o�1�w���E�����]�FR���7�^Qn�2(������	g'�}Q���p�<5U���(�����9���Ő��P|����;^����x�yw�ի���y��Ug/�s%���8(ۆ�H�W8�H=�4����%�sYs�b�s�\v�d�0Vk����������ɜ̪��!�0�[yL�hm�mXZgBZi���A���k�k�>��U�Q� �+�p���]c�"���(P� �k�׻e� ���L­�u�Πnd�Qkx�2����J½�c,�!	��#39˻�I�(ګ�_L�<����x�;x0��N��>���N���N����.� �+k�ү��N�*�?K�l�xw�2Q�1�!���3
s'�΍$���sv���'֛��B9ٖ$�z�ֱ@����ƶ�2���FQ�5����"Z=�x;H���Q2Ȝ{dMLS+����ꊵ�ƺ�F�R�W�H5[7����f�+�I�:���qh8��xn�c16����EOЩ�g��� 0]ʂOy���)����� ������"6�pwI�cs������_�{�V$�����O�Ҧd�0+��H�\`�-�B�6�&�=D"Mv�I�&��n��J���Wi?b�����=�Ů��R�������4��^���i{1�<-L��e�I���V2|�zȰ9�I�ߓ2����޽�7Wn���g#�b�	����%�����yU�i� �G����U<���?��h�x�/�ȧ��C�d�^���ћZlp�7����X�Ew���4�J1��A�E�B��"�c���L;�%�0}"�f�,�-Gs��&�y'7;��#���<�EH�+*��s�l�c�_u��oAʦQ2�S��7,&�C�O��`��i�R�Z�?O_�t�J�\�T�`�uFWŒT�I�%�+L "�[�+�d�,F���_��~늎�P�&����\�"8BmO:������~���qO�����X����n�>=�H؊���^u� 	�:!��	VYP��j�y$Ϸ��<v?K��e��4��_���@����7\:�d)��{0J.��֘oZ�gn���/+�E5g�O]~�8������Q�D
�֎��cm�)����$��IM����uX��ɖ�dR�,;\��,ͨ?P�0ܙ�֜��T!3+���E����lLXA��*z�Q��1VN�~u���'�g��pu�zc=�b9��=�R������.���Zp���k�7*��8p��/�x����:����z�/��V�6��^w�K�AD�4�d�dlI(IWj�q��R�oC"7`$U��З�<�D�k��)�%Y�SZN�{mpJ�>���x�Ţ�>%��Q����/����2�]�I�9Y/�ך, ��'!Ӣ9�~�&�鿖�H��<��{��N�T[���͘��8��s���#�9ď
]��$�(���z�1���ƣJ�D5���]I��T��!A�:fBilé�u��/������&��V JrIxݵ{��i�j�|fhp�{~1�T!��*�SQ�:�4�ÈdE�a�Oy�I���0��6 �a��/�N��� f�.�.VC-Ȉ�`�T������ä́�Ay�KiORa�G#����)���L>q���.�4��Z��08zꯣg�@rWg`1�<�l�{!���'�)�ݟ+�H�Buq��.2�le+)Mu ��k<NيE �Q����B�z͈��충f� ��[>5�4.�.>���� ���񥺛PT����R������j-Y�����a�mU;kC��Bq%qߠ�?.zs	\#�#�
��b�����n�~�?tw�7��}�JL�&d%�V�����L���K*
�jc��>��@>)R._D9۠�R+N��O~0�޷@
���<���c�T�Ν���u禘��<���\���,b��(gk�b�0X���zļ �!�ae{RG�e�ώ���
Wj��\��MY��ЪJ����/҄��-��%zY{�����SBՕ�u�����'��ˣ��ڵ�U�;�B��9"�x��4�d>�n6���(gR�.d����z^s��Ap��(#�(
��W{�rߕW�P]����Zkٙ�!��p+#���0��
�"���&JFQ�ngf=t�MǠ"��Wu��<��ss7�Z������j0�` p���7�+�!Uܟ��t�D����8#n�-�b{t�dղ��e��O����jєzޖ��" ɧ�v&�,l"�L���/oz��v��_�{�H���\05���9+�K6�ax{Z�*֋�lM���'"8H��Ŋ� 󫒌c��s>hsзA!�f�f-1����O�'*$��N ������ۦ ��[�3���=���$�i��R�/��O���V{���4�~Y�]�Fv��C�raj"�o���W��°�~�U�
�Dj���Ԫ��n�N�/����z����}���M�� Mw�t���9����Ll�wm�}����h����I��W" i;�Z� �=�t�)!��~�� �v�nf1?n��W�����2�{C���O7���+	E���сH.Z��y�9���1����G� �D�,���VrK�]R&��H%#�N�-|���=�8�:";%g�:���L�v�xBe+�s�*��Ψ��S7qŔ��nڸ��_I$@�Ĉ���1l�����c����᷹��Ȟb�h%���a�/(�Ͷ�I���o�gp�$}�"��$|Ӽ�HF�AH���z�4��Ym���WZgW����	Q�fGGY<�������j�Y=vDΈ<��p�sD��
��r��.6��$��0�ǃ6G�D��8r꺓�նe�ߚQK��ڮa| d1�2�dʪ� ��_7cB���H�gu8"2�>t���U&�P�e�V:-�&K��Yf,��䫡��L"�Ah���讽�׻�@�a�eHE��&��{usy�pиc#�ҋ�eff������k��͈{<�?/3�x��E�R�ޯ��q␨#7�����d+CD@4�����X۟nT��A���[4'�Z0���{��`R����7��*r�t3L�0F�q���$;vf�Y}^ͻ�]|Y�Xi*�X����輭�ubO���hC�Ⱦ��`W�����/�Z����%P{��N;��{����Zٛ,��r{A��������oCWu��O-rY��Őy�g�����uϠ ��.o������H��:S�ih�ؕ����������h�{���К����v��Q��H�ot��e�v?�S��� ve!��"�������>�:(}��#���L��b��΋�V�����g�ǃ���@j�tȆ�J,p����0�z�͗�D�(�1���?=S�	�Uu�<iH�'�Nr��X[dB�ť��k�v.;�ë�0K���6`�(��K�1.˿����{�V�S�M�K��NX�����6��p���n���%�
�C��iφ7_߭\����L]�𛡍RJ:�wUG�-�W��^
^b�m(��L��L�2��=�$���Y2�A��P���4{�����fvҽ�:�U�ds֤�kƑhLX�K���L�zT���3��G�q������ƙ���"_��$��E�����^�]S�e��/�cj
&�p_��9�p��qS������,���$QU���D�-UQ�W�º��X),z^��%��YM��53x#7�&2u֙*O�V!k�W�&/''�2'�LMj~���E�02ޛ���X�+��Ճ+xs^��(\�� �nBN��$�a�i͈��I|
��|7���|x1�oʲ�1](���4�	��h2���o^C������w��]�E�r��"r�OϘ!�E�>�Ū�����(��v�x��R�M�#+���O?���Y��=�N�O�gC�1�#R6E}k�9C�Hg����@8@��5�.v�/0_���mo�:{|��wM�B���,�~��~�&RbXآZV*#�z��Ņ��h%_���zyi�x>�QJ8x��A}�nuA"���豿��k"�q�d��t$����(U�,;����@cv:[�F�3bټ��j�����4�	�d��V�+"�b@~w(V�,Ur����{[;-��+h}Z�j��5�LҊN�&R���V�#X��(m���)�U��:n�S+�Q�}]�J�t���G7\�FDN<�o>_,g��^��@��k#�]���m�#�c�i{:hx��u%�S��5�l�T��Й08;z�FҌ�(WqS�3gg�����<���{V�y��!p}�}ˉie<����ZoKy�
��__��,&�F��7�4͑2�C�cb$&E��]N�����V��K�����Vť�B~䗲�F�\�5�ɔ�(C��pr�R���w�$~�}6�J�o�q����dT�*Z�'����G�.��>�H�,l��~����{f��ݫ�[f^u�_E��b���l�B� (�R:Y���h���a ��Y�^G@*�L����!�'��G$�U�K,<�nت�S�����L��jA�:������F��V9q�����Y�U��Kl�~��E�G7P�
������5ޘkg)���9X��e$F�1�`��n!����P�Z_9K����tb�n��E� �t�=�X,מȎ�/$ٞ��1�AC xNZ���v��݄�b����D�dqQ��I�ˊ��\�V8Pp��:��t~���0YY�7w��*:�%`�U[������c��M�m[t�R���*�s21�2�����44	�a���?$�9Y	!d��	�h��fk-
���w�ȏʞM"yI����É���-#���iyQN�$p�1��������������5�N�
�V8�
<�H����#׷�5�4��j�Jn� �,�$i׌AN�a����jv��"�7H���򛱹��T�w��ȢsG�P�b�O��i�'�t&��@�qK^o�س�ul��LTЦ߼ebޭ��칃]B/{�L�#1o�_Pڇ���DxP?c���o�#����7U⇃���؎>BdrC\'s���K?X�����+�rP,�/�����i�pa��J)NYa�Ɣ�m�$8!YVYW�lL��U5�����T��D+_�4E��S�ؼ�k�����>GZ���Ꭺ����	>�����bs���C��}s����,�iԠ�)�B�Qf*��)WȮjLߤ���Z�N�|ǋ�k��6C}��x���~x���2.���6��^l���{>�[_�|+��@^�J�<��w�咈�<�J+�y�⌘�!�?x}#�,pyj�rxYv�Y�����jC�F�̩��?~X��,'�Z�a�lηf���5@#�����4[��XMD��=�X��I��<E�z�,S�/$��'���ȱ�}�:��bnW�H;�n*-�+��H����O`v���	��h�s���9lC��Xwgٲ'��Q���ۑ���]�Y���:��e��٠#-�(�p����1���L�wG������k�O�$��{(s��k��t��K�7���8���,��H�Q���2G�R:�a8_,�������y\��虓��$:��ڣ�%�/��uCa��� Kٝ��!}�ߔt���TC���+��*hb�2Ϳ�q�,o���fUS��������4P��K��i��i�S������:�&���k���0z�mVq ��@o��y9G����8�/�`�6�x7ތ��?ܳ�tL��Ȕp�!��Z	�D��U*�9�"�LI��:&P+�'�Z��Kݫ�hP	H�]:@��]�;'�X�f$�X�Nj�TN���hVi�;@� r�v�F{{�E�Yb-�o]��'9�]pAi��SkB����Ч�!d�N�H�2�g�pͦ�7ԙM����M"�?^�:����/� ��$�c�`��upfV]�����1^G�	���o������Gr�h�ik=�������_�
A�
0���� ^�����g<�pi�;g
qAx4Ź#���\��O��C��K3-A�5��n��od���Xυ7�qn��I�e�U�_�&�e�!��^n��H$�u�)Oc66����Q�y}]����].x1%���PG�y�ٕ���V$#O�p�l������Q�
���/�CTc,L�A����R��r�NӺ�ѡI�K� ��f6E����"�� ��U��j���M���q��"q�@�ĩy����L��p��)TAR`	"O�[籸�mT��D�ݩyENi���R>=T?1��D{v[��8���{�'N��;�S�q�<lL�q����0h�O8��x~��g>𒻽���������t����<�+�F��8�l4�Bq��2��Nȧ��� ���M�sZ��ɚ��Ѿ����dsB��<��T;��P��4�J�حI
q���<
<~VD��9�.�AC�n�{����h��7v�l�Xϻ�:-~�XQ
�ǁ�&̨�D7{�G4���T:���H�+)˿�U�;O7U�!�(z������J�4����v���
�пj����pi��S9/V�X��9�s����h��A���G$�8�kv���%ܨ�|@��p�3�C� F�<4Z��q{���%��g�{u�MI�<��zB�V���I +��R9�����,o�ī���Y*��Bō��eVm�ҹ/�}{x0��c���Τh�o>���������'�F`�[�
��Ǉ��iy�|b�%�;nЙ���#9�O�R�~y>��K���7jg�����U��HS���~N~�Ew��lH��bFq+�b&G4�%�u`��&9g���g%,�Ns���Y��<بMtH�Z^إ��� �u�L)iX�?��pch�Ք���P�c��e:C�or��>b�RJW(2��q��+���#��p�H��jٛث��5H�-&^oH���kGK�':��޿�L�Z����KT&�ֺ��˺q�5p��@Z�+���Y��s�a�����~���-<�?�O�1��
aG�t]����$�@k���m�p�YJ*�\:YۘZt��əټ�'�X��V>��Z�
��I�) ;T�eU]_����ٯ ��{�������^~�̠,H:`���졶@�����}�TU��U
�Ec�,ȭ�+���K��U����@H�%f�4��R��4~������D"3���`��>Dz1K�x���QU����)Z |:!�l!' Y}��#B�d�X���FT#7&�};��;��S�� �+`Qv�x�C�fALX���CP�O��F�]L�q�e+��J:��Y��`�k����=ώ�j^�zJ�S�e�[���/D<q a�����iБGr�N�u�}1�aNޜBs_y;.��=�X��t��-Ri�_H���ŋ
�s��{Ap� }�Y���A�`�xJ&��K��߭�)3�x�y�����Eˤ䙉L����N��#���t�}P[w��mԒ�G�=�+gϒ�eee�L[l�눞�yrr��ʎD͐�2|���O)�E��e:}V����:����k+<�y�XlY����?�A��X �m��F���`>�����D{����]4�w���'���w���|�ߖk�V"�R���*�k��ʝ����D`2y�:��2{h�f�cxQ��R�G�e�p�x_6��:�q_ن�J�����8�u^��A��*��Q�H��=����ԣ���wa���ڤ�_lx��V�65�*bP�Z������^�u�q-��`=�������@�۴��<X�D����󣏒�]F�d���ݞ�~��u\^{2E��g��][�V��ݱ��jP���I��8�g\����¦�;��3_BF飇���+�K+�h���E�����f�0��>�9h���
�l����n=�(�Gn����ح��-��T}`gD!HFX08v�Bߜ�H�3�m|�}����UϳӃ�l���^K�D�)���|��	����G����erb��W���B��:�%�k����Ǥ��NrI���KUд�3���pJ��WF��$�\��#|)|� ������١!~U��t��}��ҫn�~vylfÇ,)&������*�(����	�FV��0�p�b�՛��3��~V��=΋�P����>B��O���E!;����{��c8B��ysI��#&TVO��É�)ռ';�4�G��e���ԥh 3�����t]��^P�	�e!���D�������w/����p3���˺}�έ$��Aͺk�>����H����<�!5�98��;e��oxx�.Bc�n����..��C2�E��u���W�Kw�]���n��ٺ�R�v�g��7��q
�7�Qs�!�ziԷ�������D����nz!"��W|A�݇[0���E��?"X��t�y�������}0g�=/��������WpD�I	e�dK&���,f�-�#���V�4@(�MW�|�u>����1!^�}��Τ1eF���蝞��/�`tPy׆��F"��Ѐ�,BUv.�� �Gð �Լ���àc�ZI��أ-��?�S�#��+��"�-��-�F$l��Ӏ4芼�F�������l9u��てx�;gHgRߪ����$��C][?Bv���1؉rݕ]�S�Vy�t�2�u=�GfV,&�8�`��uZ��r@Sᩓ<Y8h��sWÍn���v*���kL(�2W�����2�'_z���d�T��m�jК���=�S�9��{u�\�����y����h���è�N漂�˞O�,�2�)��y��pG���P��c�u#���"fM[��~��?q�����1-�B�T^G���f�΂���4��.+BViĸ[��v.����̇W��9�e��W��{P;��KR�,�Y�����:����)��\��Y���=�`�(�o����F
�n+%�oCi�2��J�y�� �=9�~��c�zrQ��|�k�@`R%ܐ��5&��F�}+���a3�ϐ�ʖ]�JΒt	bcUd�C�)`�V$����@bK��-iT�4�0�JT���C�<M�,K�'ȏ�<V���!�~_���t�Ntyf]/�T\��N:�{�k��紫��wʻ;~�Cg�U�$����cD�k�zG��������1�|��u���X�*�����S����Q�Xߤ	wЕ����(�^F�R
��w5�a0_1�K~YK��ŕ|���A����e��x�TwX��g�l|E�(Z�x�F��#t9��:8����)fX���ũ �/�04���Q���3�!e;�|��(ո�joO��!���������?�H��^u)�(��(�K@7��O�TJ��K3��^�m-�}2�F���41`����c�G�1=x�����5��UrU�\ܯ!�~����p?���ʯ򖸃�q��d+Z�s�o�+��t)���ٖ�u[n�����:v�eW�pQzaE:b&6�����>����ب�{e����c��F��/��x�͠���LF����^G��.�-<�T�!�����s������ w�7N�k#_�X�9���9�%m�����8H�6/Rm���1Ki�L,��^1��/�=eI�:��{#5]}S���x-�b�{���h�,o���ϱMϥR��K�DgǢc�'M����Af�����{UN�6p2=Ô��5oo�A�V�1�g�j����6��Ҫ1��+0�7[7f�/N���T��zU���������Y�KbHA@W+"Օ1�S��ye���x��2F %���F)���T�:OM�Ұ.^ؖ^�*��CMa�x��`����TԆ�[J�vn��	�\[�#;��&��@�����9����D2��A��S��U�m�9R�m����
d���?�m�B_&��Z�YCܹ_�����8������km4;5��ae����'�v�������n�?^�Я�p����xH򗣯�	B r# ��ole�zJ�ͩ,la�C����im��k� ��2�>.^�����`YE	p���
�&Z�N�����|L�E>���̔<?E�}׿����F���Ii��q��Xt�h�r&t�7�K,l����M��~W*�c^�U�狓�C�l׹�Y�o����,is� �>X�������k�~R�[:��G�R�ɡ���6X���,&���bE��x.�����eY��^��X�gWiy������t���Gȸ[��_�X(`�O��V�۠�:�1�j���5b}l3�Kw�*��0�������5���AE�(��ЛC����A��'$�{��bf0|u(ss�׈����3�~3�����>�F���[{(w�lŉ|Xs֎;�wkc��.,W�����rƈ/@�i:�d�a3Ajo�p�\��'�~�ךVvy0A�
3���:�z=�p���1�bX��`�4�rO0(*�^�*-���rodA��d�ʭC�/�S�UU-��t �{���{�	�E�2�ᅢ����A�_6*���?�#B28$�����6;6�*>���$�G=Up�[�ө��p$s��6�P�N��-�٧g��xOe9�����O�����y���N�TH)���,>�i`�G[j�1l׾��֗�뺀�Ԏk� �c�.~e�ݰƏ�X��Tݸ���:˾t�gB�ω-��!t5�ݵ�z�$4��/lɋl�튠o����7ԯC�>5x��n����9�	���$��*�^�YIX%h�@k�ҝ�X�EM T�N��}��K9�rNO���}��8%�P�[���iῖ�4��y��G������ˣ�v��5�w^�<�i��F|������9�'�D�̗;���՜�~����Kc~�M9vC���(��X��O��v��v�|�u)�7�l�]?������^I��g����8�����st�9عV������.��Xg�i��ڱ3�҇�O2��r-�ؕ�M��᱆h��	��s�d�	n'�B��<��m^��O�S,�D?\R3�ox�����sS���u� ����R�bw##�5P�2y�v���axA����P��C�����P�!j�x	nra���M�l�uU���������|��G	��L�窹=�l�xZZ�!���Ɨ	o㺂!�4CW�m���2�T秫���~ n�~)�=I��:s���+�+� '�x�/��B'�5�Dzas��_(QA���2�{�p��t ������ �l.�2=��Ay������m��Ȟ8��{��R?��Á�Up�ڮ�n���kќ#�̈́F��u=�)R��"�8V�SE���~fX��r>�)ELH�s`C���8�}����d�PWoS��ҁ>���s�w'+l�ɀ�9B:��
)D�|(.�Ń���N̹�$�H�b�QW��H�>�Wc��V�s�) !��>���d,���%��N�q?���8̼ؼ���`��{�F���3	�$Цuڙ>5�^v���m��L���Ǳ�4So��L ��Z��)���� �����2*M�A2���;��lGg7��������,3ּƁ"s��&�\�ˮ�#� 
2���M��RC����Q��ugy���.�`ob����g�?�_�\�%ݹN����6�fة�]�j�oQm��MG������i�Ą[��*>ͤ��f��g���D��Ɋ�L�3�e�2x��:-���俄u��'�8�ʟ{g=w#��@:��W�nؼ���ǝ5m�~��=cGy����r�{��ږ���'����p�_T_w�����]�����ܜ�eܥʕ�׼gC���(mT��e��Je������1'Y �,9���� +F�h�*^���ylԨ���0Us��R|@�%"��L1�W���~n�ꖒF�dr���~�ۺ6�l�F��黅��w��c�"��/������ߡ��t�\"O�F3T�٦�n6䭯-6θJH[�<���(ےN�_(��Vk4�_���*���n��[0o�?��T�f�d83�ưaT�JP�ٶ=X+#�7Eޝ�h.�=�LN�w8Qv���UYo�9��ٹG���?hS%@.%��^��u}oM����϶��G�畦�y�xW�۞�SIpu�T.��7IaЅ)��A�&���H������%��)�ܻ��ړ�u��(7T9�V�Z9��-��m�{�L�U��Xπ{���F{!�r.Hy��\dc���jL��+A.��4�[([��S�0�h<EVQڢ�T�8�w��x��L���8E��2���U��Q�|��C�gc4�%.�����NƗ'�1/�r�L tck�V�=1���Ub�˧[�Ƣ����r��q��~������Nh��5l�9��8�HYF�Ȥ���% ��s
}�C�V��kl��Eܒ����2�l´��@��H��S8���c�/��"���a 2�����5���������&վ$��|i��>m����@]�Ɋ�m�\}X���y��s>�Ӛ��	*�s'�}k���J�����ŨN�z�/+x9��>�"�U�xi���n�J����}���ӉW"a�.�T��
p�K�-)�%��~�p �**5��Ǽ�8���H�s����&5#]��/��,����^L6���s�;���K���j�k<�UE���xO��8�
:$7��Ɩ�&҇*_��۷?��4ѽ��J�`˰"����X�ԅE�]h!wq)����7jC v'�I�WJwx�|P#�t��h���I�ɢ���Hn0Ci
��L�����+3�H|�X����W��S �z����#��I�^�S̠\�`��+.^�Pv�wVX]>�h8�����Ә��_��hi⍦��˂�ȕ�Te���<�
�
-z�����O�sĸ�ƍR�~K8]��ì	8�G���#tlnv}�S�M.�M"�-Cj�HZ�F���۝��,��{JDZ�����;�9c��Nd��I�%'��x�vYy�>K��Z+5E<��	��VQ���iZ�O����B$ކ4i�M��r�We1��o��.��"���������1,��A�|WЂ��L=���!�s�zW�S��TM@��>�����i���A�h<I?y�����[�����gtuPh��G{oye�}�J)_�EcX�R�@��.s�X��uB���fM���n�:��т�{4ޑ���� *67y1�TK�>*�h�fa^��H5��N)�܇2��E�BΤvї���'N_��h���c}���N���M4�C�-���T�Z��KCt��1�(*MöSO	^�*n쳗����=�al�[ ��r�4E��ݺ��p���l_[�$='�ح܆mݜ.��ޕs"R.Ű�W����CZ��tj[�|�Q&�SH��邰ѩ��\<}�^������8g��ׂ9�����+X�D@Wg�m'k%fl��99�'^�蔰�(w�������K>+~��È��S���~��7��h���v���ئ��:^����W� �Y�L��Q4���^��Vݮ�|��!y���ᴬȚ�2���m��ec� � ���0����;�ǫB��ګ@&�he�B����'A�E�<�]�Ǽ@C,��G���y�m+w*�Y�]�����g�[�vc�8��%�=������wxO�K\kB%��[=P �ZM��|͉j�����Ô�l��]����X��`	^S��ۿN�u���p�Z> �E~�CvԵ����Ciu�̕�퓌�K�Js����d�Πyw���8���8�Ox�%υ�3\-�˻�}��4�Ѓ�j����6�	��g@�=��G�b}�~��҉��{uYBm(r�<1�A/>*k�( �/CM�[=��o�6;��X�"�>0�r�Yֆ�u��:���X���b�:�w)��,7�¡K*S�tY����[���H��m�kj��٩��}j����WZH_��j�F����N��A��Xa�4����js�)$���T�nfI���1*����1����k+� 8=�FW��U�	���M�:��Q�:8��`��ܧK#@�ʔ�K�S�t�á��A���+�����p������S�6%�6�w�o3"^���+����� ������YO�$*���EA����o-_K��,'C��s̑)܊_�*�w�<��**ԠXZDz�[� �q�Lv�,�0W1�~��3�]^�1�����O[�y9[��ǫ�j�fO*�B���-������;��EJװ�j�����G�a1fY�����a!���O���ֽ�LG#����o��*�i�!w��62��_�se�����Ұ���鬔�-�Ah>q�X����X���6���bߧi��g;��W(���G�%�f�X�g*��������FU<����ţ�갈�!-�$[XpO-k\�>oYlT��PK�9%oO��9�i?��*�TY�OFDv6�����e<(��l0R�oK,��)������uc���|$������cu�
,&�Mx�3����WI�ċ�Ma��a����ֈz^`|�/5�gt�s��\ƹ~� ��;���,	6������1q�*Ϛؘ�����>5P�2 ��
_p�,u�Մ���Qz��.�qbm6RM�e`P���UZ�R�(�6�����,���Z��+�ZF}C�;H�Z���b�TI�!�E��}Y+r��ԛ�������w��\ڄ��}R���c�v�����e���62�as�J���=���e#n��K�q�b�=�}<��%4JV����ſW�b�h����f�W��~2�v}�'tk�
������I��1���e'�V�����_����@�	�D]���� �]��C���f���C�}���j�F�-i��W��"���^�@N��+g3聶�E/�Yh�.��4`���K�t�'��w�b�Y��ڀ���� �tH��q �D�f���w�~�A���6*�γ�°L|F�K������"K���xr�x%1$d��Ǎ��z3�}�L\�~����h�sr���� �i+c휯�#�L�qU�yo?\��R�o�a�Wnj`���eb7gһ��$Ý��
�GĪ�@ʐ|���~#U^�w��N��:�k)Ƒͽ;�к�JTvل��in!�1�\za�_nliެ��^����HQp��8���(8�f^��Q��)�XC���R=�<T�a
[��O0J��I��ɢ 8|�$�� P^R��J3[$�c�bs�ށ�O@����)�k���c�Ig��۞�q��-��.'����Fu���P��ۿ���9dC�����y�ן�1X���a
q<E�
GĄ�T���O�@���[���W��S�[w�|)��~)R֢�p���m\��a�H�Ǣ�xgi�u���f!�z�U5�FD�x�Y/)���r
;i}�g�j�#�h�T�r�Ƀo���9)G��J;�ۣ����'x��N�~Z���j�:�_�2�ה<��������K��)��xz��W<]��ɧ����8�(�Y�Q	`�m/�H�L��F
M<k��=P�:�E[_��x��S�S�B
�dE��R\`q��~�Z�"0BX&�4�����J���w�&��|�m���;�9UҮϜ��r��@�K3�i"��ش��m�Btq�Z{��Ks��f�9}��k������pإk�R�˷Wy����0�Ip�B2,���~:����D���G�����	�R! �o�2<F���"�!�	�e�e5I��;��S��r�����,�k:�
��X�Ӝ��d�$��<�۶��!�5�w���������_�t�8������v�3��sx���ZD>���� E��������8Y?���Gq�{� �c�V<!Ge�{���Y�YGr�!?+.�E��)AB����)$�1��$l^"��)�e��N�������W԰��+"���ilH�lo���iE�"N ;�:qN��Q�]pE�97���֜�0�r�:b����|��O�[�O���^�t�_�9�#���c�l(����WV�ך[����W�F���l*��Y���Ҡ�\��������4 ���%Cv����)����:nU�+�@I9�@'i=xǪ'��0��=�ف9��}�A�S���ߡ�Bث���S�Uz&�VCTC<��-�Q뉞��Ȗ���"�Ζ�M_�R��9�6� kKĻy��.�-��sh�fF�JE�rYߤ�s��'�/�4��=�,���X�f���01��{��UJD����eP)F;p��$�*`�I3�>.����Y{�D���HR娂���P�ã� ��'x�;�Z�¬M�=�gB�L��o3��NB���6Ϭ��[�&�U��id��cvI,���͕H�����6q�0�h�p�:t�c���%Zq_M�����o��pZ��1�	#$I���RK�;�V��p{9I����US=խb���b?=C��j��!]�2mѲ�mɷ��i�W�&#�>
�Y�f�.@�*�K���VT�Ȋ�����J]�:Z��Ï�B��r���HΟ�":G�����{�f��IfKW��R�Oy!�*�O'n���ZKd�����Ј���.7����_�b�E�	���A�<���t?2\��}NИ.�"��",+�l���Ӹ��8&E6�a/_��&;�����SD)y�r�?�������5����k���
�=L�1��	�e�d��'F�����Y�ާ��2��#�F\,w�Ҫm|���F����
�.��U(�r�zq�lM&���Ê�H�?��M�������b��H#���|��"tS���P��Q9$G�I��#��+o��`Z��N���K�n!Wp�|��0U��Hf:6۰�P��0!�
-�x��gV�A�U����6#��]�㮔��T2	�sk{�o$Ѿ��BFA��=Y���.̡����`W�E��R��`�'v��@��1�?w̱x3(��ew�� ޡ�l��\n�q��yR&���	&�J���9�n�#>�������8-?���t	l!=���7�&R2��U>��yv��p����"h��yI�g��,\	&�g+��rn��x����6_k��|���&�?1�hyW2ck��JE���6��AON	��Z�߸a�-��	�Z��IR������#_L���E'�F:ƶQ����Ì$ᘴ���#č��K~�,S��ƷȆU�����f�#�c�qʣ�[(�K��*�i~�.��rq02��F�8���һ�qH�� �{�-Q�3ﷀ04��]}~~�k$���J^������0�=��K�+<�6Xyf$�� �r���������5h�w�WhMd�v�}��T��흜\�m�)ا�D{j���1�
m!��X<��^*6���h���޴�7�N[�H��1���Ԓ���L��n��[�5G͑��O¼��Q�q�(=D�$�P��}-T>��'��ڹ��0�}{vA`�rBѡ&����Z���6��z�ش��[)c�!˩��xP_Z�k��3d�<�Im��3����UU��̔�%�&W�����ʀ\�QK&E�21m�����.V�(��B'�9MՒ�`�ڸ?��^q�.�1B�a�1±��'���������t�	ˢ�r싘Z���}O3wX�{�\�.��d���ٙ�}��N�lEѵ����̯=��R��R��u���[����Е���L_�zf~$
gҒ�M]�	]���u�#md1�i��P�O�*�ư'���Tk'p�.Oˣ��R��7l@��i-8�IR0�L�z,Z�Ӱ��<��Mw	k/���,I�&e�5��Q>݀��p<���;-n�"θ���p3�Q�}/X��3+�`��{��tn�Z��VEz"�SKB奵�U�L~9���߹��p��45A	�9�ox�h2�ΊO�B21k+�0\&Ly���nRB��.�XT��qt����\�#�շ����#s��㐄v�3
����nk=��/��o�a\�&#I�Yr!��X،�e��S��{C����W8�$VG�
yC�/�Q���r����VI�ϸr��40�5��wX�%)��iV�a�:�a�"].����Ϩ���Fԙ3&V��)y \	=i��g���b�b��)����s��[gT����b�1z#�����3j
�gA C��� �>y�U��m�ߕ8���l�_+v�U�N<m

����������b��G4Fsi[&�ږ-��@��+�_�b��\8�T�:�K7H��餸���D�o�z��y\f���Wтl{������CL��2�I��B�??uL���eYI���{F[{`�se|�E0�!�5/��g�ܱ���%ihsl��}�J��Kh�-�l���oQ���(x��x_�ۉʌrB�+���-���ى��!��r�b�5t������ၶ�G ���63*���/Yq���jFZv��`��z/�x0}�Ԯ�>J*ݝ�����r��R'�Lq�9������ANsW��g�{����;��=༥��bz�4!�IØ����*�7^)\k�#Uu��w�������$sS��n��39b<�H��?���" ���b��]AdtE���1�C����ۊ�	����][�l�Y�z&]�![����l����n`pm���g�[�7e�jp4�X&0� \Yh"�!��OWC$cqٰ[���5@�N�s�5�,�4��(��"�0W$����������}�M��.80<SC�׍ݧ�$X��.(mL��S�
u�N�cy
㡅���Y�_�D�ªe�n>}�?7�#k�h�=GB�~�4{�SΧj��A��yZ�5��)���02	Zu�+��h��w]�-vk�X�L�(%�9G%��KҐ�tx�/!�q��E��_�]��9�xӯFmC��ߦ$��1Dl<�L�ɬ�#mFr�9͚_������s0�حz<
���Ѥڐ1�Ѝ�Z��/�wv��??�����G��;�����PE���e<r�C�Y�i�
��'�&W�&I?aӮ�V��e��j1�Љt���,�q��W����9f#�Ю�\�S�o3��6�)"�v{����UZDЀZ�{h������}j�(R�{�ƿJ~�2c�U��Ij�9��rA�[{����2Y��b��V.�∘Uݓx��xx�����oe����7B�)��7=�u�w��-u<d�)Y���"oĤ7DF��-��Ej�դe�0>��8B��v�E{�����\�d9��!Q<��Pp_�$o�/\�9Aq#k�#S*hT=غ$��Ф*�����!���]�|9w9�h��9䋃�F��\��'�a���ub���f�å�xM 6���ؙ������MM�=�j'}KOfb~���oa~�_(,���r�������&Y������	ޠZN�Ei�j�d����'��v�[4�H���!@��6�z�ٮy`:BӀ�D\�wiQ.,�&���}�o�Mv3k�KN)�$eǌ�0�`~�/"�������V1ru6�G��b������~ӡ"�з�V	���x%�o������o��U�q<�
� ��38՞�/�G�fK�
��e8i<G�o����#}c�6����I_���̷�X�m`��G�Z��D��οZ�S������AE�?�n݁�I��}���V�X� ���&���?o!r�C�O�J��j_ �U�\�x$N���aY�� �Մ�f5��WUB�{`�-��Kg�Ж�<l/�A2vQ;ځE��<A>�<��TBgh�\s�>��f����F��_y���h�1�Uæ@�#��]5��2V��4`�$ѬYLw�}ip��Ჺ�Y�x�I)R,���	N�jk�p�=F�sI�y��m��e��8R^`w�in��0�y�X�a�}�bʺ&H2����^�����hi6��Z2�/-$��k��o2��_�6  "�YlC�@zc(��zQU<cX� ouA�}�ԣ~�R�8]���p���%�a{�G����#�7�u�0���(��e�֩�]�Y���+c�(�ծANȲ�!&��^Eh���]����Z��0�$��;b�d/Z�~o�~
dQ9v�1�D����`��y��Ϙ}ד�
��tG u��O�x�;��i'��>zb�:W��qLV,.U�-�;�0��a!�Agn-�6%I�}x�Ƌ�٦#���9f~���E}�J,ŋ� ���MC�1	@�.�T���)�W/��#+?��,խB� �.<����1YM3s��.�i�e@54�����"Z�����\@���@rP�%4�ޥ�������� K�a�G�>B\2��ݲ�����B��L�B�kkyD <<a	YxA�u�R�_�}{��L��lU0��!���悉"�iV��7H��C����q��d�������'�s��}N[f�t�dY�_`5'OE�$���54>O��Bi�z0�0�D���Y6�9_kTd��n=��&�����F�3)e�n�~�^�|̓����
<?O�C��x�?��9�c��YTY2JJ$Ǡ�R����E�Y�%y(�u�]��e	q��� +;L wo�LY�d�q�_�ޭ�W�i����:� L�V_7���ɊuOs5p���ʮ[i��?���7@�l�>�\R[��ky�������=�{�ө�	Fr�'�x��h����nq�J-F�Q͡����-���D�R��S�0J'�۞��cUr�CílM�$�3�����g����� ��l�׹���&
����yWZ�ʂ�����!��D�U�Lc6�n���oj�	c��tB��&�u��#�u�� �c����q��P�[�,Q���+�V�zY��N���%�$cr���_sEMz�\T��c��x8���Y?������"�)Y_[�wɅU�ڵ�^��ʤ� ������XWHi�U��2�d]�j����Ǣ�~��$��v������`�7� aAÔTo�Y����_��I�Q�ۢ��+�!�ב�4J�;S�~N��\�A�y|�)C��h��b�v�ǀ�%YNƷz����2���B3�L���[��K%|KPZ��8��霘��V�W���1ey ��F�L�F�2׶��{"4~c��J��?��Z��%]4G���&�����nq��ל��LĤ�&a�[���o1��W���eO���?��7��@
�]��.�&�7�B�O-��d]W%V��=!y�X6�b	���f�2�L&)P~��288Z2똓�@����+�wn7]�|"�NՏ]r�t;�r�Qw�?�:ϕ� ��GX����6�]
�LD�[1��|Y�5�oyuҭ�o��ej\|�B�0Hc��h1�~ Nb@���'�ya�o�Dj���p�L�Xi8�)�uC�3뚺'@��ȟp�Ky�f�7qѰ�p� Ά�)�뢌h�i���v2�n��)�sl�1��]˒��pm�V�,�Wb�� �8tOZ��p_ Z,U>�T���%�Y�_#lC0�p�f�
%I��/W�j�cb��-C9�~0y��������Џ����S�K�B﹣�ʢu���ho�8�<��+Г��&%� �rC�1��'ǆ.! �򥦇���g�!O|o���R��u��}		���=�;��#ϱ�uuI^�U�7�<���1z��ʤ�E϶��57�����d}�З� '͎�}����:Y먒�(�sC=�.�Q|��Uw3v'��si.R�qK�Ve�P�F��P�K�~�=�����֊鮤��/4����!�L]�c1�lU�`�Ȱ��(C�wv��=�?rU���h��qU�>8�%�wC��o	��vmf)�sg7���d>]8�')�O�7xف��΍��2���S���d�T��V�lYx�b���5���}���?��~�z"�g,�=���,'�dX�n��z�}ү�..7��e�UpykL�����G���.F�f���Q�n&*#�S��y��\8�5�c�zPE�l���Z�\&�"7���MԵ�(ē��m�p��zB�6�p�7w�fq)�S��`�QCZE��!�j�^TC0�́ ��̤��7��xd�J�]�aa�:2�g����^(�"�?��'��.��N�\y:�����'�X*���8/��ފ�f�5�	�d�C�@�vi�U����f�AeG �ԉBb���2���S�-��B�x���A�P��p�AY��e�:a����@<��<qJ�>5��>�%
��0���5���ʟ�|q]�(Ub�S��1�3��Mu�Џ���tL��*UL���(����t,�=Г�맖�mm��4����M4F*��Q�H/���V���9+jU`��] ��G����,�+�t9i4�C@�bN)�[��"��aÎ�T�Չ�T̨[j��jT3mj0>���᷆�<k�Ұ@v����M ]�br-����\8)�c�
��i2�ṙ�/�"TBU�(� ��۩6�����@L��h%6���79��#�Mn�2x�Sp\���#��
�g�l�^�	pM��8]�]~�۷��[&+0?� $����}�?U�gV�,������"� @0М�~�-��r��_��v�>�K�,fԢ�.�H8���ݎ2�Uח���Rљ4(�Ƣ�|OH{�����R�N�+0y��=݌-��0si������i�%��;a�g����@����Է�G9}��#9�n�V�֔+S��{�Շ{2kʭ�" L��!�����y�[_-��7�,0r��Gt�aN@I�+�e�U�66^V���W�43r�^Uq�S�ζ��T�#q��8@����p;�1a�L�E�'A�V�#�w�/7��W�G��T�C������%J�'G�4��_���ýV�)lb=�������U�-5^����M��so�|�j���*������Ϲ(�rtK C�AA�1ܢ�Hk��V9>��Q���a�{a������aW_��,�=�?l���Ҁ���r&G���Z�����$!��r�R{�,�@Ed�^���#�=��������8�Ŧ�r��DȚjn���:���6��_�Y���(䄥?^�{m��{�(�/2�'�Yӭ#�flv��oD��_��SvX��]Y`�o�s�C	NO�(&z�H�12�֣����晁Bn�e�P�	�r�5�G/�@��������PdP��;{�%���\�J�y���p��f�x:-��R�ZgF@�b��o�[8�S;]���"'����9��N�Y� ���}�Pu�]��\0�W�}��_T��*֛�0�"j�QE�|ӡ6�Y��y��W���%$�7���ѵ�fI�π���K�Z��P�3,�Tb�����סk9P�sm�tGڂ� �4iXĴݙg��J�/.i��Q����?H�lё]n2�P�$�e�am���$��}���7��*�k�S�x�k8�J�m����Ή�����鮕�*|&���5�5ܸL�����Q/	s틱�-թ�ap2���}r�P�[:�1$ы+��
hL+�y�$c_��3�@�%�Z��1L1����n7�1�l��"�~^��[$W9�S��`ޯ=<���OVs�(���EYMc.��L�3����Py���S:hB!ܿ�x�z��%
C�f[���$��G�-���xd#�M�$��5�=,��<���SYg`qg�u�;7��uĊ=�o�BU";V��imfb !VE�p�O��T�<D�[<4+j+�M4k��Fr�v�t�f�=��l�0��<X���/
cG*��,��-X�*��P��m@�-R�����#���\������^Յ4xU�hL��G��X�(�L7����b00��"/H8���1�P=�葉���
��J��=�g(�f+�j4t�s����,�Fa셰﷼yD�B%�E��4�YY#���YDs�����.ͺ��Z5(m��L&ApW*qn�h˧�Zw�S ��)3��>�9����b�y���\��4�8߃�����_\��;@
v5�+@0>C�)���7!��U����~qs,��:(���^$J%g�A�%ެ񲫁��ԸH-�>��+�k\c�\�)}>A����� .p��d�����4x��C��pr�$@njJj���g�Ce���?�0|�� ��V/5ePQ�4�tSI�4MR�U9�Kc\�<=��WӉ�0E��ғ���Ԥ���vu�SТ`�Ҧ�O��bAF��nvb9��sE�Z�ĝ��U�X�i��bqp��kN�{R�6�㎛��J���7��.�W3�h�1H#8Ì�S� %i��N�ţb�-�]\�ē�H��N�V]���� �ӧ��!�?1� ���<q�h� �G���� �)T�DIts��Uo?W� ڎeV��͐��nO�b�;��<�P].ۡ܃��s1M�ȱs�g�m��̉y=���}$`g1���T����0��(󂛽�^�Hɽ{)�W�_�1x&c��aӹ�B�5�G��7��^�W�GZ��[�'��J���\>��*=�H{�"F"��U��xum�5t�zp[H��3�Z:�א����{L�����V��o�W�	B_�o��Ć�*ZPG�޻4A�d����I���x:��I�U�΅Y�йuI��j�Kh�Q|x��2��|�(�8�4H)	'ٖ6)��V�Oӹ�ͭ�m��
�����V}J�uׯ��8������[��E��wL�q������C��*Ǖ�v�b�恉pO�����e���Ti�i����P����e�Av��곹�O.���E���l�1����E DZ��8�h�H�8TE%2����}M7�h���bW�'����p�oS"^��B��	|ŞQ�����"���2\L����l��{�ư��R��/1.����1�}'�>��7�E�}�"&�6�h�I�;��Kj�>�&'�z�g���!d%�U�R��A�ϵ�ZQ5ÿ�D�3ć)�?�Kڨ)X5$�%v�H�u	�ŀp�Cڴ�M�z���z�Y��ت�Mc#g�Fl[�����	�<��g�3dO`@���ȀPdWN���r�#����	ϯ3֜Q�ǔT�%;��y�ۏ����|��X����իv�(U��onZX�m3��_C1���d���-@
"qe������9ǒ]���hv>�;��a9u��P�O��:�K��[B�<�Ѝ���`?�8D�L�{�K��o	t������3=2�kB��y<!�8�&���Ǌ=���F�iq@mFV��,"o�D�ޅҮ�{�j��l����ubq�g�րA�8�p9W�4�?�@*�h��]�(J�=��+7Yݥ�W��^�ы �����57�� ��?~� c'x�j6 �1;XS������Ƈ� �4��� 6�3�-������`��L��n!�u����8�Pc�]��W��e�??r}��UJy�c(�j�?5�����<~b�K��*��V�$�ko/�P �-�|��8T��WQ���lV9�|�W����:l�4Zie��+��x���[�� �Gҷs�*y((꬇�g�����O�o�� Gţ�8�/#�A�ו��DY��u�`+��٤�����Ѿ���u���7�\왧��L%�B�m����b���f��H�G�1giN�b;��?���^���/`�,����R�}%ExnU�1^�9����3-���sE�?�p2������'xJ *X������֩��}����ݥÞ=��Ó7RA�3�N��!�%���`iÇ����O��Eot�t�BT烵�?E�&�;]L72Mvʵm��1H
��U�M��̂��F��>9�������^ti��5�!��_-b�����E��D��jN ���/�M����)'l1A�$���	�\F��H�b���4$1�#����e�����b���@���7���^2�F<�ҝ��/-Rŧ+nA��Z�����׹���'�DY@�sfP�����a����#`��,ߌ�q5��?��=q�,�X�UJ��A�p��{F6xW�ϽM/�|�� 
�A����Xز���z�8����9@�,�fϢ���SR�,��ú!j��G4�yg��SNy��51"68��'*�.�R��]W��r��-�%�2�gE�rLt��|��o��zIo�,g�<�os;�NLV;�N�iok��&�f
�̊$��Sf�JX����=�J�A�*[<�����,V����t���1p����oiIԤQ@{@6�)�:�8��9�&4�]��"�8�.a�>_N�28A����A�tI���{���0;2�co�` �����qXh���Ɇ��$�R
�iO�6�s�40B�h �kU�@*����A���<��2���ފW?���9�b��.��Ù��� �Mۡ�6'5�c�����Z�9�{9/1��q�m]�����1�)��pP&/��ӿ�����g�|�/峺��hi�oS��|�D�U�O� �bh�Ǽ�a�lS���Av���B����Ţ�� ����ڴ��r�J��5�j��㯲�)�?�nfkd�*┾_�e���kD�
��<�?��Cߢ���s� 6�l�f𥓞�W�2��%��_�������e3+�HTʩ;��&&sp<2"�BB��>��{.]C�\�Ĕ����߉xEC�֮2e�9+��C�D�����f��������Ws5���^��y�8�(�`A�_q�7#sy�~�C����r��e���p#߂]�7���w��Јv�ՔHkR��c�^Ѿ&d�Z(�'=��&�Ct~��D��؋�{z�Wj'��H��/�;(��,�ܪh��
AQM���,�"u�+dK���4=b텛���%.Mݒ��H�!r���?2蔳~�K�iJ���3���ȩ�5��
KJ�e�m���g#�+P?��@�ح;��|R?m#�;�hڣ�.�]���I�)�w��Eo )(����E.'��{�ΣU�C�x����m8۶���DLCT-~9=�|����Q<�&��f�2����;[h���܋ӄ����`�I{9�=���7y�8���<~��W'o��(��q晛�;x0d+晢vY�?��w^dlO�����2�����_�8�U�,��F[�U��9k�A俧� �TX���ђ��o^2�����r�H�Ǡ�+ �
]���"�	�A�M��#kF���%�؇i1�*ԭ�1?��)��N,����a��HH���ze�rtrp��}b��o�s������������B�8�V~@�(7SHӀhO9*�aZ�u�o)�^�$X>��L&�ŗ�w*����R�f"�1"�	 5�u����a���q�'A����6�4��V���S8cY���og�4��Eߺ�w	�C	�����N�R��&�|�����~�E���I�Q��q�D�lm�z�+J������fgDjL�-�;���ћ�:_�~��Bن��J5@�����/�^Mn�� VY*�I�Bko�=��=��7�u;M(U̝9�8��P���0�a?�D������Y�e��D,^)�7b�U��F��ʳ���/��$R��ŕ_Н�؆nވ�
1��w�w-.�1��I�$'&��d.�8��6H���r�_�V��Y@[b���i�g�':���G>u�;������1[Ⴅֻ>K��0s�4�`=A��	F�>x��`7$p��MVm� �W��5�΄���d/\��MB�����&�w0��	��Z��~�#��<ø������E�/���
0Ѕ�&H	���Th6�c4co��dNb�I%uN���PV��H�>@a�ebq	��H�!���ȏ�"�2CH�	E�x���liɅ�	խ���	�|AV/Ce��%J��h0-?�@�M�7!+�V�X�ۢ(_\��b�S}������Vff��z2�M�X�TەEl'g������`BG�(7��[:GE�oK�C�>�����b�Z���ڽlU0~L����q�Uc�v\���H��D%�qZ�����~?�JvR��kdpT�:Qv\��0|����2�a��3'��禋3�U��%{��'j���Y]I/5�޹{�l�p	�v��f׻~����V���|��ݏ}x�Ĳ�	F^��5g�[]��f�]��47
�!��h���g�+��¾Ū���Q�-���Er_"�ܟxD1���	�d'���ӊ������x�������
�7P~�g�6-�&�5M������c�r1U�<>�iC�^��ӓM["��K�~�bcG�r�ЗJ���I��CA��y5'Ƙ���Ug�����z!a�ߕ�!�4����T"^&L��Z��,�������? ߫覌��9�ʱ]dN�Va���#�t���	�ϡ��P@��!��T����>��$MT�%H�\���
��É�M�'���Og�hwo^�����>v����R�HMt��H�H�n-��o!�>���]��Z��!��-�����<�[�^]�-�ާ?s�s@�~$�����������"�rU9R.CQ;��QJ�������:���ߐ�4��m�jsوdv$b� g
�ȸS3ļ�.�S>�ݧ~٠�em��qs�܃Lp�^xv?umOpd_&R,��V"l�f�~�Ԑ="��k�>��1]#�$r��-���|�����u{t�\�ƞPŪ_>&�y��x_ߪ���20�m��N�\��#�m���[���{��+H��IZ��PW���xJqc�&N�#�iȎ��/�hi��n �ֺ��oMN�Տ���^�IA�{���%G;��(�q� ��J��1a'��,�����kj���|h�U��|*�12V&��W�U4ƍ�V�� ���$��XPn���Iv\?�V<� elwB)].��\��j���1�	\�P!�#����g�C�Ę1!q~�������Փ!��4�� �Ë��ݏu���ׄ��1�ѫH�`8e5g$'�~4	p�²��=�C�-�����{P�6C_��������l��BKU>�&�i��-}��I������c�`��k����Њm��B��㲧���o��s�o�37�icUun���PPD��G�|�- ���K��ym���P���S�����${@��;t@C������d�⢞Brh���-|�Uߦ/JتrJ]4v�-�d�S/<���JvJ��;#��N�v?�2�p e�l]r�I�j5!K�QaO�t#�v�x�ONU�\s(��E�RΪߐ��W����s�x�]i���f(:�LE|��ښ���y/y��������s/�����Ι�;&������^�1���ڤ�xW\�󙦻 ��eLH��iM���*d�i��W��C9w~�PUoW�q�?�zꭀ#���ʾ��z��ڙD��!`�og�4�Ved�յЄ�*<9� :,�j�}�����p��7��S. �A֯���,G��Q*<��ZU_ѱ~q�Z�)x�y������ϗf�W��w�l�4恗�V�\OBJr�'VA&":i�RUI~�q7*�l6h�
�6q���@a��#%�P0�W��k�����)�8�ߎ�tצ���.]�<ױ�jd�/-}y� �s���C�C�nl��n�r������3e�i�$�P�F g�V�p>�[`A[Dyk]���]$��ڥ�Q�M��Й،T��2�g�_OHY��xxD��s��wwM`*-���'wVc8$�Iȉ��͊�ha�n��Hɮ�ϻ�����#�����U��4�0L�Z��gi35��F ��LJ����\�)7�Yx�ߧnB�:ߵ�� ����͙"��p�+G	>�9u-Lm����������j^�7�Zğ�,�1-�^���"l����G��M�]����xH�٤/��M+�-᐀��˛����U�X�QN���-L�V�����˿`�9��z�{*�=G/2�5T�{T0����k�P�2���Y8�������.V��[V,ͪ�M�Y`dnn�'Uڿ�v�^-/J���fC�������Y��D\���0
�� �xx�|**t���,2s��Xl))�A�Gn���p�O��0��P����T��u��{��,/uݠFÎW�gT�H�l��T��R��݈�Rt��@��9�(@�R��F�f��*q�:��UC1�R$��8����l���$Q��� ��[��?-<p�����0�S_�ر�1S>�`dk;��¸�X� yVHG�/�O��Y?hԪ�Pc��������/ʾ�#���:�����s�Y��{��h"_е�<����B�.���,5#�Ԃ���,T<��Z�'r�O=����6�K�3em���Ǿ\�Bw��?w�0a�Ū�
Yt�h����)$�.�ch)�Ͻ"�<4[:--[7�s��P�|C�I,��zj�#��>FR���	h�3�]�nKT�W�K��d���I&}�ޡ��D@ū/d�7q�`� ���@��m� �?Z�_c�`H)��B�)u-�����ǉ%)a�sɂPXXK�8K�p۶�41����鼂Qu�=��:�dc|1&����tIn $IT�m�YC+	�^)(��s�����������z'���ʊ2žJʶQ����9Y��v fXZ�,se�Ȧ�z|� hlFR{��i����{�ŀ�]4�T_�)�O{e"�E/l��kT�E�k��BHZ�)�q�X��^%��f-�o������]�}�$D~7�5ߋ�9���E2���5��i	sOhf�s�t�˒�0��Zw%W�����S6ft=���z�F���x^m�8Օ:�T����.t��@�J4zv�[Q��kZه��ۋ}F��ޞ{�x��wM�=����%�~u��}%	�k���|۞_�#��K@��mk,<�ᓨ²4[�Zm���R��k��N��H�	S�0�&�o'>����/���Rй�����Ǻ�ˤ>�����ڤܗR�	gYE�����|�G�N5�l�V����W/�rU���؆U^�b~�8�EC/�󕕟o�5'���cp�]�v�-̨�
��s�J> A��@�3
Y��J�~����m�hH����I+�p�&&�'Οt7 d�W���yi,�K����K���=���0���4VE�:��*���]L�%hc˹�2�ZE��А�{x�nQgSÄ�#q��N�1[�w
��L��T~<t�w���})ӹ {E�SE���@��O�B�95e��i�zI�j��
'���Mk#\5�5��Hn,J�Ք�a�R�@�
M8��������y���R�AlL_�;k�Gm�,\o)a�k���j�!X��`OA�߉+�O4�O�?��x��<�@�]b�f��p��ܾG(�(�Wa��ԩx�5�cj}���;/�Sڔ>�`���	�n麸g���p�e�TÈo����D�SC^��<����w���9`Y+��S��D�5����S�t�I�d��n<Pk��E�	΢���T�;�:а���A���
����ᓼ�jʥd��=��ǳLd,�-�G�bY�W���I�eDжӫ�[�9'��ܘ�REw����މ��=u�k���B.D�Q�h'=�{�;"fb��Y���b��?�����ɡ-5��t�
)W�����I��,��d��A����F���[��l:r&�y:�
�8���=�B�f��a�,�L�P�@�eB�K�����e⵨�qH.�F����W'�H��\�Fv>��-��}~d��w �S�ؕX�>B�ʻ��ړ�E]�n�^���/*�V�[fr�Po|����{-n�4�l, jޥT2� �@}a'v�s^����0�2di��C�ץ��M4�]^�꺲����!�2/����;	��wqy���<F_����U��4u(�t2��v�fx�:����M����kA2\��D6c�������ld��@{��-Ȏ������n���:l,XC���5�xecN��xo?��e+Q �#<�2Vrt`�q9���R���{{�OAͷ�ZԈ.���Ƹ֫b�>|���"@��C+z�a�E>�e@��ys�jJ�%�����<v�ĤD�r�O��~.��6��*�,"U��rٍ�+e��J���[
m�����	�8�`#S�X�$��"w-d�k��Z�=������Hl�U���De<��Z���i}%h�%��TG�
8�y�'�Ǉ����|����X����<v��ݜD�H��^��,]�9���ǹ�N`.�?�;�<bh�*�W6�5��׼�Aql��Ex�~��)FC���6�,.����3Hp�l_Q������\���!��yD��h
@5�,R(�7��Z��~���b�k��D�3�=�#��Yd�"#sQ�����Z��0H�eH��$���0���_��m���$A�d��mPZµbx��jq%�1Ru��Sn~�4{=#4����v�L�`7G_Ptj��3Xp�ɞ(ு&�a@T���4Ɍg��sӕ����­����:l:�ATR~����#��,��@�*E���`�sW��c��51��M3�,�a��P�����D�ֶ0�]]f�+�齕n��w�Tҗ8
Y�N���<y��9wS��y��*6����$W�%���t���埤l�L
��@��aҵ|�*�|-�T������N�B>��|YG'P4���$�`��n��IG�|�l�K�@6G=��-��Oܯ�@e�$_y�K>l��a\���Ǿ@���Չ�����%wL�\�Mv�N�:�麸��c'$ ��������E��l���0s5�Ѝ����t�|t��5�4�!��b�L��T��O��������D��6�oւX�J/��)�X ʺ�1䃍���b�:��������R�)��h1��~z�mU�ީQr_[_���4�/�t�ɿD�T��l�MhƧŉ�#S,���-�˲:tһ��ѝ�F׉��z�7�V>�n��+#U���g� �H��YƕkAn1z,�n8��9��&Rlۂ��3[�?L'!� Z-o����>�=��u%�a̸M��[׸߻x�K�[�vn�>j7���!1)�}B��|��۸�`��Y�������Rp����|���53���s�{���Oj����Iά]�q͕��dE���
����Z�,� ^
OKm��j���;�Fƌ��d�Z�.rP����\ّ��Ŧ��C�*!D?5�kdG�!K�w�&:'R�� Z�zmM�"���;p��r�w��Ә	�k�EH��d�՟�C����N�-���(X`�:�l`t7�՗Y[�b�Z ��΍!��H�w�mf�����*�EZ�H�Ǭg�ձ�b3���L�̖�#|��	�J_�gW@��bE/t����.n$yEc���U�8iv�VE���|K�X�j�J��)���+i���ˎ�3��)��l���
e��-�N���_�5
�Id�B"�b5
�.5J�1���|4�憷tQ%R��uحB7�)G5[�H��k��������N/]
�h�i��
��ȞNN�o����"N��.�E�Pt�Z���,c��s�4�@��c�]�SV�D����"X>Ǧ\و�޷�RV΍W�� Ç�&��9�2~�c6�E{�gNJ5Yub���}L�O|3[�Q����F�޽@E��[Ó�k7��DQ
��4.���W��^��\O���ƽZ�FӉb�u�B����ߵ~�����fs��<�\R��6Nv���&쒡2.�Zy&�T�M&�#����� �ҏW�,w���G�����y�U�#�8M�U��{�[�>,������g됡bBd,��������?dh#T��Y�5UN#r8p���ϮC+kL���F?�zĠ�g}����F�R�br�5߯�"��Y�T�Lr��o��*��
�36�~m�T��(��vC�N&��ʟ��˝�С��
^ayt��ڒ������2A�������l�H��Yه
�k��q^�&��>�����j�W��b����ßmA�ۧ�.=�<�*uI�ȍ^'�|b�����p�ﻎu	�bc��D�B�~c%e��s���iB�X���q������LIJ��{�q����L�ˡ>�>�Ǥ�{��� y�q���hF�,h}�F��L5mqw��'p"�.k
e�e��Wٕ�=��.�ě$b�]� �m$�89���Kg��E��ї��<����^��ۥ�A���zvfuߝ�U��#�p0��fj��u�?�;f%U���a�IJk>�gLF�F ���)m�wQ�Y?z1Y6܏y�{�l3��֗�X��D�vƫq����u?��M�a�^Ձ��0��2��r�VX�dw��^�w�t U߳/��ǢP0��}jw������W���cPz���d< AR�	L�L������|�$�����A��������xwP�r�d3
q4�t���!}�[3�w���Be�dh
�wwz� �r`tN�J��L̹M����CP�)��0��K�q5���s~�.��,9$�A�8�n��1 5��x�i/,�
��$���FX�K�ܢ�-r^��J^�����0���]f�J�p�'-�FK��ʍ�Χ�:C�b��6bLS@/%ľ�_�mV�9h��N�ڵ�=�5>��$�t�L�KW����~���T\���2��t;����<>W9�����֍AI��;tep��U��Q�����}�"FF�u�n��u$(���k���v�ܻaXZa����UP`%��1S�<�
EQhF�7H��9V
F
~O"L�j^%��KW*��*��T�l��J��ô��+��@�[���_K[/ M*B,:�~���/�&W@��ܨ�F*�T�^:�g�aC�ST�[���\�'��CN^�w����5�A�g�1��Q��9���c��Ɩ����/o�l_�|��xk���,�Y�1����9*w� v��wu���1Aob����7:�	��t�ݷ�kطԲe&�W��'�G�&�a�+q���Zl��w��J5�]���U�W�L���[� J"�db�'����2`enS%^V�t�G�wޖ�;	EQ%0=ߠx�D��UD�d�1��[F���THb9ľ�	&���)$UU��Z�ō�8� 8:���V��.�8_Rl]�~m�������>�ˬ�`_��Ҋ���-J9}k�Oy��NI�rh�n~�W|M���4&nϏ#�/���P�X�\]�CQ��n�����,���&���P��K;F9�d��݀����J����-ש�_�CbL`l��ZS����W"������+4�2qX8oa�7wX����t������*����H�t���~���tD��F?b�k_��m|��	���ڝ��O���%�ꥥ�~ULY���=s��&e����n���޵UK[���>�����`$q(hc\f���t�5P��JTRmW��F|�����m�g���8G����֡��PqQ�Cn��`{	RV�gi{�Z ����)�(�'�˴�;>dFրZ����q��|�4L	��X��e&�G-a#�i���]m���Z� �3S'��_xSD��a�S2��9�]{�0�{>��3�$+��Aɿ�͖��$�%-�4yx$������Sd�H��\j	!�k�E�p)pq��)�=zýJ�������H,i0�O����E�������`�H����}&H|3TL��͝0Y�M�_����yKy�b�%���u5p�V���NѼ�y�8:�me�����S6þ��HW�_�t��׶E���$��I��j�X鐔�\|������v�qј2�hD��3^E����������k��I�vJ����:?���I��� �xT�FQ�k�s��*�.0Ήea�J���W�`U�_�?6��.�E���5�%��h�����}�}�lT�+ř��t#i�[�����컑� �B���M�� zVk��k-���>�-��6�)!���=������W�G�J���T�R��_o:,��w���N���������=Q%����,E_H��6�s4����(�|�žCJ&	����� ��)��|��	�6 d�/�$6RHU�^�IB#g`��q�H(�ln� �+k*h��u�����O�[�	���>(�K�d�N��IR �+P��bU�YXm��'�W0�-E����7;����2#~�g�ϝ�!���kC(O ��d5�t�h�Lz����R��i�|
��N�_k��k��D�3ٖ�*LC d���#���P�(f:�R�m������m�Ta����:���:��	$�md��Mg��E��L�*!?!8�&��I|�ށBw&J���Bk�a��J�ф#eh�9���#���I|mKт��wb��c��������L1f�ziD�A}!�7&�sO���	jm�2��?`��h/{��T��.� �I�ƹ�j�_��O��LB �D����da�b��/pF�hrm5Q#[��Ԉ���"��y�:��o��q��>.��'*쑛�k�w$�r����Aɡ&���N��H�VTl
r�b)��1�����46N("�7l��kCg�����X�@�����@
gw�h��-�9��lu�A�;鑁�ޤ���:�Oϊ���T���ύ�� m����%N_�d/�z�ުl�=~HmU��7�H4^���� =)��3M'X�&Zm:��a�%����	BR�>��^n��>���lm���*���\9�V����a�I��e���r�Y�M"̟�m��#6Sʼ�\q~�+��<v�kn���)w|̋����[���ݘM�s�4�~
ӗ�.��8��M���к/�c7E�A���,��i����yT+{TdM!�v�ر3����8�9_K@"s��:qE ���k��\��a�T�L-]�� At$���]*�2�/^�F�J=L,�a'��X�j�+�~���0�n ����_�t�KD�fɴf&s|�d���`-=����:*u.�����U�͕_����j���l$ǓV����C�Ӭ��/�:��p2И��BU�6-<Twoe�%r��쏜��Q�!�:Y��L�3���7u+��}�[_(����Z �Lp�9�v,��P�l2�J��/a�p�u�m��Ckz,NT�Ք�O��"�>#qnG0�`/��2{��#��FQu�	x3��j[a�/�m�U�CN0/~=�c(q��6��<�0�W�b���C�0����{�5
�#xc#�{�	;����ܒ��$�6q��<δ2"'ه�Գ��uS�q1.���+�����k�[�%ϟS{�'��,1v(�� ���~&�^.WV����1EG-�E|oE��0�p��f��e�p}a2��{��'w�:����X���QI0z\�>4���\�c��&|��)7��%Fj:�;O�o&�)��ԧ=��?6��+��l{Q2/.|��gD���BP����F;�����?{�_����;�S����#�G����n2�_�md�?�-��c��#���=���{|�O��^Xf�gX<��^���r�_��m��$�7��&=߹�;�I4u�JTH�⇎��2|6����b8���G����E�mp�r�������z)�J����LG�)�|9�h̵+�M,��`�iH�b(�U#��y7�������Ɣ٤���N�"��[)g��`v?9Lg���IL�J�6�/fֻg�V)�\�V>S���YM1��8C�Dt\�[z\s�S',�U��LB$���=%�f��kx�q���?�i~�u7 �UE6n�e����"$����>����	[�;�s=u�E3zq��2�o����������������FkL�E�{���T��J�K��>�A>�r�>�ɱ�~Ǚ�'ӵ`���켯�2��	���]n0�C>���.1#(��]�B�m�E���$,c5��4�+|��W>�J)w ~�JAvQ�F{��Mm͖$�~�onhB�C[������j�H_O<�����5�$Z+N���J��j�[b���Π�8��5��Uǣ�\�¦�M����f�L��kc�f��e��5�n����L%R�r�zКq�%L��E��[� O��1�X�����	��
t�����]v0�"�HyU�º�X158���] -�u-T6��e�wwU00(�Q�3��m1gG��6+

������������r������@,k��@��q��,n�@�;"4�8ϒ�t&����z��C��C�R��ĳ����9@ػ밃��Zv&�ٚ`�� `O$�ğ�u|<v(L'�#���;�4]g5bE�\�����0)�A&��g���%��6����Q�8����Q�����[�ޔ���%���Áޫ�N�ΪiX%��=ƒ)�[oHƝ��߇v��'���뤓
"��3��
�XW�4�\D0{]���f���^,�{d��9�w�G|�Ӛl�Ђ��Cń���p��vھӓ�x�>R�bD[Z�3���8=��
��ZX���]l�p���������2��W��)��oJ�i)��A�W9\p��ZHE���WY.!����[�_�JQ����[Lip~��2��k��A�:�w��d9h8n�BZ~��j��yT�d�g�/��š֏74���)��b�,Q�E,5�QZx��4mɡgP'of&�b�2d����iui�o9/�Ì�fC�R�ax$G��5��{���%8c�*b�Y�V4�S; ҶԘ����1 ߏ��c^e$�s���+j�""�t�u�X�A�S.x���!.&��ү�YIO��4��܉��!�D�Z��m�GM�i
H��7�\)�L�'Tf�l�8��
�����uHS�޲��N�\��a��3�x����~����嬖�+���r�X^�)GW�G���R7��2Ð��M$��?�f�۲�;�������h��ϟf2-��î��s�Ņ�&�is�?v�e�{)=����
�h��N5�ؗ��B�}����Â���N���!~��驯�Qj⊨y���a�@��Y��j�S�&2�X���F85h����vLؾ�<'c�ӷDs��U��uLGl���?A�-�/��}���Y�5�hQA��׃}J�σ��ҥ����<i���]��S����Р�ى.�Ŀ���#;<�p�����C�^��r�1�AU)�흏o�j���3g荳u�5YOJB��.��]��2���g�Lh}1���{Z�l����cÄ��������.��d1�R�#KRȮ���H�!�A`M>����[��IF�E���^GkBYGTR:g9��}����� ҋk�u�Va)K~�=��E=�=K�@潊���.�6r���zq�Ͱ^z��i����˲"��G΄�WQp���U���H�U�&Z�[Ua�0����c�Ym�D��I�(G�~��i�g�1Y!���-����ڛɬ�N��`�3u�Cq�aG�zT?֬B���a�o�p���犇p$��KΗ�^��BF�X�,͸b�n�V
S0R��4��~���ltM���s�Z�vHӦ˺U�<��U�ee�
h\���'��0�z���3�Ű%��W���9��ì:WR[�����$/w:U�pk_����ћn�g܄�o�Y'�G\i'�c���88r7YD��s���ul0<�
5�Q�
b!�h�ޠ�Ah��+�l׊�s?���s2�ڹ;�$�=P��sd�Ҟ�熔d�Y�Z�`�����=H�2�)����s���P�=ߋ ���F��}�j/��Rv��j�����y4�����d\�k�"� ��\�3��3wb���
�;���
�T SpR!~F]�D	!��.]��!���3=�
Y��P`.]!ʉ�ۇ|c�5��VŰ�*�Y�L�.T(�*�h83&���h�:�=�J����f]�����oҝ.-gm �pE��U�^
��Gt�ˬl�\Lh�&6X�蛏�]���9��^Gѳ0�ܑ�RFNgq~q�s�2�M�٨�
!�|�
���#3�/;?�̟��x�JܨN�d*ص��U>�|F�M籋�J�	-��|<C[��W3J�,B.��P�T�����䢛�+�b�ԼE�O�u�1� 
�R�s1���yO���(.��]g*��î�f6���#s��e+(� <a��_j����r#�L&v�f4���y��C��%5�b<�@K�ͦ��.*W���G����(�#�맳�so�U��Zy�O�MQH)�T�`u�v�H`_@o	����dd�����Fϑ�6�[0�ߏ��[���8@�QqWӅ�8��U��&��h�\�6����\�	��n�������CT�0��7냸��S�lrf�������^>I�q3��k1Z��N�[�K��$�#o�G���h|g��%���*hk�ܬý#��D���-�u����qi���ݍ+ς��I#8�<�A����!��?��[��W?Hd+���CN�~a�x��>�����8��'-SX�!c@嘽�~g�L�S��&�Q/^.��ʂ-�PLM��/D���`*C)�/������V~h���h�"�EK	7��|Vx�`i_o�3�i��{A�o[4�5mdiC3���
!�Z�O��P?��=�+�S$��`�
@����J?L�7E��!,^C�Z�Z�z��2���`Wy�؀�V��[���9�ir�a���!���t�<y����kkB��L":��u�dϼt,%vͳ�E������n [�w�P�v�cE��j*ݸ;�뺧�@M*k�>����r8Y�B�/�^���Yj���Q�ؤ���p{�
�� ,iV���2W�׶��b�j��+W��m����}��f�I)T����cZ,b�����SA͌���KC��IY�'�P��!�I�p���݆!8!t�%�H��]at�l��O�?����ě�ߓ���aT]���\+��l�<"�Yx���ֳp㹆�7褐��N��:=̈́�e�:P�Fz����>��[��ԫ;zz�]�ě`�r�^�
.ʥ~T.h3lq�����U��|6��@��xR>�������6E�׾�	�]A�1k���H��4��0ApvKPja ����x�X��C7�rڭ���/*�����gG'ܵQ�T��\J�:�e�]|
��	�7�T�K���? ���7f�á��DX�G؎-�\�gmf�����|r֐�`��xΕ ��]6�N`X�#�08z	l�]�������$���W��!�;~�0Z�y�%S�}B�[�N�H��]�)�����