��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>���q=ԓ �AJ�uU��W�i�#*(B�u�S\�mL�9\[}�͖H����F��H=�a(�U��rL�y�^.\d�x�&(�0V��穰��CZOJ Λ�I�z��$V�GVV��oc�z��06�Z*݋�4�ɪ{�BR�M*@RZ;�T�Q�^�\��y@���C��7\$���d��%����#�F37�
���K��o���J<H����|ч��ү��&;2�i�����c�A��� ��w�B�k�O+z�,.��B<i*'}_����4�/:d5��o7##����_ϋ���8��H��S�N����۰cq3qaQ!ֆ'�|����yU�{��!�4����_@�V��)�4���� ��U�#>��f�z�Ydԏ��R���%��{��*�t��re�	>���e|�6c�c�_���y���:�'�4���7��oAdN����:81כ4&��L_�+F3�CSl@�y�j�$ý��
s����q׺�&�Z��w����t0`�l��d�&N�ΌEL�d��^2Q:��acx��9
ogȞK8Q����X�]��(W���}��yӁ���%G�bJ#����~�*�-��f��=j�ӕQY���8�E�(1�"n���$�LR����䋆��K���w����G�_�n��g�G�xDd Un��hD�����9���P0l6i��T�Bh�1��J���� X���
�h�EM�!һ}�uk�r�)�51�L�b�>s+�]r�©}MW����T���1��;I�ZB~�����s_<����jzs�c��l�-��"��ò���ƲI��v���dg��j���$h���~���Cژ�R��<B�$�Ʈ��}p+�$����	��}+�=ӹw�'y���vv���i���ѧ	HUN���`q�Sm`��L~ФZ�>�0�اF>�7;�������ϕ\�����^h���ȿ�f+%]������*��7�J2}�����Mh��S��Y}A�kiH����u��̖�#��Kcs<��w�����-L���y�I���c�7��jAa�A�����"6��R�&Mh�BE五�kf^o���n
11M<��!"��C@��T���_������YR�S�G3�!DG}:Qb�Y�Leq��K97W��{r�`�zr�EU��78h����2Q�1�Ķ��]GI��b�e��΍��Y+�?��:�"ylfO�%�Q7
=͗�q��K	���e�F��1#0����m��HeDmfv57V��G/�m�}�sl'nyY�@���6��@���u�^�~�<�Yl��M�X�%,D!N�qiB�&��Z��%}:��I 8D��HJ�>����(E����o��B�'n�p����_���Y�P���ϒ��
~����-Y,���n�=���t�'��v!D��mԄ��A�.�G�C7��g��zǗ����*�9>�.�P}�GԽ���3���k��D�.A���!��O��|��4���k�ny�� �����ǳ.�ʬ�(?�Ŋ���y�4=iU�����>eZ�Rpg�حģZK|�LL��-��:�]�:�P� �X����{�m�}�cE��3T��a�D�$�>���|{�iJ<Y�[z�B��L��g3�Lh������$��d�ĉ��p4D�p����s�
jx��O�U[��ܯ|	�ξ��������%
��ڂ�ٲ21���3�?j30t�!la{� �`wt�ί��������;���|��x��ɟqq��l^Q.�.I.wFB��Qc���H��0Li�!,Ѳ��$�4�w�I�/�J�rñ����}f�7]Xc����~_�na�H��oΤ�kwͽy��� � '�*�Qg��U�x|�J���yC9��S+]�v�U�v�*	؟%Y��&�cL�\�o�������(�����>@�-���P�Y�C��%�Jh�����p~�^�(o�_����ѷp����W���d��s)䶇�P>«��Ar"k/������Ts�zN�]�2�8J{���`�̌�K
Wi�Q릆n��A-8O"���xw��}<
����Jǽ��5Ɔ�����@kYJ����̴�C%Q2:��W��-�.��iP9���
��F f�ws�1�; ��n:]@h���r����"|�����߅+w
�t���;����i��J0�Mp�`!�<�����Rk�
�.���4�x��}�D)i솻����>/�
�0��#t.��cS_tm⩃J���\��������u���,���(Pi|s2��$x�^q���,.t��Ų��u�[+��C7pD�+?�o:!s�st����мf�[�)�ewl�'w�Μ�@ʀ������$�H�q7z�+��rtƉ��I��p�^N�ߩ��QO6�Jf|J]���D@��Q�\f��b�ȍ��BB�r�9���xU�������B!��
�P�\8�Uw�/���U��:C�	���w$� Ȫ�]E1{"$|?�h+i��$���Ӣ��ɶcb��S��lx��嶅�trO�K4�T��vnߋwX�T��'���F�x�Ǝ�G�ĳol�0�z����e��)hZE(>�˷H����i-�����k���� =Lp܃�}���ʒQݡ$�Z�A��F� �e,sj�p�)�c��!�uy�+v�A1l������J��3 Ur;xj��?:�",-L?��3�o�����Ie��t�Iݫ@/�ϔ�0���x��ƽ5��#a}O&U��[6�X�q)\Q1�O�\���ш$l
�4����O�<�D��:��5����no�0�(gኡ�*I�>+G�oy��|�!�r�d[����>��X���c�Y-�MWcE�כJg�\�j����7R);0�2d5`�Ș�l�`��s7�Aq���nn�:d�*�[�;�>��}>,�7������a�X�Y2�h��1���C}=�eb����x��u0�1]zG���:��������4ؕ6م�2*E�i�:�³[_l��RpC�<��2&Nwb*D��#��ϥ�����& lvt��/����C'�9Q���@��g���X0>(�&�r2�F�B�X<�X�c�h̭��oA��/_��������H�',��v:���$���dT��!��09����p�sh-��igw,Q��|m�u'	�m��s�����ځf�bZ��Nys�@�2��9�t)��>��	I�s?^���?N�.���WP�W>���;?G&y�=�3�HUw7w�/e��������h�A�i��'ؽcֶS�Z�֔Mؼ���C(K��[���iꚃ��)�v���=��A�\N;t�09�v�>_yC"�/ɢ�aR����Z7*�cH�m�>�,$%v�?(������撩�I�J9�^{�:$�k�M��[���x��|�@�-�#�� ����Y�E��g�T ��tA�c��d��4�5,���j���.fVZ���A�/��нZ,���EƓ�|��z H}�����78�G���0J&�S�*��QI>"�=x� Ǌ�"u�:v\����"�T�XmLu�(蟦T�3Q��zW�S��H-�;mz��H�Y�|	�� Ox� �~�BCcBTԂ�'�Ͱ�|�ﾮZ[	�0g����Z�Qm@�|��[��_ԗ���'���L�u��LD?|�ۦsTev��۩�%�(��tK��K������z���F2���q�W,��b���0��H}f;Ҋ�qI<��n<��i�A+.Wo$�HXXI!���{�[ �4]@��J t�!� �:H�Y"� ,;`~�7��N�צx��*�����[�(����߉�]��u�q1�>��L�;x������B�ȹ��X`�