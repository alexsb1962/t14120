��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����'���_����V��ӳ�,{ծ7$e��h���~��O.�S~��>�����u�NI�ߪW�C��·9��˺l��m쓏�����щ��c���r��}���gkQ��
�I�3'S+�p.�~��d{?񮦏�{��G��l��o���S�h�����fP`�p��VC�� �ԥuxӵ�ʒ��(m�%|�>��� n���]�bs��J�F���|i)D��OP�w��TC�6.GcJ[FU�g�Ẇ�s�|���Ǳ��#��s��,�>`��[��b�h/������K-���n�[��8�H/Y*`*k��}^(������m7�!�6���OW�d훶Uy��~g���8�3�ը����;&~�\�\!_�vU����&����y����7I�D�J߰���I�-p�X�|��̚�J:�������Z�}e���������Wݹ���\4��#��5��ѥ���KE��'ˉ�{фn0�dȐ�T Eʑ*�-�
��o4���/���'f^^�����f�p�r���v�]I*�.�xҠ���fs�s�zN��Dɸ0t�-
<�TC����V\{/�g�C$k"a�3�ބ��Bm���m.^��Z�!�g��e'T�jϵ[,���F��|���$&M�@v�e�	))�j���6�]�DM�K��5�%5 Qf9qs)\v'q��3�?�v�������%�r�%ڞc�nL�ÇeƬ>�q��W��jw�=epw����Zl'Q�$�";��|X�_k��e���Eݏ�G
��&�3�;��Iۚ+G���{�@X��Hs�������}��@���KM{���-yԕ�5�BEn2?�Q�9�^�BH���xf��Wi�8<��Z�WG��&� *�~]V���.��g��ƫ)��-���v�`J�P2$7Ķ�/����Цc�R�kkF�Ti�"���<Bgm��؆��>|$&�T
�瞓0���f�YdKs!���gw���6�@�-�a��&;�����w��a�K�j���H|I`,�j,�j�
栄{�`W�=�3=��Uy�D���[�*�������@�X��W�*��w����κ99*YHu�ۡ��V_�4a��x�`���g��J��,0ܜ�j�Uu4��⵪ܺ�o��_sgL�z�A��$œp.�d��+���`j7R��	��:+�`U#�tIf�)Fİye3������Y䙇�K�\vz'SY7��S��r��h��x︍X���<�~j��w�]��Č��zԽZ��2�Q�-Q	TA�l��������;�����}&���/��]�7����P�v�u�\{UovaZ��v'e�4V������@U�~4����2&��"���ύN��[Ua�Hde�
X��辞���a�;:���sЦ0�}�.�ɢ>S���-/3#.=�"��=6���}�aI�}������#z7v�usei�y�9aiQT�*NV�>G�]`)j�"��#�/�&��FL~x�Ӈ��.��`?1N����3�'��12�8j���)�`g��\5�9D�(D��ZT���e6����$�������q��T���!��FQӕ�َ�q!�M���M��d��8bP?�v��>�!}�.�����R-���k�Th�����J�|�j��?��B�ݎI�<��Aq���HȋQ_�Y�:��.�4�t9���(_BV#eo�8qg�ku����%6J�� ����
��y�rg/�7B<TVr,����"����F М���+���Y�+Z}B�1��d��?�CG�o ��*J����寶�Bۂ
�?o�6l���y�+)�)������<N����q��zO+�v؈1��=t@���l4ֻ\��bq������1޷d^'<�:��2�ۍB$���Q]�x���R�Ns�~f�,����8��]�
/jӖ5]
�1�����a�� z_5��H{1��W�iRC�1�X���A�M&cve.	��~�@�*z(������=i���!�lp^k�%t�g���}���+
�R�Ĉ/>�mή�
H����q��w���X$��D$�����y���B~	<�;�e�d�Wsp#Beȯ�v�z�n�Éǻ���	4�,�
>7�3F͎7jz�v���w��5�����9�B�w���]��(�jP��0�R5"��>� ���Ox��e[\������yQR �R9-�{Vخ�g!y�p�s�t�s9�J�>��B�Uɦ���I�9�B�^k�e}�(V�g���U��2�J�7����6Ω�RSl�s`Br���s�[YE��aD�nj� �x/��'�x�{ݯX�Sh����0�u��+��xA,�NX�s.��2��dۘAxs�1}E���GM
�8�^U���R�*ιB���_a5�W�û��#���� ����Xo35�42G�wpQ��^�(,��ESf%�$�5o�Z��G�/'l|�:�W����Љ�j�0d��6�o��\�.j����3�����QH��6=������)l8���������y��v^�+����9������c?��kl�n��CP�ش�h�]H�M�)�\t�\b��Sh:B<`������dD+_��=ň>�ixc�-@+�=ҫĢJ�������ߛ�髼�q1^��Qy����XtJ׳5�.�<}a�����г�pQ~hdAݻ���OWQHkl'��j�&r���|�zgR����	#�	�P$у��,fOr]Y�����4Y���Sbq�J�K��ױŞK��i�[�)�Kg�6���+3�$3'.��@k�#���@?�ٮ�%���#��������;��NQ$^�6��Պ78���[�T1Ϸ�J".��4�ķk���o���JF����T`]{�� H��s뽁�vq'�R�X��-�|�/�J�甚��П�\I���>�����zK�hѢ��-<(��Z��]���Y�5��@�	�B���'�k�°�p05�S�vm6k��ð�f�2��r0������+P X���3��@�2�եJ�w�h2����?�����yaXݿ \��ɶ�C���Qx?iu=&R rT������A�ǃ��R�x��G��R0K=Δ���yk�OL�_�a@)S<N$�-��5̽��O3^ٿ:=M��"8���W'�;�oL��s�����j2Ѓ4�~�Eږ��o){삂d?��&�;��q�5"�79�	��5^���ѱ� <�|>4}r�OcVb�*�t����^��p��]N�ŧ4���_���������u���D�*���tO���w��>\�]��DQ�Zߊ����&3���5u�7yǁ�i���HSN{�����GyZ��̜-���:��H#���� o���x�u�d�:��Ũ6��|7��%�>��+�Z6�2>����|�ϣ����cJ8L��a=N����ݪN{XcS�sc0{�����t��,���H1�k��C���R���NN�N=EY�:�,���_�
 ��:�:6���H�G�4�����*�8n�i�Ч�S;�yY =�� ֈ�ݥk9�Brh�/	K�/�]8O��a��U�O˅Զ�
gR�1�
��t��"U�kT��(�|��c9���A�q��3#+����O͸-H�
��0��>� u�Sg�[�0)!�ŷ��2zl�II�n��:�ȵ]e���"DW^i�����1��5w=D2}O�S�a"���������2�"u����f�0p��Հ�5%/)�z� f�=��Q�E��d���.�o��]�gR߁�J#��Z��� �J'ʃ�#��������0����H�©^#k}��r`G�{a��=FB_�A7��'a�I�<����\ƃ"�O ���*89��"	RZsGM�J�;�ҫٻ�>��;ҳ�u<?�º�VA@��W�K�*�(�k%U��� ��D��wq�v(.���߱R�n���7o,n4� :.9��Z�����\��љ�������DoL�ʔ��Hb��5��j�͇����#|$�n�jޥd?R�՗VG�� [�ߢ��ѯqR�����1�6\,�WQ({�� ����"<~�p>${}+o������~9z�-���8�B�J��������='��u�����䰞��6<����d
w1�b���C���
�s�&}'I?3������)��|�(i��`��r{퀃i�Е.��[�]��yR�?��������:uG��`,� K(ݺ�6�j���V�w �X�9�b
����5i��',�Q����>%�\$��������������U�L�k~ՙC5��)B��x�*�����)�N��f�v1���9��^�������������r��̕�}Wjt��*�?[s_0u� �Lgdʯ=�1��Ȉ�4�c���ę'o������W�JU���(�׿��E�2i��~��rk7Ư4�_;��l�x�7R�H�W�n�I��mc~E��`��B��Ö�V=�)���-���-u��đ]��\����2r�ѳ,, ���x��n=v�Deܴ�BF�?��2E�G��9���2%�;��w��ǉ�V�4|po��"A�)g�#�C#�_.#��i������x�]�ym3ɉN��;�<e1XDݻ��^��
ZC�d�*��
H�ֿr
����ط�򱕮NTƥ5�� 6x���}�=N����c=9<|��r�b��%B�Q�7[���-�Ѱ��Kv��a���񛋾�"[�j^���^u��.q7{h�q�W��w�f�)�5j�FG�'I&;�慽OBT��i���_�$��ۭ��O��	�}Ku?��"F&_f�5��'I�O�o���F�oށ�C�`[z40[��=�(�`-K��r�[�R�mj$�-XNW<�0��C�X�:/�D������2
�����r��2���8E��͵���T����'���8 ��u�V� :��)���A���Sf��n�y�ds�S1�o2�h ��l�^�y�����z3����������5�#�0�x��bĭ����W�rH��d|?Ř 2��ҢЌ�F�MY���[���H�g�r���x�y.�8mA�����ͅ�`pw�b� ^���X{N��VK��7�!M
���o���c~�: j����ڝx*P�_<�7'��ݳ|&;�;:�l�`!~@�Ѯ<;e��TF+�Sz!85�ЙB_d_���~���B��˔���`*B)�H��-a��U���WZ��R#%7�U���$�k?������0��R���h@5u��٥��v%��-��j�Nk����	a��$R�Rl~V�Q��8-�uU�+�� 8���8���}A3��@
Fo�:l����XJ�~tL�'i6r"н.4�؝�v��DX{<�5�d�B�6f�����۫����6�)ՠF����Y�ι=��C�_C�h[{|�#����HԵr�Gʹ��;4:!.󡞞����Έ��b���Q(���e*�d�#���̧�e��̖PX�S^yV�ů�!�xK �����1�P��/e��9N�"��dU���:�zCԲe� ӊD�>W�����<dƕ�q1?��6������)KM��L4��s.~�����g	���B;fP%	K������ַy�����ꅇ��pӓ���	#*�5Z���LF�"�NA)�)"n�wX �٬�2�����J�����=������X�N�g���|���˻u9b�9h�{���-c��m��k&X�����}�kL���UvO������#��T��E���=1���u���iߠ��
����c���%D���*�snvR�X�6�֡�l�I�ū����Lb0����ޯ�7���P��/f1��B�L�tC�x2���0�墠q��������b$-���	�a�o��;�v.`0E��_���tq���� 5j���fD�b4[37*-	]t��IP[叺,FV�׋��șf�Y�����w�#�-�:���Gݑ9�֩�����ġԛ�?
�.��������z������Ǡ���͆�k����I�K�1��\^���l�>�oU|4|�h;�wL7�#�+,�K���W�%���'9ɀ�֘�����S�?P=Fjܺ���XH
z�qk��Q�t����H"�Jn�,���pYw�v'��1�g��3
�XW"C{��˴�1e��1x�=GХ� �?r�ʰDv�tyQx���4���Ǽ��qzb�ҧ⒵���E_h?zڦiG%�!���T����k��2^%��}�!����r����l�^8������X1~c~�&d��-M�p�v̴m�\:E����I�v��p��5<F�2�{B`�-6߾�d�z Ǟ�Kh7g����4#P�&H (s] ��u^=�"��u�-#O.^�o��,���\�g�|�i$�FrG-�->{�<�T~)�~͹�qy����
�r#NC�j����I�a����Ka�)�]�^'�垏x@�kM	�/�ϣ:2#7@��Q@U�j;��8I���5�������
+j�>4�� zT�u���n�(5���o�zn4OG���'��,O*��O������R#`�q�\�o���O_,�������rf��<������V:a�{_{DV���R�i�@o��#�.Y��1%v�hƲT"vx���8ȴ3&:�-�ג=dڎ�\LuN�m.�0`�|h%�v�j��P����m�o��pǬ�04��I�+�E|�j�?�Q�ن�;����h�U��1�61m�Ù�xK�Y�h�K��a�s�K�n�鼖�a�U������ׂ@����+:�z��K%s�l�5D���xw�N��p�ɋz�z�'��%.>�[}�\6�v�Ŕ1���r������ʁ+{�2Y굄������,u�l}V�ҏ̺�|È#*t�[p�3L��8fpf��� �ț�f�D ���?:1�#}O�KZ�m��q��hLx���I&Ls1ig�m�U�C��{Q�)Yq�Ey3�K��U<���t;"���l���=Ul�[����F-�j����nnd�u���6F|@2p+R�=��r�����GS%�{1_qF��}0e�M���ǭ?�i'��bosٝ��z�h8�`֝N�a����KX/ɿ	����]�����Q�w�M@��V�@�ц5�Q}{I������1ݐ������Oc�	���VnO�Tq�<�w�ѯ�������7P��N�41����f@�]�Br�9Yx�z%�W��xBD)S���9�]<��L����(��lTgp�32���,��|zc��4���t��P�^l�1�!H�*p`u���sH�)A
2�b�����E��&��������ষ�	��`\aՅf�L��Y 4��!΢P���6���)\�O��� n&��Ex%r]h����~��uDD,	_;W8��V�	"qcz	�Z�h����
D3P������.�ɶ�)w	�᝖� 2��æ�;�(`3��� mqK�K��u�M�.ԟ�I���--Q��S�#�Y��9Ohy����S�Z�s�F`Wc�����P�e�"̛��?��>�#�a����>̪�]hq9��[��Ɋc���/z���~��}�J.�w؉��tE��\R�HJ����Ozu�T���W�(9�y�����Z<�b��e�;ގ��,�?�;��F�p������-uR3�Y�n�<���T��[�r�٬B�o��-Fځ	ܯѧ�66�ym�\b{@�*���f��s���,[v*�o�����nfR|����.R��-�)�R�V��z&��W�S#�ب�}cuEKA�t6+xU�W�ɝj��ӕ�>�=BH�`�m,a;�%1cV�2.�a0�	J0��x�<�U��X$�)�
�G>�A3e`ݔ�>ۉn�:t-�ղ�·��E���Xl��t�=�߱�MQ�p�������q����]�n�6���Ŕ2��/��(B��הf��lG	��n;�͡v����J	`z�`��%�$�@�lGx�ːgK2��ʸ��YK7-�d���Ur:RL����#�ĳQ��ް:�?�7H+�~<26O�j	e��؈:�/�ô�������D 鷥�I������<A9���S��VS����*��|�/,d�4rE�Y.�U �`:hl{�N���t��� �p�p��:�'y�R�Zq��aE���D��T��S��ɨ$B˅+t#�ꭩ����~6��0}�?V<|�Dn&������u�%cb�!�(AõD!����4arv���MO�ċs�O4�� ��Қ	ld��p G�D��s[��is8��d�E
Fu��yjt�L]#�t$U@o	E���r���k�P��z�^n�|���u��(�Xb��y��'�0��r:�@�:�X�ʊ�������.�@&�������ǈ����/�D��U�G?B����.�x������G?��'M�z 
V���6Q��ji�I�pL�E�O���,Y�҅l�����7ߡ��!=J�n5>q8_�Ϋ��.D9�Ĝ�nU��&�� fb��8�
���K
IƁ؍O܃DT\fI�g`���u"R�o���8��YFo����ŕӸ��_��)B�Za�=�촹;LV�{�"�	�Q�4QU�F�I`�'7�1�i.c�oγ�D���C��r�����c�V�/}��5t�?"W��tT�1P:���������Z!�R�s��nAK�s\QiA�]ƚ�� O"l2��}W>�!A%����لW�P.����L��L��.�v��\�����}}p��U�F�&@��˛�K0{�C�aR�)�al�c��1=�<�}����S�u���@�jN�z��p�	��i�>q����� ��K�ۺ|@����lݿ�����qe)+�)�1~Hn��]Q	b��_�w�q�DQ����ETHjT��!�l�JFI�}1��~�ɋ>3�Q��NN�F[-���c<^v�yo����J���K��7���C���.z蝊���d���8�> �C��.�DU�X	�E��Dm�RW����-���4�Ճ.9F��J*hI]�K�^B9F�i�}N���E�C���Ubӷ�r��=�/̰�yD�:x
�Y5�
��p���w�QC��|��tl����@��+4;)���A��L��:�hק7���:J�8��W��gS��xFg�L_�D.7̢��.��(ܳ��x[�f��F����ֈ�5��BW����k�˔7���]�ir*W,�0�
�r��m����1T5l]��VP�����cR��zH`8����Ш��>�q���س 5���a����+���E¼�E��C3n���+EE��4��i�z�+�]?jͧ��H�8�������I�����1F���K�E�>�Nm-i��ޤ>���`
�(�#��٭�`�c�NR�ڡ�?A|q���oɍ�8�v�w��UNզ�_7! �<�ඐ��4W��$�sd�BKa����N����X]yQS�%�-�����ٻ=n�W1�*�@�n����� �꫌��+�jd��	��/p\͎d�Ff�!�#�[�T��T�w��S�����֞*������%��*��8�y�۝�ZБ�yrXP�.�-����85e|��~�O�EpR�6HIJi�����f����q
��Α��P�Y!�[�װ��~rtp"�rm�a��J
p�Q�)���D�?�K1�k�V˴eL�?�6RHnr��y�Xaz���='td˨���/�VʹWY%W)�'�Z��xF���V��rZ��Bi�ojU<jx��1���-�č�R�VC���%�Q�����8w�{�RVx������%*�=�<���Q��=X+��*�T��\���lwIB�!�sm<�S�����}P��P����T���s�;g����>������@�0F��d��M�:�����aIo�`�t7�3'6���J_,�**�T����T
�O���~��p�����7�1�[�55Ro����}+'�V�Y?ܴi�0�@�e~�M�B��n����<�?�j�<�y+�.�M<��/�l�ΡL꿷�+-�;�O�&���c͝G��=T��A�E�ϐrL�w� �XHJy�+�Ë�~ ��p}��rld9�e��
"�� ��i�:�ﺎΣ�/�KK4��y��_e$�AY(���(��/��;�Z�a�=�5��4��9p�>��Ś�ۅheI!�� @`�=�f�����l��N�I/ǐvω��O��;�A��}$Ο��o�.�b% 		&yEc��m+ǈ��uIGc��(�]��=��0��;���1��G�m�S��t;'��&&�=�μ&���wP�$+�������^�;57=F��]�Wx���[�����w睹Di�O6��lm�R�KīW���Mu�)��3�x`^D�>���bl\(_*�~��zHKv.2oM�Wx��s�Z���o�o�:�clg�SbS��F�U�Ӟ��21[�ϊ|50W���vg�	l�ި0С�D�klV���9]L^��_�����׳���$�l]=�-�Q��������y���s/�������g��y��v�?P�F�K��`V�ﭟX�px��v���j��˸���{�� W1��s9����v�?�s��������W]��َt2�Bn�Oǲj.\�{�ʲIҰ���S�X���q�9��².Z?3��?�Kj[�{�*��2~���M��҅F��Rjo��{/όʹ�x���7]�B��`��"�C�94@Vė�Y�����y�-�?�f�ڠ�8��d�zz��l�FcP�7�)�	��^}lǃ+m;y�E--�F�L��I~�J�`����{(($ߛ͊y�!������D9����)���)�{��ٚ~n�+QW۰�^�[��&D�@n��k�"C@`�A���`�7���d}B "�9��A���F�F��>��N��V������cԨ��kɸB�şv�"��)���;�po������-��(�Ao&޶�����x�=�Wbh~��S� ��'�V���w�2�����(��(h���۔Is�.�tg��3��)����՚Xs�u���de������긢7�0�
�?g<���y���N"�5u��^��~�Gb���k��%�������:n<��ZM�V<�̀<���T��v�)E�)	�!MF�ڤz��Ҷ̩�����Y?��E;�%K�Þ}:T>�{�%�Y�a��y�A���D+Ԁ�~VC~<3���h&�Z�ݞq9V��
����ĿT"T�E�X�Ά����k: ɖ��H��T5�
_!`}to=��{�Q/�/xq�̝`wS7Xz��E(�j�Oz4��@�����ͦ�f{��E�-q$c\�^��}\�jr��tߓ�5�\X&A�Ƴ���.�Kw8�d��{�������7�'ϋ3s(ȉD��C�o��{��H��{� V��5p�����Xp���8MR����:|���2dH��d5��e%#EjĳG����W<�&�)�J�݁Ab3��멳�K~��|T����st�1x�EA.zB���z�L0�UкM��F�)�c졡W�V��02���f�8����E}�o;�}��+�G�ft,� ȣY��C�q;��{� M|˔�gܦ����
�Y(D�@�o\8m�$[�b�a�Ӆ���E�b�l8>�Rt�j�������=�}�0�=�Nk�����'acE�9)�.�bH��@�)�����<b��: ���z;,�Ǜvq�bȠ'+��%�}���5n:Q?<l^p��Tʄa���o��27��Z~�)�>�dXC�&z�6!����/#���%G|^8|c����6�rw׫)�Eڌ��c�A�~�H�{��iǄoE��
w۳��Z__#_)�p�`yu�>:BV?Go�*��C�;���|<�v5���Y�-�0	��M���m[ހs9n.�B�EF��N�&3D�{E$��]�8��Z��w6G����<�ȉ� kkE��~���`��'�Ub�t�L~YQ�*�~(�2K��f�+��.y���\\л����09j��aq����;����v�q�n�_��N5���sk��
w�9�l֝!f�hkB�3Dn�";9鸓�(x��}�G�O���-g����dk�8X�w���g/�0�W��y.mX��a���T"���Ί�Ё�gr`DK8]Ĵ7�y���O��mKn�uOPɏ���h�,2����X7��(G�Kɝ&oe����(k���M��/IN���li���ќ�eN�4���Y�V�mB�l����G��!�V��>&��Tȇ�M@��?��g��Io�i��ܽ{��)-�q���Lno����b�?�`�^rw�����y'o��fC�:Nc ��gF�fՌ���7��%."�GjF��_!�dV�Q���c�,7����%~��P��~�����'���9�+Q6�_�ߣ�d��k5���h��x�T�w��v�����8U�^�em��)0)X`�my��N�a��<s�Go7HC�S}����l⻒ԙO�k&�f���B��]t�>i���K|5��5G�[v�Of:�8A���y�`�^KT�m�Q����8�Q�ɿ��*쐕:�Y�8���HE���A6T��,���bR�����N�/<�j#�! T���3H�-�b_o�y+�w��I_���S,��7#s���}S�ڠ�R�X���9+�h�&�5lw��[���za,A(�(
ɞ9Fً�MW�m)q�9(;^	`r��)�渑�=���i�,�=�%��Ǿ�jͻ��LZ�3h(j7�֘��BS��H�tVf����+�8��y�ՐUw<Υ3:�/�ѽ����9�X�pi��v�ަ��(��+�o�f�VR�3J�F�*V����޼(^�$�7Y�a�݄ؔ��4��L� ��$+[��f����/�>��y5�J��5^�7�X���b���l?
�� mU?7��+�]�B�a��K�U�D������ x-�>:���=E�Z�[,>���yVD����E�%E�yh��� ��p�N%��W�Y�ڲ�R�'	�@lĵ<
�����V�t�Z,2^Y~�ri�m�ހ�G�<���׫�����p9�Ya�n�DīT��Y����٪[ˉ��G��O���g5٦��uζ(�[�tB�WAB�e���s!Ep- �rL����l�vi�'�Gj����|@5�z{-�2<T\
���TH	���ĥ|�2#� �����ąU�ezp �t�$%N5��x�z6��� ��fe��1 4�����
�I��o�Sb�F��ζׯt�F�Lq	M���^��f�9�J���f���_�6o�'�J�N��ɋw��ˣ;�n�u�%�,�����~�r�8�%�^��%����g�ܒ�7DOP�9k���� �v����D���lV0"�,$E�����]�����i��Q���O�E��e����� �g`x�݉{�N�g��G�K�����"h��H`�U
Uمi��e�+n�)���{񃑬�:f݀+��P@!Q\H�2ݿ���+l��A{1�L���M��n;uN�](����͖�ZUs�Ibظ����������t�Z�y��p4���z�)%�%;���6�Mm���k�Ӷ��PGK=���!y��~�O(U��\1��B��?�t6_�%M����7n�\80J�2E������#�x�����pB�&	�ʭ�ʣ�}[�ֵv_��j����<ŕRsm�ur��8�2XM���mָ���;���}�?�/�W �5Le'%⻠���n��1�s�Sт�e����U��C�]�&�15o��N�X��	y/:�x���\�ݚn1�f>K􅆖Ŏk��R��:��k��Od.�hK��{V2��L �T�����J�/_���Ws΃���)�+��gT��=��U�**�_����}�]gC�Z��n����������J����Hj��Q]��@��1�=w%�e!֔�� ���9�ao[���p�.m��S���+��E���({�6��Eg�&��@w�㼎�&N">��!ul�&Uv�ғb�ᡤ�,w8o�A+�w� }�<����PN�eɽ�P��,q��o1��nE$�vo�Sӱ툯���2>����H�Jt��xV�#_>�	�-���\a�C�� 씇8}@M丕�>o�x+�r��bc�Zd&oЩI
����a(�c{֏����D��Й��F-��x?]c�4H�=���dQG�c��s��Sầ ���� �-x5��K�	ҫ��i"ULW�qT)���kw�~�"sװZBv� @�O�?��BS���B��-�թj�Y�O�&� }TA	��R$s{~X�5Y�����QUm2L)Ğ�L�����&%�>���B�e�d�[�IgN���4�x��40��P��Y��
,�0aeS	��m�D�s�5}F��6�DA����;E>�+{�ʑ����D�gc.U��Oo�'D�	(c5� �9�g,#<�W��%��[qErѝ9������e-��l1���u�{�#�=�?d��X�`r�]k���lI�M����	��֓d�c]`���\RT�x�v���US	l���>��F�+�����w
y�k���n`b���@E.>��+.D���lv럓����w�`S�e�)���	�K�$�Zݷb �#i�|,ɪԉ��Ӹ�eu���^��E?��G�-E���"5������Iى_lG�1�}���q��b�
���kc�ŉ)u��vY]k;<>�P|�E\k|�2�a�n`�{��j�
�����w���o����1M��C��Sf����N��">3X(e䡅�:R;�yK��ܹ %$WO�	�4#D���&W�T u�)4^i��V�-��Y��[��>BE
��(��^���{AL
�%&�=*Z,�`��tJ  <�d��Ta��������Gw���R����+u����.�nگ�����]"��r�в	�1����<~SPN��Ǖ�]�72mJ0K[zZ���1aAs~ڳ�Od�2�ZSײ0+��*�/��(wemF��E�U�A��'T��(��.����4�1�d�kq����\V;��<7i��ۄ��@)�xv�zM�lu`/��=�y���H2���X�H}5��K����"�r�U�M�H������|��nš��5|�����[s��E\ ��{g;�!�v:M(<�ց�t� 6��sը��hgrf��f���:�-z
xT.����ā������5�ռ��!y(X�+��r5����o7S�YúY��n=��z�b�J�:��z�xQb���ܷB��� nU�b:m���	��n����r��ʷ
�wnd�x��1�y�X$�b
4�i_B�*߾�׌�!X#��u�l% �7R��� �
_�+�w�y�0ZqUj�4��TXO����@ AyM�4�1d�9�m�
�e����^��s�haY�",>;(^.��:�Z���<�iXsU�ˋ}!��Gq<Oڃn"�g=	~�smza�Y��ū6�� ������6���J/�IӜCtּ��C��m��UG/�L����!�	�j)i�	�Q��򛥡`e�(
�.�.t���:%n'<0;?g���c������n��^��k�矟w�����8��p�7���̍�v0H*%���H�U`���������%���h�����	"+������g��I�u�d �	<^���nv�Ь���[h��$1�Vet��iR�gᅼ���\��x���7��YM�T��/�x�eҺ�to��rA��o�!�b���a��1]mN$�Qx�K��w$��.A��b�b)Vv���� |���6A�:�$�p��r�NA����l�f�����z���5��WW��9h���P�/��/D�,v���'d�pQ�O�"8� ���@`���Ưs>\�|8@��Nȯ鋥�����g�e1Bm54����'c��'tp�H#������-ۖ~�Ņ��*��5�}��'�/�@�R��p��kcq��+��]L��4���m�MR�Z���ڎ��+�j�A��mv�����l��c�j��oP6��wT�{R? ң!@�����3���b�P�mF��(+}�Ykf?:�e�ϑ&�z���'T�g#�NHE#<oj>��u�����|@�vՓ$�;Α�_b�Ê,�vI�c����:��{�9��S�f��M����Sx$`¸��n�L�{�;ѧ)�̰�� M�o����	�,S�؄�/��Ьض9�](��6�����م	�n�}���64���b�s?L]RXw����4��7�Y��D�W��5���0����}�X�]gꌐ� y�2�+{�����
N�`�ۗ"��m�Y��C�� �su(q]���XS$��.ڗi*��J7�� L����t��s�a�z&&t��FD8�~[��h7;hUK���QմmߢݟZ��V���8u���f���a���B0Ya���뽍t����6��h�g }�8`%	7v��W����4q+ٯ��lRb�Ή⧲���z�4���sİ��n*����x��@�ϰ���N����L�S@�� �|������ڛ��bGkV��J� XhV�{c�~�Y�|(�8�<���lL��h@O���gNS��uga0<-���.�5~�=4b�:��F�v���X�7?7f��̱��#�RCغp���W�_y&�p��1��G���ʡ:�2���:�M�D� �%(���Q-�?�F#�����^H��]�; YsL}�>#�6���U���C3�3VTB%��|�ٳ�J���I�T4��_��$5��ׂ�oY�-�<�`�H=�]�9H̕	1M��;���*�3�����!��6���u�7?Y&2�˄
��4]�41Z�3c�'�)��Z��a3�	״��������Ȉ����F̤X �ڴrK���=,[����X)�q!_F�j��^Ϯ+E{��CO���B�(^$�}�^�/�9G9��h���v�������B����V�eŞwN{��GK����Ѻuy��W�� \ǐ��^��'~�N8I[W����-�.�*��h���t��@�D	�V����3��BPa[��":����">M�{��Ȍ��k�9ո���aV	�/��a�U�h������P򩲁����ю;���a� 3�Ĺ�zF����M�ã64'
4p�a.%3J��|�0q���9�=���93��ik�9��ۣ�~h�����Κ�Լp��B�����?��<�j������f&�v��L��TH��\}e�~{z�Ε(�|�>�AɃe�k��LJrl���;u�)�C1Ĭ�0��� =eR���E�����r#�X�4�	�Y���̓�`y�]�Q"�q�O�Oy ���H#}��/*X�T������\�kC�i�I���������v�lr�Sz�xl/�V��p��M'�%��[&��(�2��(������߅
�A%Т�]��.N�,͸U�˺m6�,%�f��[��ײOK��${[DQ��8<���Vr�*Q?^`�
�f4�jy�D�������.X�~V�KLNDQVgT$��
�n�e�>)��v�翁)lo��Z,�
����u���˝��	��H����m�Z�؍���r�8�g@��D�,:�j�.u3����f���0��!���b�����.S�(��nt$�pR��ґ:5�)�@�3��Ba8�|��Hޒ���{�{V�p���`ПlF0�W���$?���jM�2E&C�ӧ�Z��/:Dt䋉���^H;sЇ�"�D�\�,��[<Pueey�"VF�l�SM�[B��q�8�e����~/&�@W����l�YX�gԘ��ڭ��G�R=~5j��X�_��n��:T����b0�bD�A��E�WV�<�	�m��,CKU9'����11�$\��wsY@u��м�E
��x���tзP�/��)5��x&�S�G��8 �[6��$��g�T�"����@�9"ۇ~����nK��K�԰~�;��� �y,�Q�5�&}�Ӂ��#�i�x3��ͨNo"��O\/���`a�|�6��u]�}8?���A05�kgm'�Z��i�j�ߜuJ��G�zyB���~���v���ii�s�B	6C�!�1@�X�����#M������%���٩�����or�̺�Y��	j���l�>݉��~ld&X�y�����В��u���gh�4�*{��;m�b-I�>��q��g��QT�%J�5��(��o&b*���A���m�`>�#mH� � �<�����>���=���B���ϐ{�J-+��\�y��a���i��cAP��S���%X����Iz?��⃐�*�y\[���V]�����
Z��D�=�V�]<����B��$8�M=��`�́�7C�K� 4v�ߍ��n��Xr4k�[s��1����C,`�&A@{A �.�٥���+`7k˶t�L�C�F���٩�MI��|�mr�҆�)�@xKG��m�k�%|V����Dp�BIبS}�Ev��9�x3!�|d��|��vٵI����@2�8Ԧ�-W�b��F�;^�]�� �l��ڇR��>?���͟��}��XW~���K��Qjxa�MLG��MX2=�|��4�l[���c���Y7I��O�`�~.��ĺ���$Q,�WO�|�/�/��.%1�[�
OTD������4Q���0���e�4j�
��0 ���Lzm��c�pv�����>�w���dv����L��|�ŘǍS+�V[V)��x��cǢ�C�c>�me)�Ae����^X"H9��_FM���
J�70���x����^h��O����P����C��9�Ƹb�?W?0a�� �,��YR�%����W�Nc�����rxa�Hii���G�6���Z��^�zlQW��|����1=��F5Ч,��
n�S��v��6DR9	��i�N�|<�E)�[��.Azz�u�3���n%$�
^����Uʬ>Z���׬pV�<������h��cU�>���t0�c���)8˘��p�L%� �����`�R��{5$'*_�B>	~Y*��<g����z�7_v��L��4�؊i�:�[�v�iؓg]��|�'^*c�;�}�գ���ջ>�ȗ �$5�8u�No���T'�ې*
��`QJ����:ox�õ���6]X�>�yYlΊ4����p&���4'a�r�O	��A�`���Ɔ.�Y���#?)�P�����˭篢��"	�����n��Y(1t��/G{�)>���j���Go�J��aq�U,x�к�Lj<�`j��5���s%�w�9[��z�hjO8� GeN�`h<>�g�=R@����ˬ]�q���<��{*��tP�ڋ�ң��&��h�&h�I��k��~�+� �ȴ3b����� n��g���5���ó8�������3��Jm�U�gu{��!����7H����4���wp��kx�D�I,����QK�<�C�%�rx.W�5�?�&��-\MW���@bC꥘wQ�3b�rqg7�/s���J[$�4��H0�E8����p�wx�?�� ����V��:_ok:���ϗ%ܦj����hU�}T�w����߰�>��f�Iָ�O��.���R���/v�mR(�[@d]��cʮR^��X���=!�H��Fx�]��LD�kH�SZRY�
��i�l���[��m�Sչ�ţ��]r�+V$ُ5(5�7� Dj2Yb����G��~�k��x:��'�~�[�j�䬁:�����_ҍ��?1?�c������@���.s��3�0t�j�vLɿGȈ[�U�VKm�4��m���P�C�O~�
��q�o�v��z����RϮ���������dϡPK�G+��)�ܓ24֑w�����55�j<1z����	>4����]d vï��\��yW1��aZ��0s[�l��dy"�>NshC��?����mMǪ�@�V1�XX�?* ����n�ӊA&�B3ܩ̫�xr�8�E4����$��B-�"q�QffNv���H�a0�vT�	�]`E���k1�CH)-!�bC�� J��J%sv�"�,��g,�	����`ob)z�D���'"�T�>2Q��F�@��D�Z�ߌ�W��|{��r#�^p��[���X�N��Zۑ8*�
���}��g�!(���!^�兝y��o�������&� �~�Q~if@y�7K�ޔ��Aya0�C�	4�Qm�|t���[��l0��?���`^��o�~�<�yu���D�e;���	��K��2A��Go�}��˱��vEXI �.�Iyvg\HI��2$Rf�A�\��j��x�"�~�w��?�٪<�7z^��>���x<w�w��d%˔P�g�S~}E�Z�,�Nm��� ��	�:��#����J/����i�6���U���h�m����2����."eq��㨩B �m*f�9-,���lì��sC/��5�g]ٓ��W�
�_���*�~mo6��L���-V�Fi��.?yJ,IEJ��e;S_/m`C^�a2`�M�K)�[͡�y�)�c�]F̞���!is*=�>��|S�����n\�"��|����؄��X�i�4��`�
��NA��jwX!მM��I�aR�9$��$?����}hD5���.�%��%�d�H�^c+%c>�`H ��& 0��8��D����K��th��7<]�(}�G�ܛ�z�}�Qf0y7za6}$Jx��� 
T �����'���"%'�pK~�61rc�, �k��)��d��N�����b@5����a�$%���ݳfϒ�xQ�% ��n6Ӟ:fb��7cN�@=C2/��j_G���m���4����+{@+��h�]1��	�����|��dZHP~�XS`�?/O�+���%�Ӑ*��b��6g ��.���9#�hR
�����l4ㆯ�Q�0����c�vU��}��L��8`��A�:��vb�M�s�y�����`�:`�wo�D4��w����0�EvL�{�#�.:ُLa�a�q���Tp�V�3D������O�"�w[,4��w�XOJ=�������oF�LZ%f`��W�CJ)R�e@��?��au�7�<zʌC`B�����������=#)]<4����@@�������X��@��ͪ�'M�����U� � ��뛰#^c�	֦�EU��5#ߎ_S����u���E�=���n���|���"q	���o�z[������=(Q������U�d��F����L��H{n�Uu$��ǎ�uSQ�	v=ذ-���M;췫3������i��ۈ��!
�"���%B�Р���.a��Q!�!�� �A�K1x�)J߻* Y��E.pUuk��o�E�%|)�=��N�N�@b�N�ú��I��1J�_c�.ޝ6��D)�]��ƴ��N�C'��Pޝ4��t�b�?��u�kاb������;��w��L�ω�#�j�9���	�I�L���!�J��P��]kLGfÛ�=��Z�CW�f3��w]Wڌ�6�M�� W��XFB��i,��g�u!Nw煽t�EB��$�\����Z�v���2q>�<Iqm�p4	�%��|;G�!S�T�7>����i
�+��L�qF��S�.����z���ѿ�ha��>-��?�����vU]L�p�m>6#��7꫄~�&����K?W��9��lG@k���޶�V��9��{���Y�d�ͪ����lf��UIM�HD��ƯIS�]�ߦӈ�t���IK@\������m�t"Ϲ�{���X�ܶ��	3I�ҡ����;3k�Cwf(�.;�I�I���v�m�8���ia�v�hd��@�@�)�*U㾎@(ѿ`�u��Ϊ�8�ư?�ِ�5.��ޣ���O��a���XʄʺMW�N��lNGҮ���H ��`�����J�35���^����1�2Ƅo����1���Z]D���f��o�C��OBk��%z�v�gԫ�A4�;mM!`��3����u!���$x�t;�;dsmB:C�e�)�[)h��������uB�ꆐ-R�0__��T�O	��:mD�}�|�S��r�}���$�6(]&���%���R�C l��D�)V��> ���Ny���v�^���Se��O�mY�y�2� i�`H��58N��9��J�@θ���v��L4��S�H,��II��	qHr�X�	��0�駪���2(&�Ή�R
MKw��U��J�r}�$��y�h��9r��bED꼰�	�����I��q�f�|H`��[y�� �CEs
�K�%�Cvf���y$�K�(B�X�!L����]$��KS��߂%���"Zǋ�3 B�*�1�mvW�h��EcN�|���k��L�0y�K�s-E�v�C;{Z��x�O�*�J�����Cb ��p)C�p�Ϻ��.-v��B>��lء|e�>���iY�#ľD�)�T�*�-w�l�ᮋ�*�7n�� �c����ElV`��o��vE�Ƃ�
�8/d�NS{!o�Ky,q$�+h͈��,G�q��d�&
��N��Ѩt�͈U垒��s��ZQm:��~|8���P�s�&��W� �E�:���\��]���$>�z� %3���o-e]q0Q����]�M����.tf�R����nɁ!7��z���P�����w�!H��>�����$��3Gv�UQ�#�L���C��=�o�>	b�t�s�"w�Y��R  俇� �mٱh�p��~��albP���!k� �Z�+cDS��(.V,{�_W�L���q�K��}գae��t��������}V�.T3�E�-�����}����*ĵ�	�{C��.�ƈ�^���g����*~ZJ�A�1�5���2MS:W�)5^5q��"<�!`��ա�޶%�=��>�y��������(�)~VQ$ڷU���%�D�z�Q.�'4�]\D��if��n�D�3( !
r���|HF�I[]('c�������|i>R�_Ё*|�vMe�7����=`���7t���O�A@�fȕ���

 ��x�ɶ�5p�'���o	K���KŐ^�|[�%yn��b��]����`����Ia�0�:Im}���zy���)��^1ѝ�����|@�"�*گ:9՞���,ͭ�m�@F�S��o	(դ*'�Uhz2)y `�R����m�"@n��e(�d,�F�[1Hk����(���}�Rr�����8K�~^����E랙��x�C�2�Sf���|�l��*&?�K�nW/v$���gOk����-
�̊*V�XXj�Ӱߥ�� g�Wz���Ӳ���Dg4�3I}Hi��\���O�zK��g�J�ҽ+D�s��I���w�XV��j��v�A{E��1L�ŗ���~�&h���;6�덹k��>7�hi��z��@���a���C���{#�k�=����p%��1�]b����r@��,x�'�3p8�'M�SV��!��:�Q�
.�5MF<�<����Os�Pb���Uӝ!'�.S�$?�e�~��aY����h6ҹ�;��|3d	�L�w���\�[K�*3fG B�F���9�i�nHu856�|G#�'F4\&����~����"K�ۥ��;��]�`GK���c9r�����s8��0�^�N�x�
�=�+T���3kI{�D�B<Aks$�(�C��������|<���S�q{!fh���w�R��I�%q6�B�XA� M�p��w^�9i�+_����6���ȓ"�F�%!��i���Uj*�k,���Pݾa���zs6@��`ďi�FAgR�uE�:h!n a�x���Z���oN�P1��պ�uf�@+�뾱~��3��#�l4%��ۜ \y�Jt�6_��l��l"|4M��D��D0rg�ws�pН�?�w/�Mx��5��i�����t�����{���t��ĝ�A@_֦+�%�u&��_��q��d�w�6��&�Ν�i\�3����9�!�cp�@! $?�7�i��ӫ���J�Ǻn��R"t���?�q5c��w�l�G�c��eff�B��l��D� 6C���
]�TA�:bO)M�8���)��N^և���0�ZA�]��)vA�n	e��Q|��a� ��Ӹ��6xN>��q��Z&����1���W]}��[���jZ��7�_�e
��%[��2$��/���O�
ӔT���3j���r�z&��� 8*p�$�ƨ�*°̈́(W�̞��W2���
b���㏪��櫩H�jxx+7��f�{Fkbn��D/��0I�B�Ro�d!9�D��ݗ��dt����\_Ns���o==�=;<ٛ��X-Oj�ǌ��ZPw��<
���G�"�i@�zMN�S��&��DU�_O����D>&WTE�r�����2j��f��I4�%i�\r[�F!�G�J��A�u�����{�$ʿXAB�	6�d��,�cbZ�b���ǡ�}H��E$s	�0^�1�H*\�Y׾42ۇ�e��ǾV@�{B.U��E̖����_{��6B"t��I��_C?���5�:��6�C�W.xy7�8�du��=f�鯁O�a�;0뤖��!��LA����ڌ��)P�k/�{r���Á��j5[����T����
���	��t�v���>��e�Rv�M��:�]� >�0 h�my!�$a+�/Yc����M�y�E�x��U�-�z[]q��W�Fg�5)>��7�)�FZ���7_k��gY_�dͶ�3�@��)�0b�s:�C�*��(�)�u��&�zC��Y(oG�Ǌ<�{Yߍl�qT�Q���_pq��.�|�Ad�J�Uǹq��C8�\��:@����{�sT<�m|�ڒrk�mҐ'����< �k�N������h��}�WLܢ�2�9;Ш��8�D���)4,g=�u�<�ڄ�7���'$qʺ ���9�;���H8BC�MM�&��o���V:c�wue��hN.U�����}b�㸡�����	򉼌���0]��H��:Pd7\CL��2����-��m*1` ��ꮲ��>ӻ�Pڸ�Y�!�/���d��)�)�����m�ul�w�l0(�١�[�"�$��6˧��f��1�׵v��=�o�҈B�<n�z�������2oR����/#
���c�j �[�'��p��VB���]H- �q�W�U:��w�!�7����er~XE뚻mQ�I�%��#�~��I�\\V�%����{�E]]���Z�{0�����P]�:�+#5��H��ׂ�Th�\�R,�k����x�LI��!�~5�3�����?��8��עt��^�L�H��!���'c�R�%C���\��
��8�Ynm���6\�0�;#���2#k�]h^TZ,�� �w�O} ;�J�$���ڣ����Ոe�E��g�O��g�,�������~��"�*����pξyr��D�s�fV+�yh�	����6c���7;����R:F",��[8,xY#�ǂ�^��$3b��ʨ?f(��0��4����xT��)R��e��i����ͱ`x��/^A���M뎳F����,�,�{D^�Mwb�(�����6Z��x���.K7�FP��+��5��ȓ��ˍ�ꀌ�7�Vo/��͇Oc"32"��}p���&�Di��UJ�2k?Ϲt{���*L)�Aq��8?{a{A�������T�j@<˾v���<�6�^Cl�\}S¤=��J�q����~��)�vk��i����bUu[��ZG�e��9��\��USGZ6�>,��Y�B����g�L�9u�Y�*P���DZ��h�O_�(��ʢYiv�㥡=w`�h��;߆��'���4������6���(8�6� �E�#���	�3�E���1�hO�9�`L4	ջi$���V�i��wr���H�C�f}�h��B ����нI�\�@�z2rrʼW���ך�ӛc�Q��K8����_�ձ6x�oU�g7^�IU�,>CH'Uw��2y��mu�eB^r��'�i���뀏���?x�YB�$�M�m�m����g��Ŝ"�v��h~0�J�ց���e�؇ǫ�/G����H���+�Z"y�:E��S0e�;W�	�_̆<D�#O�w��_���٥yrX�S�P՛	�oD<+d$d	��]p�ӹ)lmܨ��]��z���<�A�̃����r����5�R�ҿ����
#��쬄��ͷ��:�D(7��+���i��y��4�b(��co:cG�"�׏f�/�]	�$�AXp������ārîz�g�1=j� ������S�q�7H��G)�m�\�~G����Db1r�@���bv�	a�RFP��UN���)��|��B���T]���B�O�E{v����h�9��Z,Qe�RhI-GZŜ'�'�I,~芆�D<��KsZ?�����C���I���+ �n��i���솊.��"}�����("���ĥ8bW�T�h��C���ׯD��~����@� �dW2JZr
�,�Uǫa� Gv_?��B��?�(Z���ͼ�b�[���"�VDQp��V{�d-�i�W�+A�}˩�|����*f��"���	U�Y���ת�~�3sC���&r�:�#���ֵ1�@bf�d~���!yE�J6��{U��ط�f�"]���0]��~��ᛮ������⬁��'V�5�@�Y���؉�?�Cd���y�$�ްC�`������朜��t�i����\@�֏$;s�]탰c��J��1W��~u"E^�,]D����`��y���H��5���Ul)�.�P��>���*�Yǣ72�RX��;H�'�P4U\-�8�_b}���H3ݖ��Q@�iք��O	�%�������r8�>93�䕫�q�C��j��Ӱ�B.���TRo'�n�]3���D��`tt���!W�_��Lg݊j��&�!qL ?�z���RN�q�S"z�lj#������kiݍ�"@%��=��x�����û��� ��ՙVR䖠؈�"A�hL�E�	~�8]ދ�KWMr�]�:�5��k�����J�N9%w&}�V9-���]��q�g������5�|��/wr��o���ߋ�ɥ��_np�� #���K��4(��S�!�{� ���4D�C
���Z��}��`�}� �z˫�Ԛ)C&����*Mddچd�}HӠ���"�wF��v���=A�`�mJp��o?'�ݒ��/Az�|B;؈���MS�W�Y�O;<�d��LS��j��S-¿�K��d��b���Q-w�E���m��4��|s��5�Be��Jσz��
[�['�ړ�4x���	k��2�A��+�"�a3x5y�"��@ɸ�8w_�M���m�X��v!7�Z��y����_������U�5�uN˺e�q�EÄk}�Zސe7�z��,��I������h���@6�l�k����a���}R���祂h�{P~�ыT�	ݬQ�:i?�	�HL���ܜ����Y�<�Ԝ�6{3%���~����;���9�P�U������	Ӭ[�9�c����� >�0���7�����p��cC8X�Zbih�/���c��N�Vu��(Z3��[u'�H�}c3�/���h�Qɋ@�"5�m��J�D��^{_@=|C�zⒹ�/����V��-�a�
]QZN�+kW��S�>�uzd/�&��| �E�ZD�b7d��H�U�j���^w��6��+�D�h���k�І*�I��YM�'����{9Հ��֤�	V#}r���l�G���Ut���׏\R$({U�P���z�u�ƾΎxR���4�p��wr�ke.�P�ޓ�Ժ�aѩ�/P4}��F�-Ml���ؕ.�v3���w���tŋ�����/�wo�0��f�(m�,箱3�J�m��������`�kT�-��Q��Zj4��&���t�Wc����."���pN|�R�PK�|�H,�`��y}���Cƈ�f��į��%wN���9Eq:��R'��0ӏdx����G|gǩ�wh���(=�
��jۅtW�'Ai
�8�&��a�{B-�����́�I��4.�<�d�3�P�r���E߇�6�_�n�M�f�i�M�_R\34%�ЃБ|�<5,���b�;��-��~5��\�-��!�a�������vG$����d��fuA���{$W��/�$�~1��M�x�6�^�@M<GYjMjkQ¶]浘Ɗ\�i/�ߑ�����r�ʳuG��m~�p0 J��ɠ̛v��
R)���3'ö�_�]�q#���y �y=�i�ߟ�+5��4g����V�N�BN;?���{�(�'�	̎;���Q��;�E,2~�L�eS�(�5�ɚcm��e�N��#��9����|���yH�:��f���T~�e3�psQ9��DBO���o�/�z�CAs>�.>��z��=�|�^��C���c3�y��$p���T����(���h6�ܑ��;��9�O��Qt���.�D`�ҖZO�����M�]���12	f.Q��*�q�)+} 3��Ӷ�>��PG��'��Bb��qg���M��&i�]�*b(W�;z 1]�q
SK�џ'��T�x�� }���c�44q���Ke>�`"Ɓ}��5Jd�I�G�eU���t)�(�B�4��>�ّ�u����/o�Р�+��.��=���|z�-Q�9A�Jꨤ?H������˃�'}݆����([y��O�Jp;��������;��֕��Jn��>�댿�_RD�[Z}%��I�P�]�2)&�g	�f�ʚ���C�^�2�lZT'$�`LW���q{�r,@΍jYX8���l�}O�0Wў����N�NaM �:ǻ��"�[�j��2%B���8)Ff$�o]��(Ӫ��9��Ƞ;	��=��To���H'tY␛���.$����`� ��{=��J*�B��~q��x�[�Ɵ��l���ȏ�mj`��(��im#�!����X���(j9�1U��	sn?I�,H*w��������N�9�ﴤQN�V/x�?-�}	�c���a�[4�-�B��]N���b�U����5a@ú�.A�� L��h@��Z�<�ܢ8 ,d�u2��k��H��b'�l�3B?��"D$����r�YB�~гt�l¢,��8DϒW((5�ŐV2w���?הܴT�فiX��%����Ũ' �Gn=�[@�u�����U�,�|��{�׳AU���(y��p�6k�` ��#��۩�!���)\�t"����%�ΠĎ��i��j�?mU�\L�"�d���;ث>�n}�8��nM$`Q����i������%��~�?���5 u�X�w����]�b!�zS��ɔo�m��M�����L��*2@n~#�G�_
����Q��R���B���_�1��ṜCf�B@pA��pj+��U���5O��F���U_ʦ�eh��`���\Ͷn�E�kJǃ9��R:&��#K�1�'�<�wK:�B�ĔOl�M�����	A�ߣ7�({>��w+E*{��T�rT(k���t���:�(�t�?�����A��h2����J#3"-ZI��ZQE	��w�ޛ3��.	�Ps´W̊�R"s~�ǭ�\X,�b����K���X1�뵺+���W�x�)�*b)�}����<�!�V>��Əc��H�/���9��lDEũ��pBc�s��D���l��T�+H&	#��c��'l�~ontmQk�(r�n��fޢ�_�yg�����ȧ������I�TN��CP�5?�]b�Ӓ�*%�p�����H#�����*(Q���f�u��yg&|����jA0ɀ�-��@��X5�߮�GP����;���U�{��)�R#�N����O�>�촧��_���}#�����l�(Øvb�<T���x���8/���ך�p��/�]�$k;ɷ����-a)�+�C8WR�}��աN�s�b��܃{ȋ�<	"��`k���Z���	�\�<�6�n��գ�
U,�o�,�Z5��z���F��u�6�������C�:/
Ӈ�/]�S�yB׺�2�[�ږ��	��D�~�E6�翚Fn�vY��O_�a��&W��.c��� �{�O�%�7�'�d�Uə�"��*<�	g�%���: ����7:���)���@���������olT��Z��iG�$.t��K7��!�t��|��u�G���㢭��S�fX�(�ۊ~iO�Ԣ,�F����ٗ��q\�d���p|��G6�:2~B+p��dB{�^��5�z�ͱ�r� 0հ�ҕ������J4E��5@6��k���1LF�9H��vAý��{�8D�� #IB�^���	���k�ڂޞD'5�_�Hz4M+��K�t� ���Y�?)��p�x��kݜs1�B���*q�-�LwRӆ������ɿxB�|�}^!��Q^�8�X���iq RT���}S�)�R2Q9'aRk8*h���Cå�l�E��j�SS�l��ظˮ���.���`� ���PZ��������L�Ic��+=t�PY&�MBn9��1g�Q�$A�$L7 V}�O�;_%����gQk��62�5�.�ѱ)k�"x�j��xm�$� ����]�mp��f9��
p��a�<n
 A����(Y��
��$���{�D�G�S��h�]^;y�R��ǻp��[/�Е�pa�6ӟ)���vo<�7�H��!9�����=Uq�e�z�l������(�2�6�P�`r��y�r$^.��7�2N>�Yn_�Th�#��n
��?)%�&6�_1
��U�,�����A3Ç��-�Bd:���ު�k���@52��Wi���fO3�T��^��5�=�s�"9{�D����x ����ʐ��ɯ���{ ���u��o�'Ӳ�&1\���m	��3�ͷ�細��5Å:̮�G�kX�1�G�'R!|��?�f8=@�+N�	����U� �"�+�v��'�L�ˮ+�hO(�<���S���� �����N3�V�]�YJQ+�GRɟWVG��_��㊳h�V�x�]���0�>7��d��O�zܱ��t���&�5��ϱ�cɨc�<g��%�/��ԥBh����n"��&;8q�Ys�}� V���Ĵ�Z��[b�s�|T[�Mb��?�-f�O6�՞�r�W�&:6H&;����6F�!��%\� �b�A���>	*�EL-Qn�T����T�H����q�OI�,��~�
�X�.gm�!�X�z�j}�=\;�߻��mJ�@���smy�E3�wC[�+(c���B���قU�;J"2�ij-y1�F��Y��g��F�T��>PjB�2��V5C��I���8�;���7hh,�Y�A"��FI�u诞�8�w����Y�dz����+nD�I�VϹRtw^w�ؚ�Fa�F�a�I�.ėH���`9�_�!��`�k��lb�����W�z�
�Y���ΟEh7_@���)n#	��2i��`]@�ſ#�nY��m�ZHs<�N��7RIj�=Lz%�P��� �@?-���Xg����=A�
W��������fQX���J���1�l�N=^��F�~Rk�� ��-јÛ�����E�Ό�3}��)g�a��9��5N��F�~�L��4�\Y�2k��Zb?�8s��0_l}��ؤkp�X��SXxP�K%����S�8A��M/��p�,���G{0��X�7�J�Hd����LW�F�fՖ�etb+��d�H�}��X�H�d�p�������.�H�^�M��x-�?Д�� }���v��c��=���@ V���aUޫaiW*�6�B��ν�o��$ʕ1ٿ�-�0�!�os��c��.���+��.�rޭ��s�K��|k�P�W�n��܃�4ƅ<{�ɰ�pŕ�F�^�9d�N̩�(�Կ������z����דҤwƃ��-�+��]����ӸBtX��7��#f6�b�`;��[j�E�fB�Z���]�ҭ�s���́5����4�Xs����q�MقY��*Uh%��԰Cט�ƬYz�p
ܑ)����T�8��u�B��L�b���w*z��*6��n���S��l�!�H4%�'M�e��v�f��
	��X 
%\����:�� �r�o�A�p2�Ơ���~��Dy����m{'��?y@��=z�ӯ�`�Hn�r��T����B�K�4ӫ�'�R�hZ-{?�st]q�ظ'��>��D�_��D&�19�z���hoS��:�XT���m���Kx�H��
���ɋ�Y������?�e2�D�¡]��X�!�t��Sh��E�u_�xn�Fd��X�_ՋP���1��cɞ($�������S3!R�iXs�X�n�c@H%�?����_�Y�%Ps�w�7���Bp巯&R��HK��*�I ��gGຄ�V��\~�ڇ�v��SM�] �%��';�!��4 �BW��s�WC��o�u8��{f�}��s�1� ���e[����䜆�6��t|
5q)�2��1������e�}�"鳷���9~�����#V��'@L6�1�=;uT�`FvY=ڪ����]N�`K|���t}$����������;y��Ј�2Iم��WT�`=��è2�X3]DX��A�%��,�@_��b;?�L��1�Ru����3�L�J������W�hHR�Ͼ�5�^T�l�����v	�Ekb�`�����
l�5:z�X��@�����o�JyLmWY����,���y�Y�1*�v�!�H����zS�ۆy��A(���/kA�b�����7��¤u���g`�8a�!���K�����ӅA����\���/�(�(`��Fwd:l��9��$��q�m��h�_;#ᑛ�^��d�N��c��#��)�ݣ �&�X������U��T��iPO��>|�5cm+DD`u1�ie��`h�$|�-x�KQ�� Ҳ�.�,�:����ﶔN#VqSB�Ѕ�@�K_W;Gck�!��y�v�����K3=о��2��K�
�xJ��:3}�aQ���3:������1��\SR6�Ž����&$�ٚ�X�}5���@ac7�2�
U�t|�}��U-����u��q�Ae˥Z���U\��	�μgP�G�R�y�R��[m{�cG��^����
�2�^O�~�'�/�-�����*
�|j�B�&�� ��V�K �Ed�/�@=��8����z�\a�]���BX���H����L�~�9�fӀp�jL�W?~�j���P�U�������u�[��PV-\���#�T���}��8"q�_�(~��>	��J���*%�b����>�4�Se;�_`�Q�j��!��W�E�3����&��n�K�lu��!�k� /ɿ|��`�*���`��l�bD�[D�^x���.�f�<&=)�C��#K�/����.�s���ʠ�њc�����m����>�
�m�$Q��CCM�$����:�	���p$�s���x rG���'Yh���S�z� <n2�F.��[��?��v�	����P[�O��v���y��7[u~��V��;ݼ��� ��n�P��zޅ�_miǈ߫ �v��w�'�UR�7�֪��rG���x�
F���p�g׿��<��{m���!E8�d��m_ �N�������8��s �H�ݎ�x�K�!ԲD�YC�w\�"aľԆ�f��S��P؋�Wr�{��$���o�E8	!����	�ơc�zm�� JY��"�s�򇽛�E+*e���v7Q�,��(����=!34�%���q�IYqܵ�BC?QF6��{A6�if���|�7B������ ��)~3���Z��mz<�!	 ���|J�:�:�'�-�P���DŘ��j�i���v[��Yo���,�[X��O5b��M
��bL�V���F��^k=)22�䊄z�9|�ߔ1e� �\7�v�;짍�,G�v�!Ȕⷌ���h�����C���0�qs���7^V~�eg�TFlL�����|-�o�.2D*R[3!-���D�
�b]>��;���v� ��xV�R�I\��(����VNOZ� Ĵ4�=��cIf�m�[j�l��s``W���c����V�)0�X�rk{տ�oX�p��_��=�%]�+:��4�>���YLI@�*�p����2���N���'�����[�dM �C}ov	�T;����:h�s��(��u�����R.z��ꍱ�w\t"k�V7|ۯ�2^ɔ�O����^�iw���ޛGWޭ��{��P= f$�� =I�r72һ͖�U3B�����`_�If����gO��^P��ε�^&L(쳋�OcE�^w�{,u�f�E�3�e<G)��hC��̆�{t��v���<�,�M@\�>�%�8BmZP���0S���,'�^�/�x����C �#�,<�*�����H��'$�>0�.�)�����<��D^�ƈWwh�FVő���Mu���0�t*e*D���Y7�K!0���D�ڥ�uK4�2�d�a�̒���OsW�b;�.6J����璟%�L�ݿh���G�v[n���,R��)0��N6JP��zBm�K�����<�5�ߺS����7��8}��o�1�_��3eG�uF\Y*�}~�Ǟ4 �|��=�D悻?�G@�xS���Ez�y:�u7��������� ��&�`(����~K-\�9���=�wX�*8מ$s�}��c��.�9�W�I�m�7��ޡZ���e
�+��8����Z���s�/���<�9�Nq8�fY}�ޏ��	2A�	gp����C����$�B�Pq&ߏ�r���H$���b�A�ʇ	�oEe�7N�RŰ��99�",��L�P(&�jc�l�D����5�[�,�;.�t����>���|䎠�Ѩ��)M):W����)L����C\shљ�J���bl|�b־;��G|�̊�~K��e(����JG^����Q �TR�5�c^M�S��ӎD�q�ЉlS�Pe�zܙ����L�"�׀o1 �U>J.���[U
�3�P�����X�_�m�=�(+�B��k�en�i!�`,a�t�ๅA@Z<&3��`��oiG�f�,��ClR6���#�[��LË�K,ӗ@���3G�L��^���_�����Θ�]Η�����H�3}Us�sE�pq���B�K�-�;�x��f�zR{
��t�����B����30�`4�	e=�[�Ca_ea|I�d�SSC���紌��X�8�q�g!�*�U�+ɝ���%��D�0`��S��DP��q$�>� �����V��K���E�`�����d�U?߁�M�R�l_�Ɛ+�=)R0OD����G̣�o�7��q�Тհ�e0:����k�I����As{q@)��N���7�&���ѕ� ��zM��]�?�Q���M�+c5L;��F��.�Ѧf�`pZ���;�.�)�������&l��F��N�E�iL}<�W���S�;��D�u'����J���"���|/+d�J�t��y�3���@N�4���	3l���fO�I4��6E�uAm�H���!����q����N�-w�f��H��|�V:�� �*���Z�}z�7M�ޯ�:���O�?X�Ji��|���<�U��"O�i��S���B�	��v�R��>6��kWZk?Q
N�{V,NG^8�!*ϟl@��Q�C�!�Z#�b2�vq�v�A�vE>܀_*يJ(EZE��D{*����D�[g�&�,�ز��Fh�LE�,�J#�:����x�wc���mB��/��i�� i˪���M������d�Π�:/.�����:�V�%g������ok�E5ĕmPB�������؋�V��yI^^��e�j���4ؐm�9!'��?����T~��1*]U�{�-��㮁����]ְ�~rX2yz��ܱ��E�c�VJ�C�f�)$��~�"���ξ`��i��l�p�w��@/ŐS�s���;0qQ��b
�7;$R�ہ��d���.��#�ϕ�@�f�:��-����Z�O*��<)�_�����0�$ �����PTYʻ�[mJ���A[ξ��>K���uI���k��|j���2	odz�}��'/�a_qE�A��2������B��{��P��]��V��dH@"�4c0b�2����\k_���-y!�$�M���,����$��F��9�6����|����(N��r}A�ƍ��{X$׿4���&�'.a��R�7�DV>�~��Uӿ1T<gE9��,��E�=t���#xL��Zn+ZR���"���6��m'�w�?�c��Z1}5y!}�ݴ��/��Km��L���^�t,��B�z��(�N�+|I4�H}��<�V�������ZcC��if���7�� -8(Z�ad$�������{=t,[�6"	"P-Nk����ӣɜ��S�^�QQ{-=a6N�G�����ڎ7�V�4���z�P������Pd�`�E6�[e6�zL׹#3`+� m������k����i�__ô�R�ώ"�w?(����?�}���$�@w�i3E�)����@>pwSj���y�]{x2�p�@��H��?GC��̨g�~_o"r�&j�fj���M�о�}aZe�5���)hj����n�4�>D���2�O�/��j� d_Ȝ�#����\+T�$(;�s��dV��^z����k���6-�o�j�(u���x\'��H�����-�|�6��cVCYӏ�U:���]�5J6̙}�#I%��"�qV��~�u1��^��;͐G�J�
����->���e�y$h/�T�e�����w�hj3Ԏ���R�i��i�z�����<�NXR
P]��퍩c���/����)���Xfggu���%�ѓT��!����ę%�m���2#��x��i��r�����Q��,d�Gj_�u�t�F
Uk�s�A�����X��g�<�%��Ԣ�ـ��[���T�įpP;u��u[�c�
���DÉ��<��e�������f�Jɘ?�ru�����Z&����C
�2WMr�^�2�Hb�� "� 7�1A��;R��PV����s���i>�`b��$��Ь;���A�;NEV����ɳTP�V��J��~[�Tˍ������Z1�~�f~܏F�i��2td��{�7tQ�����)�2�E����x"�s\�;��'^F<�<)$��&�*4����f�=A����	�؊$�/��շ{"��U1!������]#"N��d���V�Y%���v�{��f�V�[�yv�+�D�~T��:H-��ҊCj����"�r���2��=Py�mO�m۲�֗;K���#C�G;�`��N9ܵY*ͤ��:�42� �<qZӵE<Y��/�x����١�rs{�(���( ��^�cʐfYQ;7$l+?�ɿ�K'�SF& �R�=�҅<rT��xf��],D��h�fZ-�Q�E���g�@³V��A��]�aBQ�*t����>�����)��O���+�nJ���}C�;^�K�j��]���5o�G	}�s���n&Ƅ.��Mg���Shۘ�KI�H�8n`�r��1���kA�4>.��)�A����N��EN�5!Gd�!}5�������F����`=���F��Հ��P�0%����u:�����8Z�<_\�r��#��1 1�z��cg��ǵXkJ���@��X�b�$kƷP
{R�8���֢�A���ž^к�����unP#�|V�|=I���\4�2%��=F
����aN���;
jy�y�V�����"��:�}ݿ�P���$��)��4���b���Ȗ�=�b�(��j�]ٜ�����Q���lF�k��J�Щ��­�m���`_��\�c�S��-FCr�ݹ��u-��yF��j��o*ѧ��>���X���Q0Eʑ_��}kt��j���%���:��X���O
��;�Z��>2ʷY�" i��sW9���L�`�UA�ס$���Yp@HVL�XI�@@�&иU�a����x�����Ujْ�Ft<�N�؇�$Y��W��:�fFZ.�<�5e�]����2�D�_2d�V�pb>��+x��"�p�Q̠����bqL�T��,�VåŠ�x�9}��ZqĶ����6����N��a俖��
����a����A��o^|%��xu�$��:$�Xw���@d�iC9�����ps�@A-�S�հ.#UeG����DLX�Ɯ^yH5�3���6���U��
>D��r�9g4����|��,�3�%[�(�刖@r)�ɢ-c>:O)�F�L_��C�Zt8��!@�D�ɓު'ICN]��1:C��9,�C�|Qv(T���'P�Z�Z���m��؋�7�:3�
�4����טK���)+��f�b��τ�u��Zq�{��|hz�]tؓ����'y��Fgcf�P���%	0�u�̋�(ϐ6�mɌ͔MK�ZW��|�ڥ��~x�JO�faA���XZ��pW^�b�o�)O])�څ�B��j�n�P2�ѽ�u*� �9m�$�/�.[��i��U�:��L	"D@)�ş���^�iq	z�#.�������hJ;ʛ~���w^Q޶A��7J�"�����7�1�+���F�}��_7��| ��4��C5���޴�ҧj�������fә�1B�]Å��^E��x�&l�
������ӓAb�H㠙a}`kp�VP0�5G�������|�-�I�lM<%��fVoŭ��nʱ����J�Q�`��@�y�@�Q��I�N���s=S! |���d�3�ځ�6cZ�蠗�uh~���)�#?��ZM��$��\z.��E� �9�<����L]y,�,�Hয়�':m��W3 �h�s̆q;�"�wp�M
4?/��Q,���Ȉ���\P�%&������Ѻ��k1�\ � ����ѝ���O�Y1�!�������ws6�`�Ù�l3������{��%��)��ǀ}��qɍdAЪ�d�F0���J~����Ml%��(@:~|�V\	�Q�̈��_�^�D�[�I2n�q�4�n'�ÿ�Q��`T���n�ȁ,�-�T����2�������<Lm�p��L���d�����js'o�^K�[��z���n��)�����{�zː�~�m �:�#���Ësh6Ռ���g��ܑ�̹��e��ZG���o ��:�Ta	�� ����y�¬o.�G��4�6 ���:��vn��	#E���h>���M���!��A;n�m�9�P�T��w�R�a��.�NX��7z��SO�2�����k�o_�z'��V�~��+CdZ{,,^6�]$�ڴ쑟�J_�� ��Ա��g��i������4��eN`'a	�I��D�nz�BNЖu�6y}͜�If�1;A�piv���+�&Z(�I�y��?~i��(��nIT����;Z��:Դ���IK���;E=�j�W��N7��ftH^]�Q��P��T�4�cbCr�(ڿ�l��ŞI�.l�~�u�Qл�I�Oئ��T�Y>����&�ۮԤ�;Y3b�i5��P)cE��@�}�s�]0����:�.L�r�:����N^W�龆D]p��_�'��1�l��V�fS�gƶ�pt�K�d��g�mO�K�.�5Q I� �<-�.�_T�h�gCn>���q7���2��5�&�����:��I�Ϡ��/����c<B��Vd�w.��Ѳ�_���2�9�!�.h�O���)ϸ9�5>���TKz@0�V���Fk��H�'LH�����.�&W����S?F�V�E�b�}|�k_uZ^�L
�W���_��7�y(�����4Y�z9��$�5b�%�F.��p�̀�FB8>��$�@2�I�rF��tH~dn�@�+�Jz}��.6�Tᚖ�IJ�^`��)<\-�t~_�������.m�v��&��4����O�$'lE�a���*��F=�������z�.c��wD�_ۻ%��/� �{�Yk�H4��؛�U�����i����ߛe4��z�2]���!J�n�j���4�@孌���/�#��������U�޶G�H��c��1��S8�[cLu���ٛ����OfV�3��zk^6M���r��7��gO�hY�,(��NA�'���w2eIj��3��n��>�៭ɪ8yǡA�����:Fc����7u=�:�Y�E�UP�K�|���0I6�9؟�'���I�Rz�S��)f�ִ`Tw��5W�H6��	��`�-S�����H��`ȫ���M NjG�O���@B,eE�x�޽O����t�K�.?R�PX�|��}$)�a��m�`K���H��,F��S(Y���q��s'�M���K���D��1�ݴN�T1��0�N�2�c�������t�C�Cm�ǋK$0��u#_���Q�����4��czY ^,'O#[r��R�{vr���8�Q�|�/�iK;�Da �c�)�c��/�<�����Q��]�T����#�&��ʥ��%�c} C)91����U�V�a�l 6�X{M|*x��ZHYװ��^�_����V����l�e�>�����
:�r�ccK�� �f�.0�F�z�+)��k9��_�ȿgbm�򾰶�-����@`D,oc.}�QSe�df��0k^9q�EM�k"��o�=O~xϳ��@�%���X��^|��1.`F��S}����9I����R�u��������x��mr���Frߍ'�Ս>�.�~��q|�	9�g�RKC<D�����W�+a��p���3�*@�^�����i�2� r�1�oA�G���g�X�ሕ��t���h�nI�z��y�NO&Ƃ�R-���I>���,��9�K�ˬV1�b�������	(#�d���E�%�4zᦻm�-l��y����V%nS�O:��e�TӾ%�5a ��L(*���$l��Sf~�����$��Q�T�냲���c�G۾Qz|AC�D�h��Y8���*���4�H� ��2a���uU���:>��
��gA������O�
�|ET�$���=X<��X��u���Od
�_ʸ�M��BF^/N�|�w��ę���=�~G�V�*�q��к�s� ¸���剝w�j��d�.���:g��0��Fp�!����Zr0c��PHը-���{��9�E�?�/�(�����вO�Ƨ�����]pƲ���vTs3�F*1��q{�{�1t�������7]�h��zr5d`�v���wu�E�er}��,QY��� ��%8�*8@���9�kY*��:W�c���{�E�t����Ǽ��s�Z�ϼ���
�жLOA���%td[n� ���	�W�G���8-������R�v�B����-�|�{a�_�D-S!���>����~�Bqz����ӆ���r\��րh�v^�-��s�����v�#�6�%��& �9J�7	MG
�h��Y,)�� �G�M^��fp���^]{ςI�^Uo�y���"��q�Y,W�]�eq�<ǜE�Hv�"�p;	��&���i���
3��C�Y�D�i]p��9�f=��R���-�W�\L7ʭ�u,������x�-�N�Ƀ�LY����Kq��M���Bχ��oez^��yy��[��������R�b+>��%f�|�\ VǓ��b�^]��2Ǽ�;�
n��/p�x��+�iݗ��F+��>U������mU��q\�����T
�.p��E[^!$K5�����򰘯S*t��0��z��CK8 #-�hY|Ln������Ԗ8CP��Ŀ.@;�:�����f��������w��q"���\��"����&,�l�$�r����� 3�G��'I5�%��p�w��b�v�"��F�7����^T��Ц�b�K�XN��A{�Y��iVڅS���%L�ˏ�+A��d1�lǟ�W�.M�"����632�g�lV�-4�o�M��Y	�R�����.����j��0gs������.����P�NWT��=Čc�$��.� CJŲ�LUy�r��Kk��7[@�NC���f]��C�>p��������[���L���N�-7� �$���r�m)=��,�DbW���N&;6�
�>�t\��Ɩ,����3��TѺ�f[?�� �V+����q����x�$���ߢō٬���� "Փ�*b\�J蝄�P�������3�/�p�,��[�M��?ڻة5R�������ܙhl�̻�(-e�?M���B��g���CT��6C.�d������(����(��|p�R����$��08��v��^���� x�0[^�YnQ.���UR�����uWY���wz��� 5��roW�Ge����lMi��2S�QN�ɃČ�c�E��+�T��UE+���mA���Fh�F`�լQ5WGơv~�X���%�i�9�K�����j�����l������閅�Ȋym_-�b�e�����^T�
04������L�p�o'�$>yV�θl���v�X#��͓+��3'vg�����M����hkv��g�``5�v'�߯]f���jc�x�;ʭ�L-'v�8��+�@��aDD�Vꜱ��5nD��'cc��b 	�˶%�(n�F�	R��1V�߇�3� /�+�v:s��x.YM�K`g��������h�~p��y�K�[M��N�<�~!��A�(6�ʷ�R�N��Q14>k_+@�tnV������?�l+bvx1��aQ`Y�3���R�U2$�pP�IhD$FI	���n�\2�F�_��߁�Q���@����>$�5���2E��ᚐ��H��>m���y�� .n�����e��}�+��`:�����	�>)˾�}a�AO�}D���=Tp����ϙ�$�tN��d����x?�p����S��w&E12E�	i

p��к`Vy�	`D����,�W>���3��B��Oi���{���~X;�T�0�Ɇ!�B�1}��S�u;X:�lq��?���n|&L�J[�L3+���{#���6��K4�@=�7!H�B�%�+Q3�d��#��WIL�̈,��G���7f:�w|���D"\Y�bx5�#�nE�j���3]��y�"6�� _\2*Qvj��aO2��;y>'c��J�et���Jϣu����F�G�).H���=��&�����Bמ�ܤ@P^�o�kK���\Z��>�H� ��I=��U����7�}w0buvQ*Cd�zäL�q���K.����::�,F�栟3��a{K�6�K@o4q�ޚ�>o�V�{L�zǫ�̛Y�pA|��	�a����Ӥ��*�fDSUދ�ٟ��/�sʦq��mɐ��S/a-�"���ѵ�ޑ��`�xN&)�"T1��r��V��i��'*��e�"�)[�3��0r�V�<�<�s:Ԃ��j�~2�����vQ���\\}�����R�����`�ž�5zލ~@(m����1r�m%:/Y�O�i�į&Q�-��H�5�X1������0$��T�^�JqI��{K6�d?%�G\�2�Β,Pט�l������O��G<�`$Q3�v#u�����*K19e��i��+xY�L�2K�K_��ԅWY��s#�De4�m��۬�K�g'���g�1m	���f4�:��K�A%_�����m��-���jP}oǝ�p֖�s�"1R��0XV��h��(���x�	������}�1�!`D�Ye�Q��
� q��OGm 8��<E�D��S�>J�N�sdՂ�]h��Z��h�O�.�3ޯ��͜m�妖O7�>M�VV`P�2�$�2$�GP�C�ӃaI���{��v�c](��[������\�;��xdd�� ��'�)�9;�����c5����ų��w/C+�'5��d�����؊�5�d������V�a�̶m|���4�8�_z�z���#��R=�$P���&��-A��V�F<m�n	vh�J�ѥ��O�Q�㖜 +?Y�芧����F������e���YF�,�#�w��R�hFQԙ55m$���L�;��-�����/��4�5��ODu��a5)�JZ�X���UOI��m&���M�&:�Ld����,����lB/��H�]kM��l���5
 Ҥ;&MFB�N�a«��C�S?����wA05��CV>�`��ŕ�_�4���q�F�]���bd;��*P�V��ʐݷ���ҧ�������>��@i4��[��>R�2j�?m,�dc1��1ʌ��X+1	ᴺ��[z��$k�W�]Ï�>%cS#�¢����u"}�]�י�ꪶ���@I��/e׽��yISŷ�P����sj�`�O5M��$8�%yi�.G�e�9,��n�9zЕ���p�ǛI�<�V#��0�I@~ �q�ok{�"@8���9��ԅv���;'AL�P"������`�`V��_����M҂��/��/�!D?�i�&}��'ʦm�l�n���h��A7;L�W���=��S�����gj�vH�d���!\��M��8�9�6�Mu"-�6�·�>	��F�B���=���1f�'4�4V��%q�U3d����=X���8jx���$���A��Te._#5�|��n�cO�J8�?�Y���O��>*�1�B/	\c�W�x(av�#aU3��O��IMq|��+��H*O�\s>�{f
e�� �_�`�gz��o�:@P�-7,�P��;�e~�b��ІH�4��WD���mYH�1��>B��[��:gx+#\�f���E��u*(r�>��4�P�	3ynO��K��ï��Y7�Xכ#�B&i���vɹ�F�ߞ?v�<)�⤂��t�{s�	�5��"���z���1J1�}U�&��i�V��%dq�� m�;�Q|���pU��܈�j�D@���~p���9f $Mp^	1t6��O(Q|�H�m�I�X�E�XL�O9�v�\�[g���+|��m4�@wD��"�t��ȷ�v\	ბm�)�!R�~6�Fn?q� �ֱ8b.��D�o�ͼ7�=���x�H�)B?WV�#.d���gLT����+T�M�z({"
vC�������V�ٱF�I��g�E�r0�;�)��y9]�o+�<��`eM�XQ��!���AfbYI��"�Z`���2z�L�J�ɷ@M%�kC���^+�܌�~2eQ@Z����2/G85���i��%���N�ڱ���鶖(j��,�ˏp�vKG��q���T�7x�N��LU����E�x-�����:VN�i�O�3�#U�+2�Dm��^_��b8�#9G9���ثp��g�I�z���Q����{"�Ȏ�S���'zSk"p)FQ�
�����v��d���*m���E<$�=��bůN%�`"�l�����O4��
^�˹��B.�(��4��b� ;����nh㝆�a$�:�99�Y���Ƨ�F?*ol�RzoO��Ͳ��2,��^��;��:0���I��'���۩��a���abu��s��4���Jo�H��()A0�y��p�s;ڧ3f�Sf�����@s�M�uF�iFK6��lΐ�X�V\y{p���\��C���w�F�E�� j\3�f����>�D0Xs�i����}5�b�	T}�>`������Q��ښ�ByY���mB�|k�����R��o+�&M=D� �N��>,��4�N��Y|'�풲d ����wR���0�إ���[�W�-�ۮ�kBˢ�;�
�U[���&^)�`*��Wι$�)�U�ط�ʌg��j����z�?LM��'�H�<e���R�A�B�J��33���2��.�k��i~���*s������&�}}�t�Y�٫���R�#��wEal���X��l�V�� {˕�*���(z.�d�ڿH|�w��u�=a��d�L��H�^%;~�����Y�I>��O�A��m�Q�8�PU�b+�y��Fvs�`��d��[��̻JgS�9��7����s����	5j��R��S��8K�6W�����������p���d��>h@�Џ�>��_�W�b�<2�[F��LZo��浏�W�čr���g���y���� _g��>��Ӎ���f��Fs��[��������4T g�}o��rѐJ��ip8����_8����Wq�!�q�r��t�N����͆�t)'��RFoFC�=ڐ"����.�J��H�z���n�A=� ŪC��}4�cFyZ%Ȯ�"�CTk��qLֳ!�a��舸��o�c�4���^7"K)���e�#���w�PD'=��W���O�_�q;βƁ���_]7Ӷ�"A�6�g�q�AHq� ���'����Cȵ"o��u<4�������
ȖI�$(���v`��X*�#Nr����j[<^��7�U(�fz*F�+ �x��[�^v�����6=	�J���̈́����B������""�P�N���C��m*F�?�;YÜc)Ci� �z6�ն�n+Z�9�O�uX���sK�,
m�b��r��c9T�����*~d(�9n��3Do��B�f��v.%����
�]���u$#�����\��$�]3ś"MclӐ���u��$���u�W�r�����n�����@�w��
�y�*��t69S�e���>s�V�l�o�y-�"�QQ� ��xV��sSa�T�[��-��^7͠Xff᪵=��T8�4]�����c��`�y�Ph�8�,�۹d�����'�����]�,�@'Vxsl�*!P�=��J�U�߅�i/9m�u5��*�dQ[��w;ËkI���9Q�ڵ�J�W{�b]m�JP	v�	���饨���:���yѢ�(��k�U���@��^~���Z0��E����i��~="͍���gî�2�٩��@���r�ھ�q���mI&��@��#��[v'azA�p>�Ai�Jq�tO_��!�t��/.��ƶG��sz�~.�k�m���K���eH<Va-#�܄u 
����D���j5�8����;���'��SH7���8q�ibqR�듨��pPQ��P|�L�z��u�,�}zQ���_)V/�ͨ�ʓ��0�7 �0�4DQ"��dr�+LנS6BR�4�L���к��L�?�����H�F��a�j��+�5r�:��r��$�`3�Vi�EU����ʩRੑ�Z�z����ڧ)��!�0~�(G��ܸ�B���aP�?��'��'5����@yڞ�a$���:�"��"'����>?��yŐ��&�/c�����&��#!Ϯ��/��y���A��� _����n��մH�O0[��S�H˭����ܲ��
=\��,��fw��!�U��Y�XHP�Ս:��y��[i!�˂�AO�������Y�A�3gi�A9���E��*0w*�:��m�Ԅ�2F5�.A~�R��N<��f�b�5Ax�wH{a 
(a,�)P���z�w���C������ ]���`��� g�����d�ߡ�Bg��r.]9E�%L�g�B��I�#������1�x;{���c�㓶H�O���K3���'��$֔n�;E�3I}F/�p%�E��!>��l@�o�^ݿ8'k�\��h�.=8���d%��[�pT��R��SPDR�zr
�9�KV�����%Ҏh���'懙����c��[��eԣ�=��&��%�Vh �O�f��dl�Xi ~��w?�w7a���{ݚ��K�/CE,�~&�5��0'YYI}��}W�*�9N�j8��?s��:��1]ԥ��y���j���C)�U�G�A��oJ��ﺖ��[q�o�m��ǩ�V+~�*Co�BQ@KLl0M���j=h��<��q��lc���ދ��;���=���6y��X�֔�����1XF��l/�٫�7075V��c�YB!���
S�A��I���>�qp��3ZIvڇ�]`�X%�G� )���p�7���#���5���"���ʒn3��vz_֌�u����c4�A�s)�U��Z�2��������oƫ���e��R⥳�ǟ��L�]���������
�W?�ȕ�ʬ/0�_ǯU�ZX�A��(���)��E�`�*��;�Zѵ7� p0���,6��Sg*�3��T�_�nʡ���R�Cߩ�z��~�5�̡tG/U�C���p�AE�*>a� �<��=J��E�C��-��oԭ鿰���cKZa�nt�sY2ɗ���W>���^�ͦ;U�.V­� y�i�x�q���3�	��x\���m����Z�b��t���,%�x%�'�%�9HO��F� �
إ��8�z�:M�^�8V5-���z�=���HF��S���z��p���h����[�V9 *����gi?����d��� bz�W�m)�s���
�w�o9�����%��ؓj4im�ЀTR.V��Z����
��?�6ۼ7r N�CA�엮0(=��-�d{���Y��,&���,��*��/�c�@_����b~lL�B�����h`��LWn��������ߕ��	]\�t���J�I�T��ϕ��5�i9�!�jah{XF��4O�󭅯U�����ɰ�3R�oe�X�#�` -	Yp���7R2��g��*"ކ��Vkd�4�r�B�ߍF����]L�?�� ��P���4R�W\2>N؏yF[ئ����ٌǿ�$�]�(�AK�Y��"��k�.��^�!� ���Yi篦������!u��Lu�����NUG;ķ<)��������SV.�{ۃ��Z��Hs��[(��{C��j��t!w�q�n^��3[�K&�ׅUSz�&������"�F=5����Z��хp_��"�u��&�4������
�[&χ�lr�pC$�W>�?p�&"&�;`�B�uۊhvR�P����a�t+�J�})�'_D���h�A������G���7�5k�㩥��N+�O��Y����~6��0�୴�*����߀�BdW��%��p|)�(t�X�Q�>m!����C�Q]$O�˭�(e`QH��j�H[^_�n뮚�0�!,��dCD�>4p��9��s_�'�4Gi��4[�r@��`�ǊHq�Q���	q�M2o��޸�(l�X
~W���5�9G�i��loާR�9���A�J�O�K\�H�> ��{���.�f��aЂ��m��UQc��C`���I��:�j��YO9[:1�'Ys��e���` +ǝj���**N�A��0��'�F� K1�}/�7��D�i���Խ((�t�Χe��`�[w���z�.����z7��V��9c|BN�
?�N����}o^y�J���St��(�ݦ���$�3m�Jll�����9�)m��V����흁q����7�a�mb�ʄ���{��l;=�%i���9vH�Ă�a��4��ŕ��p!��Z:����'ɄJ*�ތ�%5tw�
4Z�?+�4�"���.���_�\�����	r�к�<�h����a��ɹ#��A�e�f�O���Er�{�n9'\� w�W� ê���:��"�W�(2�1�0ݧŹ����qÆ�aZ�F\s���")�G�s�rŋ�>�Nkxܥ���rf��.���)��]��>�aSzc�W�	��sJ)(���=���H6�/�������uu[��Q��*��V��Q�Z� �YO�=����I9���Bz�0?��ݸ�C�ZF�="��]2�ޘ���]����T�Mo#W���Ж'�R���z�U�^oE��-"�C�g�{�ͪJ���hd}�4���P 쟺����7A�N��r^�4�`8:v���snU��(�8�w����%�:Gf�Y�N�,D�p��ӳUcs��P����pK����D���;%��}N*�Y�SّY* 2]0��c���d�bp�|�U/�'$��M$��vmm$��r}������:����Al�4Ј�L�E�Le�O���2
B�`���c��3��q�G���3�����:�݀Qoq��`j1�s3G��+�ư�&��_�0R�B����/����!�4��u��S�@pW8�9u�����v@}��<�<�. )���&@����)�u��V��כֳ ����v\I|f�2i��Ͽ���uY�_��ߕ�%���=�s�����8 �D�d}MH���93�H��ՉpCX];�P;�
T�l8��W"���+8H>+v�C�L��;�7���"�x>��
�Ҁ�"����� 0ݚ��Q�1XU�^��u6+d��C�ӆ8���u�ZI	�I!�0M��C<�Hr�g-�3��&F���xh��I��О9؈y7m{� T��7��rT"4�xh�f]F�g�S�s
�6����D';�w.�����@���*�7���F�3ڊ�+�$�|�Z	E�����3�K9���Z
q��R��C��Ê�!ZX������G~��1/����][�r ���kq���3A)i\)�o.�d����*�Ա%\��;h͒��)̂�L����� !*�*��0�%8~+�m,�>���K�:�vF4\��P}���>[ٲ"�4n���a����@���ز�����'CŬ���'���h\#���vD�N)��{9�'���:c5S���!tA�?P�#)���� j��v�R��ij���>>c_�����+кȢC������z���\��o���օε������G�Ҧ��SOA�[�N����y�hD ������m8_���[9�hѺf��6L��rP��0���S�N-axQ��B��n�b��{��j��}I����ѥ:*T������6��-v�t���mn�+Y���߮MIz$E�����1p2����H"��;�)�wo�[{�r��q���M1�T�N�۞�E�V��`9���[=��\�ق�=^:i�QV��q�1Ӥi%b^���� �~E@���������)CJ'�����D�_z���b��c�'xY���F��ͤ��?��o��U�����޽���g����%_-F��Չ�
2ݟ��S!�;���ǻdG5u��aD��fE|h���̏��'-�������$?d���X�pG��"���'���5���Y�`�Vݬ*�,�}��I�S�HǜMì��-�5 R��P7)p��r�A�w�����e�X$���罭���jŔ^,[V���=uHP��_�s_=Z����:~�D��蠉�`��w�D:��r��� --��l־�OĳY��B�m=ӱ"�٬�X�P���P6`��h7stp]a0i��A"�XrfŦ%���u���_v���U��J�Ϥ5P(�^W�+d5/\�E7(�h!��6L�O��q��"�k�[U�slu�$D�5J�K=��W�>u�B� �M"���������(K4����W�ꖧ�>��p�t�=5g�%�U0S�/�[lf8T���cqn[���x4r.�az+:*��6~N�
`�j8����a4y.���W;�>�����7�����.�>�yVL'P��=�/����?pEmZBw�CB������6�^[7B�2�M��sQ߆ݐ�w����������B���a��10���S��g�`ߐ��:r�_9W���mM�T�����3��=ߏ���P�r�.���  >�r-�x��@⦴����q����R��97`4w6���j��N�f�)�OM�N���%'�?��H�Y8!�;���_�ej�N�Ґ�P	Ȫ� �E�N�KX�����&��Q}4�Cͭ�}��J�/wyW;(N���L�=' Kf�F�Jbnh_b����)��|ݚ�J,l��@I�!�v������mko�j�F�fEAL�Ｃ��DZ����$���<�W��`Řci>�����|Ԇw%�b�$�	�`[h�F��ԇ���^ҙ]{Ү�{�cV[��eQ��w�v	���p0@�`B�)^�9�˛�cP�Аb�����Q=%B���}iǚ��B'�)¬v0ۖ;zk���ڤl�P�Lf��2�[G���u�?m�����^؁�8
���>&������r|��&z���(���l��XAt_�܈B'/=J�F�{6:)$π�)?[|Z���CC����	�� ޫ��\a%XL�#���pV�!B�B}��+���b��rG��h;i��T���FMzd�L�2D��f[�9�*	h�wm�F��}Ȯg�7�޽�6�L6,�a�`�V����a�e��*�12��<+���poF�7خs�3v�ߋ+T~�OA��>J����l�����a,�߲��Z�n�ݧ����l���}�im�n��M����W�s}����5M��W�������!x��G�5{-�)/GO2C�1�`w�$CV���C��䗺�ZfT�LA
��R����8�	��
����YqE���jy�R&���zi��lY+[��G;�/��ˆ`����S��'��D�:�D )�?��i9��
��A!���]��`����UT�<~Ϙo13�ۋ�R5���GA�VA�07|Q�3s��p���m�$l������!�X��rq{V�Պ�}����	W�.�.ß"��.����V��#�\�ʕJ��ʊ���V�*�D�HO�/o��/;���DH��9�/b��I�����H�t��*vބ�Z���$��q`�e0��ۚ
��������*3K��r�CD�G�����V���G��` ?�F�����ؔ��ϫ�l�k7�fqxg�-jOC�������c��"��4ԍ�p��F	����vP@L^%��K���V��<0J�(qAC��N��!{Pn�< �w\.׸��D�R�u�qő��yR&�����z���4J�Y"���$����t_^�٤��1B��Y��&���J:Hb���*�Fw��:����B#�3g��2wG�p:Juu�;�E4�=�̤oȃ�|$ŝE�4m�C��Ք�f�����[I�� &D�mE��%a/�c�<be_3�9msR��4e�*JƯ E���m��mo-/	@Q^�e�/Qs"{Ƀ��m\�����Ӡ���L����������˳�7_�$�A;��v	�5sd��=Շ�?I��č��c	d�b�T����gY��g��
���*��W�਍S�*.�)�ԐU�Çe6 �ܺ�H��,�B�b�	
���V`�\�1˦3(԰�t\������g�A{K�.��)9��"��Z}􏝦��Nތ��n?ً-���Z[�%��Ӹ�	��%�VL���������x�e
]X`[�\Փ��]?��y��>���BJ��J�όC�U��(��?��+�ѳ���s;V̋	'Y�P�&n�M+6L���r���A��$�z��|���~} 
w���4�k�}���#��y��<����:UN���8EP���oZ^ƒ����x)0�iܔhXlPM5L!���UUԟn��Q9{��WQ,Q��o/y�P�����&�Q<]-���h���UZ�����gȐ�<��R:r� �ܰ|��Cvy��b��=��L#���W(�{i�#�&��0u7b�k�{*:�n<{��IN��]c1JuW*!��tW����^���3��-ow�M�恣0���$�m/e���د3�^��@*�?Ӽ�;<b�IjL�.V��:YJ�h�1؜:�s��z��.__����Z�x�H�Nf�K�n�������^���F=t�ʓ�/ӹՒܿ�N�Xi�*V�yg�9��`zOp�����S� (��n�n>.3��U	�u�	LI�#��׻�a�HH `l����2��AȌ���]�S�s������&L�'��~���g%���M�]˵��}-<M���]��y�I7˭ac��F���&��r޷��\�� ��8&ͤ/h�g�MeJ�h�vK|��wa���]�@� Bc��a���o��2��\հ���.|�{m���D�Хx߱t�r���{H&�	h�oý�Z�ȶ�\�B�/C>P���+����]~�s6&��a�x9��b[�X�!�yQs�H�ld�����˗>�KZ$Ņ�ڼx��l ��i��d��b���IQ8ΓЊa�w�ʿe�8��U"]n��	�)�݁������W�I���'[O�G/�#q��B�$Ɛ���6��:����A�X�/I�<��}ʶއ�B�.�����nW'��{��r�r-�����`��Ԗ���E�^9S�HC��'�[y\����pR˽et@r��.�.V��J�H�5�k.���]&�*T�zV�ꔔ�3H�!��c�ŭ��?ʜ�_�A����6����u��cF2�M�����q橞X�bCj��^AHJ�"]/aR]g�ܺԆ(?�[�G�VF]���ݓٮ��k�������(��c�7�5L��e(0�R�m����IX�!F�Y�M�1�Y�ƹV�V���@�+�񂧻=���b*�H��1��d�@m.�_�:K+�k�S�T�e:c!牺
��9�)�h<y���@�9���e�TO�!o�q��я���N�$�"+\����sT��N5J��̣!���N:���	�C �"����v�|���p�,;��G�r��|aV��)�Q	�]\r�"2|#�zUl�r�g��k��L��o��Q&�`~�p@ńp����R̸�W�҂Yx.��5i��0M�K��Ø��ڝ�J��4�����@�p��2e�g�4�'{���淚G���G�0^�y�?I�f~��s/����((�q▭Z�#����'ݗs(qpZ����x��vVr4tm<v
`�Lp3���H��w[~���b�{���&����L{4s��_B�+N�����E�ޓ���������x�ֻs;F�U���/������q��e8�2Q�me8���P��c�*��0��YwɁap�Q��NH<h�/����M��J^6v�3j�[����[*���t�8��!�yB5'�Y��v���Ռ,hÈ�W��@A[X�� ��
M�[��f��؏g���8�����F
��I]��s�V��K�����ǟ(��[�e����/~��_R13�j{��{�:���X&q����{�{�7/l��
*��
��$(��x�s���W�<j,����v�8B^{�u�v�������aR6�0L~��,���}�W��쭉˵-�EL�v�h���E�6m���u���$G�֭C�q�����\���l(B^�{\�p,�ߣP�2Ɋ�E��(�E\~�wC���*�[�|�,1M�V.�
|�fj*���i��/��W�
Ǒ�-�o����]*.��ᓢVn�bN�i0:�b����Sy��x�_�4,�)z��,�t�1oIm���cU*��u�0���A䶕���m�.ɟ�%a��G�V��5��͸8Wf���P϶)��7��,��|�$,*�dm�F�t[�i@uc(����Y���|m�
;ۧ��֞N�|�wG��ߦ.��_H@�Ki��ݝ�-MX�������>Y4��)�7;�mj"ܪ�	.�\W��\4
#.,�Y�d���3��l��@�/�*ˣ]�B�?>D�B!�[p�q���YN Jmn��|�3` ���5@Eс!)P�!�Wn|1k��\�&�{n�?�� ���|Q[���r�b{�;�F�m�A���ڬ�i>󠢤*j�o��0j6�Zh�a\ڬq��o5�Eg�m�O�5���uc7=%A�+��7���D4�guM^e�>K���j�g�Ӫy�0�"��U�z��C��V	�@�*��4(�`��{1�8�Q�3�v�#N��z���z�L��J�&�|!3'Q�ʽ !�G'�a�}�p�N�E�-4���ϧ���E�4����"r���p!;Wk�W�J�Y	X
.'b?���}�w�1���4ݛ��X����;�����ҷ�?��mPXu.^�}E�m��V-@ ��#[����Lv1��>�v���{`g��ހO�R�I��,�{�*�u�WJr�
�i[E���mV�13-ܢ�P���A�z�Uxؔ��v�Cc�����	fbzX��#�����B�6�~������M��q��B�s�w�g;�;��U�+���Բ*pJ'e��u��XLz]��L?U��477�?m�m�"D9�:8ۡ {�RĤ29��S��f��0�G�<��X�l�l�I��(Q�kə�Z�n���j�ZByjnvx�e�1���2�����s�@'ך���5h+	/�T�.|6I��Nm��Q˼�w9��޿e��a,>�	C���l�V�O{�8�I=T <�hJV��u������rG����!�σe�L�?��m%��������3G� 'NNP�;�V5����#t}6�Va7���p;���#BVh!xJ�9��x��7� 9�w���ߪΉ5��"�l2#��ҋA�Z�����|ܺ�%�O��ޓ���WM��:Շ��%\N��Z�N��7�5��׶���=�!�"0��9Ļ͠X��ۿuh��}��PWH�A�k�82s�8���]UzrVG�G:�o�=q�qw��5��k��@�u��$�zl��pˁ^9�P��Q����"������a�� H��%�9Gyr, 2V���4�@�唔�c@�.BUe��I��"S{���wHU�o�� a��E�l�Z�9��$U�~9���9ɰ�o��s�]I����8���1y��N�$n�Z���~�p���k�po鴤�>r��1��n�A��e�A��	;� 4���� ��R�Y�y���cD�R����C!`mi����}�cAi]Gn/���R�X"L�0ݾߖI�H@*Q����S+ӡR���5aw	��ߺ��k�\C+$L���l1`��$�Ī�$W.�<9��Zw$P<4N���px�����$S0�`��4��i�e�Ύvu�T���B��Σ��n��Q�,�[lЏ��T�_�<C�6����3	���`&����k��YR >���K��srOBͿ��{KZ� ǅ� ��_XN��S2b}g.��h�>��f��R�߮Y�pz�T��u�P�\��pN#O5֥����k�7`׋�����N�0�M�(T���.668�����b���M1�i������nL����>7|;�x�����7`ul��t4[y���2���rp씕��,�  ���g���b6-m���Ʌ�J��E��Q�k�����,���Y瞃<Ь����B��c2�КD|P�&R��*<Կ��ޒ�KڄD)N.X�d0������'���C~��簽�ۀ�:��`���H��37��A53Ƨ؉d��4��8o��H�9�Q�	�M!	��f��\�Sκ��y��;��8���p@��}b�7��촁��Ɵ���ع���Dl�v������ (��vm��&���|�1I�#sv\�/��a�x��r���l7���k\;�2>�S�?T�;��N4O�@�k�>E M]jB����)0)X�@�c��'�2-5Pt*V�؃���"����߳�z��8@Um�R���H'H�?�\λ���|��{��6�E)}�HN��Ɗ����;����2�*c�wZ{]�R��=����+�����%ٕ)��c�Γ�4v�(E!������7�'�|qX����@����_������]ѱ�j�4vĠhU���6d�J(�i�Na�(�Y<]��|dC3+y7�V�#�!�/n���-�	s�f
U�'!U���D��;��c&zP���z ���O�\��ĳ�rk��g��J�9��m;tE��h>#���{�p�j!�O84Q�Ĩ�Q���
�<���.��Х�?1�'�30��6Kܻ��ɭ3�1Q5�������.rl�4~��KR���CE�ܘ^U������Q���3	�2L
�'Z,�Խ�FU�-�2�&&�e&��&�)|EO���s`6���d0�"or�})�HH3�ρ����O��k�
���W�M�<<�4)ƾ�B�z��kL|b�j����ȿ0XU�����]Ҁ��Y�lUׯtufh`�<��^�ʼr�GpyE�G�V�;�Be?�'
�^M���Q�e0�esB��Fsh�H����vj��w]���#Fi��a_�	�ɀ�k��
�I�޼bK��;�p+k}g~���:&�{�Yv�i'����2"j��������W�&�߷�qeck=�E��G��ܔv�`4��������w)���H_�X�$���3��ǆ��� -�{'�	7�la�4�t�w�W�+yl[�l�zN���a����>�XH�0�_FI�3b�� �_�c��?��ޙ��t�8�g�Ds7�q�4�9�u�����K'�r��3lz3̳r��8�Ǥ����;)G�3�36[�W�Z�$�����Y��f���U��Lo��sK�߳��E��p\��5P�'u�u��N��B������/�=����F����0CZ����N�|�C-��hu#�+\��|8^��.3�/n��W��.",eҞX�;��Z�C{�q��m�4�������D�sܝ���g1�cb��\�l��)+���0�+�X��Vu k��X@�ݿ�N5��bo�E$���`�&ًf�Y=�'�S�{�]�5�)���s�EfՐ*m�L�Ϡ?����>!������(�)7�3�D'l�Ik�0�!S h���	���QuBl�W��+Me%ɴ'JY9D��_8I����p�_z�&p�#XI�;���IY���Q'�=� *L ��A�7�JFnTi����e5��d��q@ �FgT��@�D�H���'�Ǌ�l���"0B:����� S)/Ѷb;���[�(-�۴0�'��˱(��i�͓A���	���2��r���4o��I�^5{l����\^�{�'�P��zED[W����l��'$�r�I/�u��~�}yO}&�ܳ�km��'��M�r�a~j� �tJ%r���M�i��5�gie��k���4LuY<?��NAOB�h�BK7�c<X�X>�.F��	1SE�tٟi��łS��2l�-E�тK�Iֵu�-��d�Y��@��V��
��g��e��nqm3a��ʸ�v��-O0�.c|��z$b\�e�~|%��HG��g$C�Jz�7�;��2HQ�ڔ�'l�7��aE0V�����Km�!�����z$"w����[�ఐYct�X���ܽ�]3���=�H	����Gs�c�"}��=~��+ZL�_$V H�t�{�0D��?�e�ɲ*���%�Zʕ�HF�[�d���V��8�UP�1��E�#��绤�>B�|��������^���IiL�LS��3�Lb.g�#Jc�ͽ�}�+ؖ�X��&5�G����,y�L_�����W	��=�m���"{^��xH��^�ȵ�G0e7w8��
F ���l�،o3K�ӲoX>t�UC��+5�c��]ɐY��ࡻ�f��K�鋯oĆ/�1-�s/M���?���\_6T�+pH�ԃ34y�8A����Vu�7���T�\���j���-�����W��`p��<�6Qv	��6D�5 ���WĬ�'Ld4ᎍ�1z��|s ��/kg�q|��㠟ѳ�8���y�-�����HF�3���'���f+�����LOB���n5����]X'>��^Q"P9�P�è�(�뱝Wi,co�N���&��ig���6�ܑz���)F����l�q5�v���]���x����&wni��QM�A�:5=���?�B���2G�߀Y\~[U�r��iA�q��x�0%QC�k���#LP��e�cɣw]�s���Ae��<�z�f+�J�;)1��{�M䀹Hͳh{�G�v04���W����)�[�����IU?�-��TZ�D%@�GN/���B;4]-�7ڇO�(m �`�5�r���@Z7G�Қj��l9.��������a0h�5�����2���+h࢓�JC{�* ��X�s+��/r�W��]�<F�o�w��z �m@����G�Hڗ�u��i�n��z���B5�4'F����mҕ�������)�+�j{�����B{z�aۺ��¡����R� ɹ��H� Eu�\ز�OG�tM�8��"��rNģ��"V"��j����ي���>��M":�G�l�KAU}��}(|���r�}N�6u0z����w:�n���~��}�#�EK�~��d��29(��_pZ�r����F�r�1��=O\@
0X����� �N��;R�yc��m(��������sMU���X�U�KAE���E��VG)�u	����$�Q���:�M���OH�A�^���rR q�.����!�vn��!���;��D���ç@�+��q��]�܂���[��AϠ��C����>�ߡf3ha�ww�@S��� (S��:|V�̇�d��R��e�?H+aۆ��m/����*y^�8��?z7;��0`�tf���|���fק� 5XW�+)��RA�XA�6��m��lQX�gwjU02���ʞ���;{�{2ʱ��γ��<	��C@�	�~������3rq��۩N��������������k}����w��|1���^M�(��a/���Ȕ-��h��y�@�����*rY�mA>n�}B��0��o�m�Y��9J-�i�Ťk��Sj�X����ԕ�<�����R�h�����)47D�Ǹ\�u��s�����!�F��z�O&�JI��|)Xd'6'f����l�s��̦p�0ĵ<�%:����<9���`��\F&nb��Y��}K`
�o&��*T��M��S6�|�#�)34������%IFj"�^�I�`�e:�\OF��� �m���d��lz�sA�+�F��`�x34�|�)��$�YgI�[�d�mk�ն��t-	�Vqll��d^�8�,��ש����9�P�S��S�-��귟
������s^�>�L�I��dli,O7>��<V����L��V�.����)[�F7Ѡ�7��a�%�B���
5d�����u��R�Ͽ��������_<�U��r�RU��"+������,&H�۸���4F����(s�\�ګ;9	�\���::�Rٛ\nHlD��p Y�5�Qa�ϋ�������I�ٿ/3{�':�4��z��=�c�pϊ�tܯ���7.:�Y����QL[�޳+����}�]��p_�T�%�6#M�GyV_�:� R��9zz��;�����.j�x��jשEԸAԟ�0���B�!�҂8�� �D��(u��&i���L�ٸ򉰘7\a�v���B��B�5n%֮	���1�Nˤ�	^ƽ��t�ӌ��W߀+��n1A��"��f��H��k���U�m�-�,��|�XN��
 �FT�c�� W0�� ���i�6֮+HJ�E��_��ғW�oG�#�/�:��%��狤zB5PkSB�ͭ���˥��J�<�*�ؤe�hA���T'H���0��C"\n��2����\h�KB1�R�7}�G�$WdO�P#t��WA>g��#e� �.J�=c�������!@���A��/���M�w���I�#�8�E�ڿt�c���A/&�2����#�G�4��^�h�c؄k�C��;mq6�}���@�9��������DI��}y�6����	!|b������	�:���>�
e�d�Xޙi9A���o�^3�P�x��%*�l����q���d��l���YT�s� K!:��;M�i��hI���z�bvL��<S4-/�C>��q���<dP��,��$�N�Z�F����Έ���!�0xezʱ��o�j���&���h��<\����b�z�:�I�7��ӧ���N)/��ӄW�j�K�UgJ�U��>	C6�����+R��d#KTQ�6@�K+o���C�a!8�j���Ī��1�%��B��� &�-k�' �I NUw��-W�ZĦL@�?�๳�����С��]��f��6�N�!ÇyŕY��C��=$��[�NT�1����8sSR/\�~Ѫ�њ	�$�j���������KY]���x��ɷ:�E�z�v`/��|�L5#� �p�N��k�q1�*�Dw�����	���5�I�q} �8Uxn��͔���H��X?&zo���s���-����O.oX��[�1T3�����lU���ߧp�H�]>6v(x(��K��<�L:k.�z �}aL_�a�nn9�� �?��si�?ٮ�Z��Z�l�%)��`��6R�.;@�nm,�*Q{��-E�";� ��V��$	.��}|�:l��"�>\�������r�6s�ߚ���o5�
z,u��6�m����G&ӫ�5O(g�׶=�8���ܢ�<�>Aܕ!�Q�o��.p���[a�<ᷤ��_�,��+�TV���]]WI4 ���֩�=N��0]Oy��bww�>�?9z�Hci��e肱�gl��ݡ��B�c�tҀ�l�ı��!z����EI��n
��PQm}d_��9�E�>�C��W�b��e���WFoI���33.W�Lؓ�)�Iq�"�����1�k�(	�9�iZ�=���� p���u���>bj�n����!����%RZ��&�`�:��%���nT8"�Cw��ٰ�r�6}�,�ϴ�ts�S귴v�Ҟ|0���o�B���N'Nc�2@*(*S�0l��"՛�L63���`n��_ԘST1ֳ��"�Ņ\����zoU�$��_%��9_���{��ԋ�^���7�R�$�叞dN�m4>>��!�z��3K��Ajܫ�έC�1�'c�Ʉ$]���R!w?[�e�� !�HZ�n��.�CW*jf�3	��KV�$�찳�h��"M Q`��U�n[�	FjH�~��GG� ��BL�� �q��d4c@/��kT.:Ejܿ�^r��'2����5��A:)���uu�`@-$�H�Y�	���Ib�U��gĩ�`
��laHq6�ֆ��E/��r��ʴ�?n�/��啲�1�B�1�J�Ω��Z�;�뽔�ŉ��:�㒈?u��"�'hi����E4VP�J��b�ܙ��WdZ`�4F�.Q��]�-,�;�T%Mr�>��f]n�V����C7��NV�@�/�5�a3�r
iTX5���(!�x�7�.�b��Um ���xe�������Mh�˯k{�A�Ó%����!H	R?���o��mLF��?��#�m
_1�4�w��X�~X|
�8�}�����|�^̈́�%�2,��h;�܄: .. ��L����N8��!i:l��Л_m�\Ha��x��֑80-}P�	�v+6�^�0�D�eXb$J��d�v���.�o��:��nwK��l�������)�IF�s���M�vV#��������sH�� l�:ǋ";�
)W�
��� h�����/b�ʳ�H�ٿtO�c�������Y������t�/H��a�	��w���k~�� ����b���[/�_�#���\tC]3�0#n�o0����/�DZb%��m��h'�����}�J���k�\�,CY��@���{]���݆	`��BpMb��o��=8�/B�/�C��yHJK�=�;ה����/�_��ɺ��F�,���ʯ�Xs3n:��bk�z�Sn�Wȇz�혒aL� �j��m�#��g�˧S�@�%��'�n'!���X(>1sMm-� B ��]�t�P���O}ع�S�/3��rq��a%r��䪿?V�@ΰ�ǐ��,8&���/ƞ��`�6�)!����P�����p�u��ߙ�;� v�mj�p��J<��M����x��ވ��j͔h,�b�l}_�ںf�1��Wz����dY� z%��k�R�s�RQ��G�w۬������t(e�@EVFw[4���ʸ���t+@��t	G�����I�(9?߮�E��� ��xyQT��t�D&{����KhB:��9q���3��c3mc���y(N��"��D�ϸ-�4�d2(�7 ���T��l�#o2#�C#��"B���9��y ���;&p�h����*t����>^7X��L��Cx(��=�u��A����R!8�<�~f��V{�m�DM���Ʀ��F��0�eYDoz~	=��Bӂ:y-��#	kGS��#k��u^�>�hs�/����vh����..w+�Z���~K���.Ź�u '�A/�kK��L˺��(��Ĭ�[2d;��uQ-�C�񖎤[kRK�3��>֣#	���b����� ӈ޻�������^�Ԇ^�JÞ>H�E��`�0^�0v�t���a)h��X�J���DgQ��,r�)���B�����U�9𤽝�T����%����6�l�\D۷��
�;V�):r�sٿO��N���+^g�Gl9$U�^��o�/{V���c�~��몭�9/˧&+���ݟ��������o`��-q�Ҝb
.����a��D���Lݡ	��(q�g[a����ꆆ�[�*rE�U6�������;!tJ:�*xj.��.@rm��?�B78νsyh�z���߶�WAT�0Ld�M�P�Tu�Pe3�ӿl�_�	��j�u�\{�PI �]�FI� /n!C�n��]*��:z��H��:g�����x�8��$�W=xP��1��l�m�DD�m �݋3����e�oT�?P�V�#_<���^{�g�#���_��C'��Bo�A7�D9&�Ռ!r������Jp�����sr�ܯ�dg59���M�];>V�9��LF ����@�~�_� \� ~�ȠJ=����M�T5�B*��+�=��
��C�ӌ�:��Dk���,�0���*C��'�c�D��&���-�o�`6p^��l��<m��F�)
`f��n���-5֙����T(��A�6+�R<E�ď��R�9Q� �uuu�Ln��/� �Q��B�s,g;m�in���#�Y��#�=K&�/�B)��:�fL�.Rmqbl`�_/��l,-`2����==B*A56׎u�6$�{�!�cr��P��w�D9(����Q�Ƃi�rK9��<U��A"�Rd�#�u��֢�e.��_���!�U�*����$J�(
�a�f�"\�*������R��4�ѿ+\Ԣ��[��Aމ�K�k���A���?�dp�>YXp��ٓzA""��%s�y-K�0���c( |/�*<��I����2ս��'����9鿀�i��G�U��edF��|F~��l��>�&f����f�[%��(��5'��N$���c��wq+:�xG�Z�m��`��'�TL�:t�:P"u����7���,�n#�q;Q ��q!��&��%%ot�S��F������|�yꙦ��Jm|υ�`ϕ!����"R(�k�� S�g�3%%�>sw����f��U�^I�,�U�� >��P��Q`�VgL�Y������-�+x��C�/��aAJ����T/G;��l>f��UM1�����w�M�2sz�o��@.N�J8,@V���a�N'��P"��l�k �\�A;H�d�`�?�u��!~�������X���砙�>����C%kP�Ŕ7���`�
�K�a�A~�=�?[��K��ϟ��	$+;����܊V��������� �"��P�E��.Ӓ`Gd�Q����q݅�I��نZ��a���ܭ\��r?�����L�N��J=�;���%Tx.QK�,8y��hB|t1�gj*��]_ڒq�Lc]ج	���Уy�fԛ;�|��*���l�M���KX�Ob���^�(gm�
�K���M�f]$�6pݴ��
òM�Z�ce�z�<y�"e.�p4�α@"lM`ǟ�Gcq��\�O>��ϋsҝ�t�̍���ɨ��:BRR�̵�1_nX3�XE�+���~B��'�&�3���p6���ZJ���K9�J;!T��r�t$���$�$�ymu1�]�Z�n���c����VT8��G܈VB���������k3��Uԇ����*HO����`y�p��������M�n�B��M������8��(ʭ���p��}ug�"����}$�������R�E���kD �2�nX ��_Dҁ���J��";x��;�1���
����.e�� /�d�!n��")��9�"��;�c#g���Ջl�uF�jz��B�H�����:%�-�M9���6�g�V ���@�q�(o��v�^�뱫�ڹ��x�8:J�-y�{o��I"�@V+i���+���Xb= k��Ίu�Su_�Q5��S|��|����,D��B�w���yUcʻVC�|���4e���긧1#�]�ѥ��ň۽|�|yHi8��M�	`�zń�ogɑ1/���.�G�y}�.<7E���������Q�Z�D	Q�5/=�^f%���Cѻ�����뼉*�����]b�-�=������0�]Ѽ�il���S���Ԇ껵{���7G�53> 
�*�;[/ޟ��#�h�"���C]�aPgKP�ī��_�{���!�PڊwQ�l�	�zU�S&͒3����}
���N|�L�3f���" ���5�|��5��@�LY�X������j�cF/�h�:�WV������O߷���B�\�e�K��I����%Լ��Ն���m̀$w��An��a&s� 15M��g��[sնv�O���
8b�|	�hk�K�Ln6�)ڳ�k��V8�Q���V �~���$�n����j��O�.����β:xl|�����]μ+��l����uJ8�(iz� �z��}P<56yt���4�=�޷T�1���py9�q�@��T��ێN���3�3�F^�Xh{0��j�=�2���W/c�{l��-� "�@t:����nρ�F \�o�t��z
�h�� �=�~��pF��"��mO�KgR�F	a!�sb���sMk���)F�2�7&/��OC�Y���X����>�us[�����kOy��uk��������Z���V
/D��=I�@'��9���]�R�VdźC���]I�i�q��YFEƂD6ab�:dc��owR=G
3Cx�a`>\�Alz/�U|�ԋ�o�!$�XW�zԱG�V�ҍJ:cn��@Ǣ�Q��se&��c���������]����_�/�Õ<��}���A4�������HxHK�����s���G�зiT>�Ӧųbӡ'�N��K1��M��Tɑ&cT\��\��Ф>������֕1�=�u�ϼ�gF�jo���t?���{��wps���gw�����t�&G�=0Zf��ܶV�s:=�)����{��@~�@dA�H��mL�4��͉��:]�����փ�X����i+(.8�3��* ��}Z ^�>h�	e�kTV�X�0_�*9͛e����GZ���R��9b�@�`Md�����v&��~����n�?jC'Z<�������뭣�f���ǺyQ���!�1@�M�V�01o(#����#�nRm��0���p�RCc�_�K��a�~(���0%�!��݉��.p�W��rC��e*b�V�<����W��~c,����Ъ��s��� M�U>�ׂ�ƥ����f��w�;�r{���-�X 2���DPV��3-�F{80�g�57$q:(��3�x��x��[�Ik��W��j��0����9�mf��<�_3��w��ϟ�_�b��4�����`�k�?_m�^�Q��J6���F�C��� �� �O��p"�p��"y	� ��n�gj2��`8w��;�!�@���ɍyd�������ԑ��F�k�[��w>K�-����7x��h��'H�'�ݧ�aץ�F|���w�0E�3��x�����6�������3��w��l�y2�ѓ4����au�N��nJ�%��/���:U��Zi�V+����[�74M݆z�b�b/�<k}�33Rf����"���^w��0�uZVV(z�nFBm��cwy��e���u*���EXH�D�Xt]a���z�%�En� ~w��}�ԋaiC6E�9X�D9d_���d	F�	l��b��l0�q�n�Z�	b�o^��b�?4(Rcx%��!�MؕtĚP�s��̇rm�W,���?�0�r|Uk[�+��$��I�D���YH"������y���G?��4���(�#7F��il���U��f�Ѐ�F""@Rm�>��xB������+o�Asu`�b�����A`ʆ��^���ۛ���˭�ט��G+}�Ə��լ��+�'����X\1m��?�\O��i�q�)oD�J~y��|�F������2�^�!{�+?57!l���Yg���� ��!\:�U��Ly�F�ҺW�b�R��B.�S��s6���#�������_�b�r-��5W�p�(a߇@�r[��챙���Yy�ҝ"�IO�K�15���~�QҪ������N?2BCm�����T��m��n��{�a�K���b�x\�\?�]*V�l6�8�)��A�2�!�7?�'C3��#N�\L�vЦ>�Jdۚ��E���ʍ�QS���Q�u:T���KHoղ-s�c}�w�xe�1
fvC�,����O�F�)U��yϵ]&��cWE~�m(o�z���_W��SG�eӰ�7���M	ř5�y��{��2<JCJ�6�?�ּV���ʛ���ѭ�nU�s����)�&����l���| ��Eo�X��+#ձt��*J�o��jP��}'ͅ���}�5��!�Q��m��y���{���5�Z�J���.�ٶ�rC�l�T�w>����o6G�C��T���_�z�=J���Ys��6X�6�b��%H�B���H�|���h�������$�vj�I/��r`���q���|��K��q��e>�	���Ȳ������6��#���Md�'ז%t��aE-	�i��-;����pr��� ��Y�X���g6ᫌ�C"���B���?�t����$
he�\�>=����h���l��܈�cF��G�M��,�Ė0`��v|VM����w�x7���g�ž�����o��i�oٕFG����� ��"(�$Ҙd�VS>5_c�"j �����~�?RrD6׸D�)T�5Z�2��|��8X7�Y������Z�lx�㘢{\�7L�ɷ��e����t�: ��O����J�7%�P�7����h�h���[d+�l�VL���3��	;@uT��1э������k܍��~�yK�m������-2ׂ�Dg�[�7�?�Ԃ�x����0���)"�|���oY�p�~[C�u�Ɍ�c����>w���ͮ8�(�C�@[�(&�3|Ӑ�Eu��l��N����H�����B|"ݮN8�� N�;�A`��+�ť�6i���.=��YGt)7S���.���kp��e�]s��Iʆ�d�RӽE��U�UdG�$�F��f<0���oj��$T�|ML��e���7;�D�N9�S��ք��(Q5�Ц�߬�{��Ob�G���e&�fz.nUY�Z]�T�*)S]ZD�t�*�Y�%l��B-�cb��AtBX�Q$S	�/�}���SD��29.��E�<�k��D@
\�|HZ5a���� �� e3eOO�`���j�׋��!g���%�;z̽���[FJ�ߔ2��"!����Pz����Uĭ��㨳�g�i�ϡ�d�����������q����k��CG��üM�
�u��a�̔�.B���HC$ix�襕���$V��#�>��OA��ȱ�s���L��Z�_�;��j�Y k�ʷ���'�x�k�M��6P�S�7�G76���R"[-!��g�9��;#��ˢ0'��R� �	�QTB�V����cQ����vA��B��'y��Ƿ�P�7����__YF��<�[[��c)�Ñ���b"%W�x��E�Rd��C:�]##�q1��N�IUrFkO���NF�z3��Hx��T�2���A���	P���X<���3_9��/��R}��L���s6�-6Es�y�?�V��T7KU�hO�|J�UJC�iy�/<����(U^�~��T�s��5�-b9lڄ�݂�K��������L�3��^F�	gER��U}�;|2���hL
[e�FrS#_�jǾ�L��� �x"OB���~�-jmy�_�,�ٰ������z� �;(�<���
s<�i&�W��l�'�!^ '�����1�\[�K����WQ#��K?��L4t�����SI�s)߁Η���-5�w�����c���H�a1؂�QFgy�dC��W��ý'�I���|�M=j�_���j���$�?����zė����$H��5.��G�T�M�cI�Fs6H�WjR<�ө �?�7Z���ж��
o
�D���~�4�o���0m�Q�}��$���TFx�G�W�K6)9�I��*�l��!E��L_E���Y���vd�p�8EL���ګق`��5``5�_.�Ӹw�C:z�`f
����sB�aX�/Wx��<b'3��	u�`P�!�3�s�33�2n��*�oVȸ�!���,QC��<D���23��C�A��#��,(	��ε=$B����5�v�36����ܪhO��6�~L>0.~O`�%��5�Pu�\�/��XW�O��ءcC%u��9-B�U�^a��L�G�Gϻ����]����+ǔ�:���<�d���!ѐ�����DܾG�]t��|2`�p{ZQ ��}8����}����]�{Tr�������h߼�<�@�\}�c���g]�fm�^��Vv-}��K������,��{Ӣ�:��gܼ�`{tډH��N�@�`�f���L�k4�6�cl8Sl����ѱ�\���J���E��6^<��wfV�<����� ����嚡��2��4^`d�
2�AA�߭'�N�x���撥$Z���Sa&���Ю*�De���R�L?ǠE_J�!8���$1�t���F�d~�,����t�v�!m�u|Ax��%�|���??^-��P��%vF5k(�}��SUF-T�I�e�TT���@���uͥ�Q$��f�2���v�A����}��^y �M?�+
���R��6���j�����i��Y�7/Ρ,����_��5l�)�HS|4��U:����B�8�:,�II'�������ֳ��DS��Y=���x��B{�lf1���������l�/f�!�:27���)o�C}����/=S��*�����5r)h���J	����<���M�@����P��1�!#�h3���h�_�&눙|x��1�,\��z�w�d醣W>2;2F7�Dކ�+(y�,�ꅪ	snP�^�����ƹ<9X�ͮ�UF�R�"�A/uҏm	��ct��2�EAt����)?'ƾ�������'A^��7�*5�{=2�`<	}O�����@rm��p����]yh&�ژ��Li�o
[�֮d�����+�O����cH�&������R>��Ԥ'�>$����/y3�~t�"BM�����T'���{zN)��Oϑ���W�uX��E�K:7�$����������T�"�z�i�%9X��o�ԧ�H������ 2X
�������?�o���|���4�U�)��S���&�:Vg�3c�M�^t� ;�Ð�g9#%�Y[��{��]�x�����<C���>���� � T�m�<@S�r ࣍=���pt����_Jr�8u,G|/@t:XXO��A<~�ކ�?	ʲ��ˀ���q�t��&"�Fs䰂F!��j��3�b��>��g��?�a���������v�?E��5 }rP~c�v�/x��k�����!�Y�%�!�t?t����f����ȴU��X��Z���6ib����~�p����W��0����d��ݨ�j�V���Qzi�x�/�&kG�����/�4��1w��M9}�ٷỤ�`��³��T���dT�H�\i�/�1�S�>���p^���\�l��k����w<с2=�<��nmp��lH��
���Y�V]��FM��6T~랹C_��`Q��8�z���N�Kp��q<����PcS���<���H�\�Y���O&I/,��Bj2��}%��;�I+��T��ilf��k&��@	�XO ����%�\h���o��h�����'���?W���K���8٧ȅK�M{�,��x�KX���"+-�{���h~�gN}8 ��VxY�y�ӌ�=��>D������}iLD]f)&vd�aK���>UX��Au��I�V�'��O�6�0�*(������M������D�w����g������^���}��1t��������$f�W�VɟH6|�~��ӫ4ߞ�R��T�aĆ�o��c�n��h;_��n{�#R��:��$F�a��Y�9T���� %�Ձ��/��0e+��f�e����2[tQ�� �`|��fy����wj���:����=
��qiS����g�e��,�@J�U���lovCȬ|�7�ڶW�.��O�U0��Zs��t[B^՞�V193��|['�?�E"�|ʮY���s�n�4��i����a?�p���Xj}ݟ�=^�N'�6a�����Ne;�E0�T��(>L^�~#��s���\�tPs¶��9مı3@�O�]R��I��U��h�Vg�8DP�3�6j�]ֈ���1�p�s��At!3�1�֦+^�X�]��&��H�h��!jf��=(I-5X��p/����5���ߤ4'o��xn�⳪�N|?�Vט��E ��"��*{�|���CRuuo��x��?3��cZrl�W7�Z����5�\s ��ɲ��|��*��x��<"lpL�_f:�?����{�4N�-�˄¥AH��b�+�����C���6}Ƹ�K6����*���A�|�����屐��'�C���x<���i�..`}�S�%c8�s����l #���l
��������:��@��Y�x��6�L�Տ���n2Ǫ%4���A�y��kb����kp�U�۪�V�� O�-]#������ҷ�����-�mQ�
ˆ�6���c)[�C�5�g���K����4E����.�����c�,��&dA��l�y��4-�ˌ.1_�4Ѵ�A��uȂ�Ϫ��/�9���̛�ޡn���"! MU����Q���"J�q�d�Cd�; 17��{%��k7��p$�h��A�zrL��"
%S�-#	�`/�ݙ���rmx)n�}8[5o�Β�e
�ԩpp%S�X%���\y� �%��K�):*g����P2��B4l0�X9��b��[oyZ����k�걐��P_���B��2�2�\NG.�(hK�=����_������Z���=CJ .|�s���["�w��x;��,y�#�P��A�Z*Y�(�>��sW�\��n�4�#p�`�u������*��J 1�ɪb�+�}#e�� _"	�l��{����-�ufh�"�\����;�b5rZ��ْ��إ73�D)L����"�e�!�߀��[�5B�QZ}�w4�����r?Y�̈́���tl�Ù������&��uL
.2��%!��3�k����<�,�?�X,�����􃱀#&�>��@�<=�"Z6���.�O��ߋ4���R������N+���)��;8�4%�e��P�6�������.܍�����7p}Df	���A1�����j�1�Pj{�q���h�Q�8�k�ǌ��I��6��&�zG!x��Gѯ<r. E�/qd�f��F�y��ݽ�h-�W� )�>/6�.(���ڻ��wۡ��<�r2�@��w���8��nG4�t��\����(��i�%��Ap�|�d(-0@�<�s���u�k�&���'z�r����/��㹙���7�l~���׏76�^A|����㴎�-�C����uFh�&?Y�R�e���Ȉ��'ޫ�Kj���d�s����i"�w�Ivy��	���OCk���+�FvgѺ�����9yt��Q�V�M���Z�7s��ܸ��6Q���{�����ۺ�g�f<'N�<�_��d$b+�w�57���y���؛|{վU�J����C�[��Б�$��.{])!tt�E.�\���	��w�g�g#�~.80�����ݮ5_���{*,(�}e�(��9P�2�VZ��+$[#�[1w�ewn���U�?��-�$�֑���da�>��^�;Ku�W���K�M�]6b���o�Y����~�vE��w�\���C>�SX��1]��)y��u��&("��`��nV�);�D���;˻�,B.�&���R|9"���{�s�9���;dI��#b}�Oc#����!<�'ΫU�l���MӢb�%w�pb�V��i���>�.��+5����ɫG�*ŀM��[waF�ç�z)�q�e�c��>��L`�EmT�q���uOU��)�<�av^���ml�U�.,����e�z��a��<�>��n7Z-T�A&R��5��(���	r��SIŐ�Ƌ~*_�GIO �7@N����:�`�	�_���w�2҅~@��)���Ȧ�%�.^=D}J0�yT�>����4V\ª@���ك�y\4�]Y���6E�l��d�/�&�7�,�Y�6g��Y��S�(�[�B::��+�<���LI�I���w{���1DӖu��i͌L���>nNQ���2z9�C+&�K�];zP���h3!X�򰃩I�,Ɵy��b2�&�"��BgK�[��0�jJ;��~pXC��|0&N1)���vL��; 4[ȆM�7	W��(!���+k(H2��`��k��2ј��(L�C�kQ�J�&�C�lJ�3/�^��u��k��|]�VS�lN�
o-kgUJ��D�w��: ���E�.�#���y�+&�~�3'�qɤ��/���z��I�NB�N]V�/Dm5���M�xf�v�Dr���偕Z�T]��/����(G���xS��ӌ;z4��e�5
�*R�8�3��Pxf�@#��ڲh#��%�k�*�\X�R$5WC����R1b�]75�;�Q�����nb#� <Id�AEsU�t���Xą�N���!�Ip �	�1m�7x[r��.c�-�qb>#��ZJ�V�Zm��P���$��a�9��&����aj���vL떧d萜�Ǝ�7H�9�ׂ?}c43]W���~C�|���*��\�$�N���{�U)�R՟'I<:Y%@�reʣX=����D�G�X,g��Y�-�h4�a�|l�� Rz"�EV�K�B���jJ��Q/��y����j)��8�Jr��>$���"�4��q='j�?V�cvb=�o�_C�Uy%�J�Ί��w>��Iq�ݠ(�\KlC1�&�8�<,$R�e/C���NT;3�9�em��.�������VV�z6�e����]B։ɔŷ�U@��u�n�]�*����˫�R�re�]t�bɊKG�oW����Ϡw
���ڠ}7u�\�pR�r$�B�뾿a�:q.\|2Jv�K�s�RuT���v�J�r&D�#YE����%�����$�2�b-������&y��k峂ݏ-C!��(�N�D���"|�Tߊ���}�f9z�WxZRטEh��8��t>N��o��B�!���ٓI�9�̝��;���ӟ�xSc9���p���������N��jթ]�#�nk���+߇ɢ�A��p������{��yˣ.�9|��tg#O�̯k�_�6��|����b��6R.h:-�!,]�%
���*L��=T�]��i��M�B�o�n�����0=.��V�O����mUt����w�� ��N��tC{���Z����n�0�Kz�����<9H���nĩ�xj?�_C��eR�,aH�Wd�Ur/���kp�����BVĲ>�í���d�$�O;��j�O:�u��<L]��p={���7"_4Ƽ�?Z�!/\3�P���}���.ڽ +R!p�&�J����}�NsHn�?�q��v	�%�ewR��'�X��:S���`!3&��Af���v�� ��	��׽�UF����k�,������+0ƅ�����]8Ɛ[�M��r��>S<����Aq�\��@!�X~��oZ���<���ݸlۛ�z����/���1_���v������ߜ�|/�LBE���)}!:�H,�ߏ��k���`����gq�*$T�ϐG&8��g�߀q�k�U�l��\�Ep���Q��;T5Oa��s��4��C�"�* #燐�~�����BV�zoi����ju�B�Y=�����Q��@"w�x�g<൒�JN���%S�ؒ�,
�=HAT���]
�N���m�n����zT� ����^��(R�K6�j�`.� 8���ƪ(�JA���� �x�7tP�"�`(����hs���]���~�<�|;�M>���c@���)( ���ԡ����gļ�L��Uϙ�<��
O9>/��bL�;We�\�f���s��p�&�w!'��jzk���v�Hq)��t_Ŧ��t�k�ߒg�хP�A�k�1̽��a�t����9���Ǣɚ���Z����?�]���ek�s��3�?]�\����$��"�ׇ2(��w,�=�ܱK�����;�	��j�2|��F��f|� ���Na���|�� ��ݐ���y1���v���!�-!͕8B���ݻ����&�"cg~\�}���i����Z��EQ:a�lD�-סl7�?H���ng;��:�q ��_ѹ��~��I�sz)�u�7�u�^Y"�Xx��F�ɩ�%ᔥ.��[6�2�������|�F�C�x�˝[^���	jI��'+�!�!����VTT%h�[�\����\���b}%��A@�z��*����'�a^�����'�$@<�4��g�w��o��L�6*��a�rj�������n� ��[YU7��;!��-~�3��j����q �����>)�st���)|�b>W��wU��D����@�t�ي.Ť�h���k���_�VmT�d��l.�6B[> w�9{�{��j�+{�'M̯�����n�09~p�K���=)I�� \�t��fQI��jzC;M�Dï���|������� ��s��7L�H�+,��a�$� ؅���lE�&7�~Z6i�k{�3^��[IO�g�n=��&t8�A��2�.S��!#S"ruYD	Y�8էL�\׿O��>	����N{��p�]�����9h�\D��5k��Xک�£�c!V���ZFbw3��oi��1]g)B��®�U���̷l`��Mmtذ���}-���-���Æ��!�
0�m�!ٹ� ���-~��I~L:��v��=�Kb6���-��徥�K����g������N�	ڥg�3���ܱ��<�퐘�#�� �Y�Vٰ�&�_�������	�֦?�׆Yyy�%�]o�jfSv����`�BQcE�j�K-��av��.�<�� �BS�'L�\�3��ǯ�[w�'�Y���׼������`��tc+Ի���?ŷ2�M"�м�5 %D�km�u}�K��bq�L�^��!,ܰ`����8.?�Lnf^��uɣ&���#T�փ�C�nu^�E+L>]������dZy�vmZ4����VΆN�;&���]��;��SM�X|��$����M�"P���Ii�4�=p�d�t���S[ix�5(�E^��|�}���[aO}c����*R!Iw�U�GY \=�D���(��WǗ�|���+`�����X�P_�N�P�I����{��yk��i/�c�S�anQŒI�GZk �?ґ\'F-��,�@F�93�'��-���h@�X��̦A�ZMS�B'�e�<�+�?o�R�e��z@(R\O��&0��� 9���a���s!� ��HF�ڍ���]�K�����Յ���4�Q��'4��������n���a��'VVm��R�vD����~�P���;�!�D	ic���d��{�6�x�+���}���I�������[�p;��1f�������d�ʼ��ۈ�ZO�"�����n�G�6:w>=�	%�Gp�Λ����Ɩg�Ϟ4M�1��Y���i�^����`����[u����z*	�ùQR��9�oL�?��!�Pm��N��
%P�6�"�01�S@�\�Nᱡ���\W��.�w��Q���T���Y� �
U��#��l]rfK���Ӄ?�%HSO�i�?\%�}oP^&� 1!_f�ƊF���}�AXo͊#f^��7y�;���n�2��GOJ��&�"oYE{!�p#?xu�}���p���tW!�r[����֥��%q{/�=Gf��C�tv�,Ţ�zr���kc��l��	ZHRm�����i�����ՙ<�0g�	_�=(`Nc7bAV�9�'yN���*S�-�	�fl� FƸ��������-#�dn�qRok��]i���0g�x�Y�6W�� 0����0'
"L�xD9�_��߾��[:3U�T���B\ ��%�_�p~�X��z���M�o+����kG+|_!l5�����$�]���=פ�k��͉���#ܙdN�?�).�BX�%����O�ةb�<�}�)�rK�����|��	!?,x&� �!8zA�J}�ȎиX=ɱP~��q%��iV�,p��1��0ٿTW5h��"��N*�m��x�A!�%�*&C�I:U*:\�-zaG�	8�<�`��6ɗ,_��F<a�1/L�Z�?��4z����6M�K���00Ki�c��ۯ5
]��ȧT8|�n�҆āf�,#΂���-��tVs�#e��H;O��tMb�s�K��N����؊���/X<&1I�1#�k���p��"��>�9}�΂�bv��Q�,�T:\��$�b"ʦ�� ߨ���*6$s�( ���,��ʮ��[eIOY��с[z�XJ��e���oMv�E�"�������j.�f�,��n���ޡ��,�b�CN܈f6��Ű|␲�0�qhe16S%���;7���H)���޿]c9�Rr�2�h;U	�r���������,�4'��]�|�K�p�H�n�G�`� �:<6�}��N�������euE�Gg����!�R�aw:l9x��{N��?��z�E�n��xbv��-$R~��d�7�O��v������(T���
"��=� �C֭c��w�7}�C	���+�0��L�*�djx�.UD�oN�`*�6V�0J.�,�A�u�Pݞx� T�ƿܵ�I5w������v�vǾ�0, 2�[E�K"b{��nq��R��u8�gGE�)r��g��B��Բ=?�Q�W?5Z�aR��w��P�|��Ft�33r�2"�>���`+���	8�i��JI��2e�Z����"ьpj��*�JNjy��;�u),n]�dI@9�Nr�}�#r��4����\�Z�W�P��)�#�˺�]e,����y_8���̗}@��<Y��+WQ_1(�u��c.--�q/)�B7 [�~2�q��OU����dhJ�5�����X�c]��n��
%A0E2�"�,JR��EM�ݵa���_B$�M����������F�&/�N��4�x]b��c��} @ɿm3/i���{|��zYcw7��[�f����U�Uo����+D�hJ���iteM(�`����d��;�Ҡ�erk@�t��3�&Z:gl���݈�����Mb��r��e��(я�WQ����l���ǎG�ʌ��>Օj:4�r��S�Ê��i��-���a�0"2�H����r�ɷ����'eΨ��l�b�bA�a���U�����ښ�cL�$2rD>Є|#+��!/��gdU�U��Y�)��3Q�]�߾b�fTN�whx���\G c�x#��3}��|_[���#TbJ��x�l����Tb�>=�
�`�v^�%� �@z�8��l�7j���h�ɫ����T<�1�����@�b���v�C�٧0{�T�����$�a"ݖ�@ ���ctu��x=Bp�����h;��Mɯ9�� ������X�K�lMk\�鐕�0�<"�w�^퇋b�9�I�:`폼��>����h���]�k/��Ъw�ꏞyD�.���#@Y0��h��c9-����{�ѽ`D��y�.���2��tG��n�\$'��m��W�����f3�%�=\�Ώ���9T�f�h�$��@m������3�l$����K7��R0�Q�m�pԟCK���'����`9/��g:��p܊�ʕ:�TEA���O��b��I��mt����,��am��:8|oiK�X\߳�!����21\<+��|vӁ�9����Śn�"!R�@
i���х�g�����"�1C�V �E�ƈ/���C���ѽB� �M�ً�j�I0O����Z=/0�V����u���5�.�0�/z��Jx�`�K���ا��b��j!�،���Y^z,�$է�����a�)����j㖥���1[B�P�n#���Iw
?��Z�8�S/]�2$�d �� ��|quA���>9'o� �V<�n��*��F��<�_ށ�yKP�ˌ�$6ĖcɲXy����/U���4VJ���*��}G��D�����x�>�63-�G�J�;5�n� ���zI��$���>�Hz�$9`{�(//4p��$���BN����ۀ8_I{�'bm���1G�0�[e$�R�uRZ�Q�3�����b������6n9��j{����wj�-%c'j/��vh2�yX)5����Y�\3QQS�ҭ	H�*��H�ū�G�Y�9π��|G�=�
δ&F|a����ڕ��������(o��zMEn��|�9��ג�99�Ѭ';�-��v�P��޻��l�61��Q�ZˉhD5�,�>R><����v�C��B���vtr�*��6j��\@��P�C�p,Є.Қ۲,��yjt
!�pO'�yc�棶��x"�������y�&�bg�w�k����4y�l�OZ�j��/$��nD��������u'?�&N�Ɏ�Щl�?���BP=��78׌[��ˑ����� Ѷ
Cش{3z[tr5��
q��$�?����PT?+z�A��5p��D�yI�Y�B�RଳN� 	�?ش��S�6�?��2������Z���/���d�w����h�Ѝ��>����~�U�S��<��1k7�O��phb``;���A�ñ0�k�ֻ r��o�O̖w"|�������Q�t�M�$�����'���jym]�'�o�������C������ȪB��ׅ��w+qb�[�jCRH�X��P�}�o�/������e�l8��Ҁ|�S�
>�̈9��q3T�E�H���y쪈L	��Q��V�,�}�Ѩ ��e���U���TS2�
���6�������|^�+I�f�S��\�L�N�g9��e��)o�Ih�����ETD��E���VwY�� �u�s-iU��c�V�c{p۽M@�A���u��w˸�JƋ��w���7���%�%r	!�\�0$�"+s�����-I8I��ƟN1� ��r��;�5T!��tF"��+�|mԳ�\��iI7�����<�W)���w]QG-�w���2��^��Ӈ�X*<N�Pmk�rhzz	�9�mZM��3������@jb}��% 4�ν������`�B�����'{���'/
�����š�5��q%gD��@��2��e���#���	����ؑ;)~¾�!��td�#t�*	`��m���[d�(C��W�[�����Y��u$�����'
<l����q�r��Mչ�	>�C\�g�։Y?�}񽰗L9ֺ!Q��m�-w�yQn�l�m�b!:1�ޒT1wW�N_�mXk�Ǳ�B���Ʌ���^��v*�A{rA����Lr^L*˕�ge�!�|�},`ݡ�r&�z-К��b3K��3�1'H�@�QIFT�侑��X��f�+���2�֤|�b� [��7�kl��1��fH��vJ	�T.g��X�#�1��Wy�fڇ����
���߆�� u]"�;E��CiT�:H�� ����y�O�S[0��
��M�yЌ4��;O�9#V��f��.�%Ef��~.Tߞzv�x��U�T����������(��!�{�cT�C-j��+�\g��[ƽt�qՃ�Z���z�abi�C���c����B)�N����W+�2�4<�2� ���T:��^�������w�w��'V��?��%@@68"4j�#|�Ǭ=���uiP0��e&�rmK�f���9	�u%zҸ���^lxj�HP�V�y/rd�����V=aQ���d 9v<k����T܅ˮ����p�M���T�!G7�qU�$zU�l�%B3�义�����Xe�����R�j3�CX�Y���^���s���V�����<ҦyA���T�dK>����*���*P��lQq��.������0�3�(hL��,ڲ�����-��#M�C�Rz�r�b�&�P�)���O�/���̯7�7f�*5*��vQ5)Q���K��0�n�D$vw����E鑙�ͳ�qQ�XG$3��9O�
�*���o���V��}��O|�N��gZ5G�;s�/M�q�j�`2\W�ʔBS�L0��%�055i���*-�a\�Քֿ��22�~�!�ӫ����2qU\�#j����ɾ�v��3] yC4��r��|G<K)��W�/U�j�[��e��ϟ㨦w�p�w[w�C��{���7��QdNˠA���c��z@!c�*�N8Q���ӓ��a,T�ҽ5ȁ�P�����H��{+�A��A�Ze��t�Yڲ�q��@26��q=�MM�ot�� X�7DYr��Wg@���t���Ļ��w��=@H��r2�Y���/���b�����'��%���<`�7n��s�[�:0疠�چP;�V��� ����al�H΄��j�
�H���:�x�dO�t��.�Ĺ�>�~�I$�6؊$C�A�(����i�p��}��CRH�J&
�v���X�iY�/V:o��t���R��4��(�H�J@����������\�C�<qئ���x��p_(�(H��rR1�',��W�ѐ{�C Q	�v��]2Y9p+9F�>�.�>�׌�$g���0Q�<D<���[m6e�~s�j�3������?�F����p\�=�� 馎�Q�j��ʋ������h5Ib�`Q��E/c�R��C�cD�4�x�жG��M���oih��ӾV:}�J�+��}�h��pnKƿtt(�hƆu;��Q53� a3����,,4�#ځ?ګ�3�I�wA�Fn����$�#.�4��=�Z���9�K5�A�����z苂@�`��M(5pM%ܦ��x��UL,�6G�RPh�=(A�����;���+�h�C�k5��)h��^�����S�������$_i��m���"��Z��l��������S���侓���DQi�y��S�R�Y�F��J�f>�d1{Ԋ=47�e,E��/h�!,�7�����N�,)b)P�Ǉ���(���Z��8W:V
١�^�����q���Lj;����Ӵ��\h��2�G}��y'�}��RZ�Ԉ��H���;�0���h~����M��� �Yg|��o�9Zh$Z�a������д�� =ߛM��Iu�ʉ�L�Ͽ�w����ԗ%`�mI(e��<�v�����7�l
>N���:�:���w����I�Lg+�Qf��AUS�3W��o/sWt�sJh�klx�_�2�&hb���K�U����,-f$�d+>C�{`�khh��P���J�s�(��N�	��Y��+���g7�d�`���.4rY��� �s�u�W�N�4fv� �v�����-��0t'ؒU�	v$��H�^Pt���7i��}[ˣ=��Qquó�<�p"MGZ��"��R:°�5�t[��FK��ZD�㌉�+�8ŀ?S����dL��~'<o-�]�	o�ǜ��	U��T���΢���&Q2���Wo�=�Q�x2�j�G)eS0@��Չ$f�~�Z��9_acNfH�K%e����<h�hH�jctg�9	����:Q�[�l��,]�b��X�|�5��l�hlZ�H&'$�Ы�l�0��N3�e*���ʤ⼧��;�]�O�z��`!�%�jl8ю{�f�3���ڞ� �%�#B�ۮ��n��4�kY2�JT�.FW� V��]zF)��6���
�=�`�4B9�i%w��2�ys�j�S�8P�ZY<.��hwRJ~�����X���j��]qE:���g+�B��6����/�Ռr O�A��P6�~�7r �h�V� �ȭ#E�ȕ�&���ۄQ�F��8���j8�_����`��B����is&�Ì�㬳�NW����a�(Ύ~����]���*�ȭ鑧�҈qXq��)[�jhO��G'�"eǡIyܾQ��I��C�iC�����C���1��;��$���ˋܪ]|�Y+YC�{|ޅ�j�̪��"&ID�'�X�jaP"���f�//����J��ud�y�h��~�.�����ָ]���x�}�9TEѭ�(��lhP�2}�T�M���˨"D��KRhk��g��.�Ƚ�p�]���d�[�?�x8S���N&i�C>iI5���`��D��c1ݘRj�G6`P�R��쳠Ds<�w�|֐��F��o�
��kK�"(l���9bĥ0)�纻Ó�s�ͤ,$��ȗ7�����2ݘ9t����5*U��ф��6�%Oh���>��r�{�-ԣ����~'2�I9�G�	J��D�Z	��)���������~ I�e� �PNY!
Z_����Ϙ��	��L���
B��_%��Tt^n<�ǔ���|���Wt�"�� q5�%03�'�H�����~�kd��Y�\� �=l�ғ`��6%���e-	x{]DU��dS���?2>o:�F���n�5Ʈ�=���F��'Ş�j�e��&�^�~�)�{V��`�Џ�A��W�F���x�]^��건$��t�5�q�B_�'���8s��㾶i��$� gw�����~�v	w �'�#��a��d:�x�4.��;�	�^�rH��'$�sr����}a�/d���ڄV«1=���t��'��^9BQ�
CuhT�Q�|�V��`���va}x��G4T,X�܊i^�5c�/�q�5���M%�=�윸yA�s��ޡï�
�KlQk�SUP���}��O����9���KgJ�u��aȶ�JUT��DFW��D�n[h���n?Y~�BY�7����:��d�T�����)N��� u�Q��4O�u?�6��i�<JMlӈ����|�T�A}��I/���R�0ky�+:��$[�����W;_���x��4ҧ����}��`� p��+�"nq�n����]џՎZ,Eს�9�/��Let�MͿ�=�!Q{���*P嫡��$	{��+h�4�74�#��/�*꯫ק#TV{�D�l�e9���㞷p}v="^ 6�?�]����J��zV���3e��Zߔ��6e:(��#��,��@`��@#\����o#�8sQ���1�;��I��B�~Nnj�쓽�L��}�9e���Tb�͌���K�z�Lp��>�WO�x�Θ���s���ęn�)p<y�/R}{�Ez�f)a���!.�.]��@�����%O�M�����,5.��ѡƶڲ�Řj@��5� �L�u��rd�hҰ!UN�.����W���C�ABC��;�A���bLm�sjURpi��ׂ�=���a�x�F�#������Z��Q!���}y����yT��O%L�"�`˧!�u��m����������wY`���Bm���j��)�`[��>12DNMQ���W1��vإ�X!�u}KU�45+Q��眢�|F�Z86�{��!�)7��ʅ��N�!�6���8���_��A�ϤcE���3 H����fz��?7��TN�p�f����zI����%,�y�S���3�V�St���b	j��;�A4���Ѭsv(#��tL|�3���^J�**ѯ�[���(@�<p�~~�ׯ֮ܦ1���2��z��n@�`Q�.0�>�<^d�QH� ����ޠ�iud. Z�^�x�>5H���B7_�}^lL�'�|��.[JE=h~(	�~L����Q��_$i������E���m��0�^o�jh+UL�GO�5͝׵F=zm��"T�O3����Q�13�����xҼ�kk�:|�rTUk�'E�S�g��V��f\�,t�+N��
��SE�����	�s�(
�� ����3o�?�"��d����#��+�2�A00�²v�b�G��p*������(��'�6G���8F7)_*���D�Wj k��]����.�Ֆ���!C�W��8DSx(�F��!I��L�r!��g1��R ���K:�נ��-��=��'���;0.�j���:���()�7ǹ�;�[���Ag��?�:���CKt�ˆ9t�sP�x �!�����p��%�0^^!k�`)�*|g#1""b����#�C�����/j3[���!�͡o@-?��tq_�Ua��&� �R�?�)��nH%���N,�U�#��f:��0'�1Es&C-����O�-#�O�[�?�g���C����oL���˙�x�n��tj�U��U��#Ƨ��w-��Ǽu~(���J���Z\E�%��h�_��NM��m��_!Ȩyգ�� �@�U�%�2�̇�8��[�����E��\�׿��1�@3��֤�S����ȺP
�+�~�s���W��r�s1O�_�Ƞw���[ V�VF�/#��p{c�+��*u�M������p&�Sp�8Lt��|��������X_�/#�U���L��}đ�؋�^s�P���p"�JG=�В�8�O���3�M��7��HATtܹ�WN����0A\��?F��r�W�_�8E�d��ne�D� �a�A�I-��g����Šw��?گ�y����l	]��4OR���$p����E��^������B��o�[<��������I�z��/΃�W_��߀�D�'�ģ+fv��O�Z_U�:�r�ʊ$Ln3b��¢�.%i3s�1{�|�Vub��PͲ�վ� ,u���%��x���3��7'�N)8�+�Z�ӆr[H�l�^ر��u�Q�c�@M%�jէ�A_N�ᤫ�Y�~��<���~�V�n��"R0_R^�-��޻f�{�e��/��$�.>����5�l`,����3��~@����u��\~PrA5��@�5%���K���m�R�z���a9FSI�w]�^���s<o��I9����'�D�	�#=g���=��LZ�;�6��q���;O��j���C�z�X�R�f��.|8�m���~��O&����+a��I�Y�z�G#$�ۊ�Z$�+ he�(̾��&\�8ZF�z�|s(h��H�w]L��b@n*sʊ�7�E�g]�S�X�+]�oj���yTC�F��Iv� ���$2� T��7�.�N&a�����Y?>�"����ol|�[ry���HʞYƐ����w�g�l��
�%&�ţ��Fnˎ*�U�H���QRJ'����w�;@��we�����Ï�g睠��q���k5��*����Oڡt�83X����Z���F���۹��,=b���?R�+����7�{�]S(u5�Mi���@���F����}���	�Ph�MW�U�ꏫ���t����,m�ܛʁ3����:&�q��kiY��|\�Iq��[�染��R����Wc�"�˳�/��tR,V+� �:)��x��$P���8�ٸZ�Zz!�2�J�!ҰC�ά�s� p��^�fj�i5�+xwr}W���<S�7��ֳgA�p?��l[��M�Jm!8�����In76��#�:kUi�뵔F�m��|��Ig <y[].���U�5"]@O�^{X|5�x��C�(��C3o�&�����4I`xP�^��e�kCTfL�C�
0��BOB��v����� �Iї���c[Ȟ�\DW��SS� >���C�M`m~��0����*�� ƧD��H\ˢ_��Y{uN*�Jz`^�&�_����1����A��;�Uq ��=�C��}�oZzU+�
Y�L���CD��PC�a���~>1b���-;:n�� �2���h�V�_���Qy*)@o�l��v��	��iT������mX9Y�p�����"�[��ŗt�y�;�B�eu�8g���ҟ]Z��i$�����R����r��on�x��_	�QEvڴV�٧R!����!����&��.����6@�����w��D%?P�m������0M�?+�_@��gU +�0��{6�,>kR)�\{�#X�N���Wo�r%u12p`��ٟ���0���-���4cҿ�Rs��eF5cTc�^'�k	�
��:6#�\_Ո�l�q^GYyW���Lc +���L�W�����.����̯�pN����s�m.T�,�jZ�F�Y�S���_,�I'H�����#���c�FW�k^�XVۢ{שbOX'YglY���oEko���L�M!&�X�	)��	/���'�?zt5��\��<���oåԱ�pE'��)���������w?L��XʶQ������}~V &��
���78?} R����y�/���T���G�!KJ5N��iª���%W#_$( f�n��>t��c���	�R؀!����7Tm��ّI�Kl1��2R�t�?Q	+��u6�x��D��M���C��Yވ��M9���޸)I�9U�$+=x���ޗ29G��O"�[�X���&x�ғ������Vvc�TqW�"9�6�ӏ2%�X���wP�	��ɬ���� ��2�yjӥx ��V�d��F�$k�����h�\p��\��F^/u�G�&�.���)�w�E�A*�h��O��1*�fIA�x���w�c�'�o��n��� �<I?�7����Fw�Yv|c��i�L�Oջ�/{���,���72� ���øF�+�z�p؏O�E��}���K�-�;g��8���3Xo^�dH�o'K_ח���
��^�
�mʨ�/l�-ʑZҗt����:ݜ���H�|m����*�{ư�F��K����Ŗ�	������<C�MB�9�����~I�(�$0�˕=Li�"d�d�c�\��"��B;%�I��'��~ m��K/��B*{�"ƣJ�V��&>����&�ܱ.z�{����;�����3٧!����D�����҆�q�7(2pʬ4E�{/���%M�
�mx����yz��!��c"����c۝?��d�����K��uW�\�e͋�O�<!�~����e>rzM%Q���}S�0S_��1���$o��x�����M1�d�*1��}t7j�x l�;��8��u������-�7�o�0�*�=*�3���z�C�H��{�{l���
�Oԫ4�J3��0zG���	�a:��{V����O�ĉC��2o;�<�9y="A�ϡ���"���j�DU9$���y�P[p�܍-m�em��
�%�C}�\����::��,�`�5 ��@]X�l}A�ϴ�BB6��aA�9Y=�sqB�'��<^��f�?������~���6��8fA���xk�L�m9b�L�b�2�/3���$+o�n4x����4vrZz�|最wkjp�	!?�U@Ԕ'7�m���%��΄mm��Kj%��0��G^��ۜp�+��v��`FLo�a�f]�"9������aP^��/2{6A�M��$[��0	���&\��	E*0h�����c[�4��ꮵ�X��ɴNΎ������`أu�gaC����G���0st�Hy���q��V �L����;�bԼ�_��S���@�󺱢�E�mr>M���zL�ut�������9�k�'��[��@�Lj�q`iE�MM���g�V�j�R��5p�.�����o���=�=b�ag��۪N�QR�"�:���B� qs�z�n�$3X�`<�lM�gf�lȩr��m��z��Z�<�dXu�hB�h�6�\+���֞8]��f,��K ��5����"�"�5�(	ҍ����f�I.#�L7��z�Y�C�oJy3��������C���j���~�b5Ǜ<���ؠTӣ2���U�Mg$�e. �ɝ�I�0�[<�TV��m�@�^"B�L
� �}��5�L�C]>�R�9��"��G^�,��<SJ�՞"�[�Nh`�:Ǡ\e�0�pz���I��m�g��b��z��_�̽��>����J�v�Z��"xr`L�[N2�m`mV���������E��i�FV� ����#����Qæ�J�l�i��v�%�P��7j�m�5r)o���%+!K�l@��=~�?��v�嘑��%��s��ٷ��Ӱ��YWpp���QPVT���D�݀#8^V�
ǚN�S�|e��{�Ôge���\�!̻K� ѽb�)��A`�U��h�z�
95�w������9[�־�i���}�%*ꖦ��3}q��s�H}� ��J|a׺%�|�3�$%qp&�0�C,x�i/J�_������*�AL�>%\��=|���Ó>U�0Ђ_�����%)�
ā�{emG���aU����-���b��G�2�'�@��}�O�	�k�r>���B:��ht\8f�� -������#n�T�هNݢ��G*�U�� u� 6�,������~^"�Q
��Ȩ_�^f ak⦑�ܒ:�#i'͔4?����"��];�e}�B�YW�'r�8���M��\�h�0ԧ����b79*�G��S,c���G��q۩�}i.�6��X�hU�����˭Yl=;��P~�f�����b3=v����Ep��L�z�T�x���3�W`����u���qc��À���a�W���'%TD��c~����wQߦ�#eDR��(H�:̈�(7`�˗���	]v5�G�����8����)�S]J	\�_h�hzI�@����/���{�,�cEn��u���0:��Bg��T*hk5��5��@�;%a��Mq�(1n[�u�'��F��w䳈�IW� \��[2TL���F��"aH���2�s)~�ta/�������4L0��c��,�����6#�*�^��3:�Q���I�� ����i��j����u�K��̈́� �O��R��
ǳ/r���|�U�X@�.�Uc�ԅ�Hi���f���wٹj+��?���V��m�l,��Xٹ
T3��v��j#�F��z�� �bD�ddh�&Z`C//���~a��?�E���Sc�pb��Ҁ��/
����Q�_�|�ټB�'�I���B��|N:��@h>�v��<tu�o��ȃG���,��5�)�4ʑ[�l�Kb>�8�<���j�$�hj�IiȘ��i��t)�S��]7y���۱�4��<�"�|��ǃ�D��>�'B�?��N"c�Sܶ��qK�#�)��{�8���Z���X�3��Ʈ�s4�L'���q��	��N.�ӌց����x�5��'�.��`�	x^��� 9�eD���C���9-(1��j̎O��^
��%:��d������\�£%yd�YΉ6`�2%��$�;��J8�W�-�b!���?i�dQ���aNs���N��
lg_�l䖼�	�}�5T��r9U��W��7Ѳ��ǈ��j���!C7İ�`��E��t��ܬP���Z��x15�_�n=�Ry��	m��8镩������	�ښ�p�p1��b��oO��9��gs�7.Uh��>���"s��	#pq�DmA��3D�8�����z����ad0'p&|�0,�V�����+mJK ���
%�|����_)b��7��>�=D�[��YIBW�'��Vp
�D������d�c�9�5>��WS���� ��{	��1c �<�󏚭%�:��8����qj��f��Ϩ�tվ՞.$®'}B�̿����u���xp�7R&��;J��B����A�f�?�X�
Q遒���M_;�_Q6��s$��]���i!rv�����7�6�SܢJ�q{9�Y"��7F��B�a����������^��o����Z�����mC @�$y��g�ˆ���}��E�F/ ���i�)� ̟�����]C�'Um�^�p�h�85١/�)�j����<�uEjʜK5�6�<��������6[��FT@��k�hxKJK���%�ђ0Auѩ!A�Ƿ�_�?�o��y��G�:�}>A�v泷��]ia[�)�p[��bf}?��c���� �9�E#&u�:L�nK�o6��ʫy��6ӽ`̉³l��*{}��S`��W^�7�#�{�r�V3�%72��J\��L:�������\�#µDN��.70�:���"0#�1s�O����Ą�l�#,ļ.Q�򰁃_�Q�Ԇ�i�);b����i�������ӽ��!>f`/4(�i���}J"3����&�v�$�h���Y��e4�����(Ң���-��󄥦��ITύU����x;!�̙&U�SAS�ۃ�@^#�����c<�ᡰ��a"���:ĸ�1%{���ER�Ŗ�㳅�8T!T_�*�`��D������v�8s��/N6�J-�ը�q�:�E��8=�?M��/�Mb@<��mL���OZ��v�6Dh%�1�ë�ּ���/yQK	��2TY���������	�4 >ʴ#Y���3�X'��fOO(���-hv����~L�����|�V�l�9�y��	��%���
��G����3�Yv3P�$t����y�tp/�����Q�X�[U�)�Eӝ�Ò�/f�j�Pgː�mv˂Tn�zLAv�I"������;�õ0��������w�1��?�{�g+�Yz�i���Q��Q�V-A�?�2�}�E�I����4@�	@Yٌ���m5	���OT%S|u��n����ۮ�]ѿpmXи�_�a��(��JS��ۖ������XK�h˘�x�y��9��
7X,;�s�y���F�%��B��4�r�s�^{,i����/��	QX�D�yi=(�j.�sS���0�(w��}&8�D��G����c��0����`�R��B~IT�$LW'��0&?N$,����Ͼpu�3I�_����Xs��`�OpC�D��tPh�q�6`���"r���4h�(թw��
sm�~�?ڮV��y2=Q`=]�U�MG�W��7�m��2�0�n��{��G��Kz��S����i�_.sVou�\:�<:��{�C�[;5h�D	���#'����޿7�R�+�'3q�ҫK}���K++���6z>��=�p��Nd�`���}�}�!07[�|�I:8��$��;%�& ɭ`��C��%1��%�HؠX���b�sŔ.���z
:]���dzb���!@,�cHg�~ �K�`��SF ������;��� 3��&Z~/���up�������?��
 c|:�z�5�YGr��q�wv`���8<B��V� �>x�� �7���ܭL.І��� �W���.A/#�U�M�I�b	�6�������~Z#��t�'@�4��B`GJG�_�̢' =k8�'���BTW.��#b}֘Z���^��ôu���s;���Mhc�\G.f�Eb�rh�g���5-�
B.��h���D[+�+�`�o�y�bu���[�E���h8$蘣��Ǭ�U���Ti4�����^��L���%O"�(,f�K9��/6}�����g���Æ��\�`�CЄVGP%�Z*n��9�ϴg��Wθ�`�S�;�8�FK�ȫE/.Hac�>�C�����[��[FQʨ��G1�S������F�!���/�(���[yF�?�S�O�a��ϴ�&4���u�/���lA�]��T�DO���֧�K����^W���[�:���lD>B�~T��Q��X�H�,���ɨ������k΀�wn�\�I��s���5���T(fMB��#j���o������v�<���z�:U�yp����|�ow\�+��3�Gϯr${��qX��Ej�a��7(�»'>ؾҌna =�}	�P���-�a��_뇽^#o2ʱ�2�/!h��D�l�t�b��r�_����Z"�ܼd{����#���"^�\/l��l��x�8��\�Դ1~N���Ŵ��Y\�TR�C�?�o���j�WM���ȇ(W��� R�є��o��?��t�V����������!�q�<��+s�j�Gd[�3{�X-���8J���s�[6N} B��=$�2���wtr�