��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ訯.$W�7)�v��_��F%/���٨���)��?_CіP�XEmҪ?��������[VpQq��H�#�)jo�A;^7"s �5�_��R�_��d�&�՝ELu�|R_��u�D ��B�(�����߼/�.M���i�x]�n��+����aS�Ȇkv9�9a����YN�܏�-�#[1}]����[�$0@���8���Q-D?�s.w���ݩ���v� �lNȈ���]�4�^j	�1��6�j�D�W�^S�mxj��h�J~>��#����G �
��a��G"/i$���n�sɆ��]�*����~�[̬X���,��TL�c�n�;�:����x���$(r���|����̡l�߱�2�@v�b9��Te�!�#`#Q�~D<C�J��iB�0'?��~Тu�� w��J�y)�����^�X�����m�X�_Ȕ�BIe8ߕ���.ZKF�⾓��R��.�GڃK���)�`��B�&.V�_c��4>q��n�c\���?;��h�^[c��,ē�17i�¿�C	&�QZǜl�B��TZ�����pCT��0U������u��Q���xal��E�2XlN�T��2;f�2��`�%��`�v�igX(j�����T��a�\�����^֒+]ܞc��e�6Y�8���K�-�E���d���y>y=��M�4�K��F}��qx�[���R���Ĳk0���*��\Gb& �tԌ�Y�9�wߔ�b`����/]$��]hx�{��ڷ{ig�s�c����ۋ� ^2&���	��V�e[F{���/$	�fB<�ͩ�9�Q��}��	5V�S���c�������k�[�����0���q=�e��8��k�*��.o�j	�;=���p� ~���4�n�i;����J��fS����8��,9�,(�%� W���yU��޿�-5��ʠ������؀�1qgE�|T��M0�i��C]BW{N	�}X��䙊w�ѲnF�Ck��l=}�*�?0�E�CKn�"�Œ=mC�Ɲ!�<5P�����2q.�~Cb��sǜX�:`٬t�B��,�cUV,H��i#�?/ZW��V�<L�\���뵂�Uk�5^�jY���'�๯GTEJ��S�:����j�qO��u�k���숶-@�{�����F��A2
!���iA�e(�-|�gO��
�nL�����H��mKp3P$�ؚ�� �h�+���?K�U99y2����;ވPɮ[��`S(��1�l�΂��wy6:�k������r2���[��>^(1��o�j��y�:{v�"5/%��L����B�-q�(���Ze�YK=J�q�̀�@,(��\��N�B���?<y��i���1B{��Q:����c?�Q��&�D:f8�����T_8����Q_=`�4�i$q�}r�Xd�!]����X����Yơ>�G���wO(juJ"1��d9g�BP
5ۦ�c>�R�vC��R�b������xb�O���m�����,��?d�lg��`B#�eq����Gn��<�.Q\�Ҹ�ҫ;�9[+�FS�e;��!��K�F����r�������e|��):���x��NYu���p7Ӯ��4��7�[�[�-C�z[��|\z)�K�ޥ؏��	�_�8�&�b>��F�{�)�߃-jd퉰//�_T,* D1j�@�Q����8F�j��<(H���<�9�,�Yzw����������O3�6�}k)Q�[�#��~I�Z����ll���<I���� l��He_B)���xt��N/i�PM�+Ď"N�k$x�?�i^@E?��D�2���̈����5�g���1D�ѱ�Q�Y]���s��15 X�eA(.�sMޏ����Ch[{X��Q��E��f�2b*�"=�����I---�8}�W��Ʀ,��>�:t=��G��рg���9�Km��~����CZ���Z���M�� E�;x���J\ŃXQ|����<�c����S��5�H��eN���%`-?q��f⪦S�ޡ�!������m�X|fA�����̷`�+�!�ϑ
��h&P�\Q�P|�����'{�}1U��X�L�{öC[�Ќ���Zo������Ţ�#b��s����^���\�[�g���=��uن��@%
��P�S�
�P���?>���H��&\���[GHH~��=� d�J�d����
����Q�_�x��r�H,%��;���G��w�t8v��{譓m����9Tƈ�ȋ����	�2W������>�'k_Ա+�k��r86�$�&����2k3�@A�F �UH�y�����A��i��g7G�f���~�g�$0uvEv�4��a�*/�o浤E E�q�N[s��F��Nܰ�����cH��F�5���s���
ԏ�.�@��!��\�͟��i�����GҐ-=YKxi6Wѩ��7Z7pE�K���p�<�S�mfߤ��U+N��q0�Ǒ`1�:f&g�Dd��AE.	dЩҿ�f
34?
"��_.�k1���Y��s����sR���)����x5Ȑ�0�7l˪��x����ﱯXm��%��H>�&��w�+���ؤ"M�_�f׭�_��v�&���}��u�uo� 
t���c�5��\WAu��%(i7B�ә(u	\0�'y�th"P�H�����K��1aMvS�}7t��T&\px�3�b���?hL�=�R�pa���WzM�RWx��$��[��%�LSSZ\�/��ڱ,s�Р�����c��WH�	M��4�sW���_�F��q׎������?�k1�٘bmf���-�e�����u���9��Q��?�h���n5}�fJ{�s�;ϜBc��Yx��U��07t����|��I�/lt�=ō�a�&�^���A�����W�i	�����Sd�0	W7�7�%:`��A� 7óv@��+l�!^E]����	!��0>�9�%nc�y�f�6� l�ЋL��(�<զ�^�}.I1t���$v	OJ�� ��b��7�Cl��P�شX�"0��8jط�ܬ\��L���ȸpGkl�
d}�<�;>�hF�j7@���2]�b�=,���];p����N-c�B0ŭ�,e��'���?��<�7__�:��_ɭ/tHS�0�R����M��OEݩE��YF_�:|�A����gCo��-~QH�#����)�/tz��	�����i��褁�	���%�Xs�yۻa�uL�J�´ɵ��\󽏰62�Z�M�k亍_�e_*i���r��N4�Q�5�[)T���ㄼ�?�uǉ�+qѷ��>5Y.����:��#~#à;�M���c��I��&��<��.��t����05{�߆�t��V���6�3?Ӡ�,;�5L9W~o�]�pT��u�����X��_r3u�fT�op��C#�A��ɇF��ǂ
1�7ļ�����|^�!�� C���@��#��0���6��HJ�(�=+'mGc�����Dm�ٿ!#y[�6Vt��=s�?Z����J>.��j<O������,�/�����~*�+���M1�]F�
\��6��������,-�]q���Knk6�(`�Ȫ�~	�>���|�
D��ҬY�����vꙉB�12���UO�����l:�P��Mi�
�l}	�M�)>�G^p����lQ��N�T�"�@"�:�:�髏�vr�d0V�l2]�
������ofd���#�k�҂O{���+S��D�f*�ڻ"���Ws;�V���k�كGn�A���m�ê 7W��`s�uz��X�Q5f<���f[,�k��#0��In�O�*L�|_��!�꟡�� 
�d	�c��~�%��;��D��o�sA]��mU�;����VgH׶mx�NB��i�}`�6u��RSIR��߲F�f��/KG�;� ��� }��5��;Ͷg_]�$@���
pK��=��� � �����,x	σ>=H���e�a�9>���������1�#q:��U�UH���w,�ө5��z�ex�.���І��xj۩����]{���{����y�G0ޫ'�^k�`|�"��Z�;~ϣe�х,�N�2c#�a-�z)4lV��$�)n������M���Ґi��HbJ.�cs~B%�o�����y����/Q����j���*��?-�G���Z��w;��/�p�/s����ˤ�|j��g�����զ�Ԩq�_�^��@��.#.V:nUř�/�ʉ��صR#o�����_'X���Y8���<���{�o�;�h�������%o-=�95	1b�����:[�r
p�����Z�ĵbX���y9�x���~.k�YU�"��g{��w�4���F+�zx+�o-�ėp��1��Ή���#�[l��Ӻ��qwqFd�Q�$W~�M���x�U �f
���ѴEr�`�Ҧ�0V��)o���K,��_�M��}u��l���"�Ba2sپ5����T�g[OM��%3Y�TL��nN����تe[^Z-� �RM�X���g���,��㠢-+��x�.��uA���T;ؒcl:�"!��)(D���i�gI+�c*U�nN&|�r�q1��t�L���Ϣ���[�^���r��S�ح'�g��F��@}y��9 ��8 �YD�
�rR��Rݠ[��.�W�:�e��Η�'h�
��نߝ��@����I�������=Jx#��껤��g:j����t�!�P"\�G+��y�{PM�R(�Y�RNw�ì�a��4�y�۝�3��˴>߃�$u���g��=Ï��g�M r=?�3����M?�Ob���F=/��n�LJu��Q���h��L�3��yCXI�������Lw]�F�Ի�KW�o.��.�$Q���%������N�Jn��'����d��{
AF;���W�@*CW�5�ȩu��S )O��[cv}C�Y T��e	�e���f5���R��}�\	�In �'ܿZ��=@���i�V�������Oz�I?l�g7}d���ST�a�,���$!��b��\%*�0��͛�9@f%Y��G�Q	o7����d��ח��g<I$/��14'7�s�D���I+D�u���MM�Wm
�k��Z��G(80A����8��]���z�Gs+eߧWQ.1�(��rMxU���4�  �i�� ݑy�`�q �l�f�-��$2��K@?�x�#THI���-�u�2��S�:���M�?�/!�jl���*ϩKH�(�4O����6��ӊ����4Sj	)p;�֟��^;9���$f?��0#���<r����D^2@���@p��tb���Ԉ�?��zM��o�y����|��U�L�3v��0����X)b3�?�u���: Xj��+�vy�&�k�.&�]ro��=�@1#� ћ��-E,H,���^��^�x,�����僨U$o�ww[��X�x�C⨁��@���i��8#&.��j�c���~f��K9���Cd$6���G5
,%S3kA�i�u4����+:ܑ4�={�a9ۭ��<�Ր���=��I��k��0�I+�E��i���?u��q�
��"ܩ�³h��'�T2�,���؏ˁ�[�ӿ���
�k͔�����Q�����D|��d�AbR�khu��6>�M�;��❄R� 	Zv�aÃ�a�'k����P�&$*)5���Y���
-��+z��0�R��u��|!���9�t���"F��1z����+##`�2�@g����j
M̸�h��K��FY�(����ˎǸM�������1�|n4I,e�!R�;,l��ђ-��V��;7%�hX{3d��[��߭�;��=�ᢛ�P�h(1.0I�z5��:��~�}\�L���VwT&������35ǑX1%�IL��K�ES�'�ߌ���Ы���^�}�0)�Ͻ����������w��(��>���Lǳ�]�-�_r��>L��,&>6�,wvt%�~t���Ѕ��|h�3�#�;���U���a+�i��E�Ofp�jd�Cd|\z �Ť��ט�7#s;���6)�#�S�R��[v<�#�[�G�_��9j�`�mq�/K�E
K�ۿ�w-�L��jE���>(�9$H�s-�Ŵ0�l�,�&��v�C�9�/��o�'�Ld���]2�eJ���X���4�T+�}=��2i���KX�W�Еu�ڮ���N��+�����yH/�iq��Qz<�^8��ፙ��[�����s4�%��۪��W��}��0��!���7�� H[T�m��?�S����
R��3��͝���c� <ol��ưޫ��n��Y�,{X��JF#�^�-+Q\E��/�(Z����z?j�.�	���[lz\P�(�<k��6:y;1G)a\�[������D.q���.�\�z�1�)�TچNt}�u��p�=r��u�.�	M����)P.�F(�/�u�8d?��FGƔ�lvy -w��l����4�؉��U��K'�b�h)'M�؃l�o�,j������V<�5$��i��'e
�T�t���s��̴˓'�i�������� �/7�y�Pc^�&f^K���953�s�[��������i���������$��8��I_Wc�&��nz�]��3���W�cC�X�;QV��	��c��Բ�4L�( �C���Zq�N��ε΍��!�o<.�
�q�;�d�D���`nmFv�D�N����)�!��fS�~�砙��b���Ғ����~�.��EnOeI�n�/z/�Z�mɟ8�(���� ����~k�:��.�*��E`��w� ��c�
��pN�il*O��f�i�4��4�`�o��X�X��;b�Û�L/���N����)�;ּ4�<�o��S�r9�X*h�lb���Ԁe����z�Sͣ�����Ɉ�ZH!���j�����'+�W�����֣����=R��\_�?O���5��B��㒩,�aB�-/D�`8C�Mķػ�K`�}��o�%U|�ԍ0�D��V�Q;�R�bA�7�vC����1�/�i�	{ǘ�!��`�Ls�Ϻ�{��&4�ȑy��qڼ�b�7W���S�|E��rB_�G��5�Vq���������+Q_�X퉭�1�J�&#�,��o��ݿ�?�%��bA��O��2&x�@H˵(���k#J<�<ܜ@���B�@��":Zv/�Φ�Ҭ՗�ʶ?���9�$�a�.QZ'�o�+7P�����@W�3c{�#��kM�#��^#�o�S=��x�k�r��Ǳ0ƿ�P�W`�w5��������Z�o�y%�9�@:�����Q��8�>_N:��7R�#�!�tL���hW#�H�j)z�_粒����
p'Y�;=NMm_�̗�]��t�X6IYa���eϖ1~3n���M����0�-��9�g�X�+��OvO}��\1|��8�8'�-
#Be@�rD�=�fZ�C��&�T;�~�f�e��;��*��A��P2(B�^�L<���!�73���G��.�C�Z˥{�o�X`{�����I�K��/KȰ�-1d��Ү<^�]j�/y������-vsb�x�<�:�KO�D�����w�`����TI!��[-����;� �Mz���l�0��L���y�=�������˚��*�:*�! �@��� {ͣ{5�uJRZ@{�d~k��ט\��;�Z/��*@7�ʷ�g�,�R��������t��L��+��pj�U��Ay'�e�P~ͦ$;��ԯo�D
q� ������]��ǡ�j��a/48(▱�etgJ����6��$Q/c'G�A�eq{���J�/(���au(*�'LƮ�OY�A�'��2��rh����(F'����������x� }�^�}#E%�6��`����C�"tN��!/mJ/��I���3������C<�AH�2�(��Z�8fR��M3Rw�6b~0��R6�|���7U�<�����M��m���`ē�������r���~�P��n�~��VF��么��Ȧ��d�w��8j?`]�РK +�H��#�p괛]��4-�����ӟ�r���l�l�������b��DD��Dc7�i|��K�.����[@���7} ����\'��~�?�����\>W��O6��Ki�����
�����3�j�i�[q��D�YӢ��X0�Oz���\ۚ�l?!��Ơ�{5�hvQ0�Ϟ�#����Ӎќ�%�I�?���`��,�f�F�T��vOG`�X�\X�Nu���I�{���m��H}q)�z�|c�&��_����$� S9]:�9����T:C� vf�no�*�vPVD����>��t~(ۣ���`��ҵ��1�����dz8g�D��wtp�G�6��TS��}E��ȑU�[�ܼg �B$H��稳�(`Ԍ�����^��͖D�fq!}}�g�V�V�"t�>y:N\ 	�=�rZ�W~OWgᑞ�Q�K�,�	z|�3��#;�1v�[�� ��t+�~���+/;[�,Q���Ş ��5m�rU�T��m6�cP ���֛D��1�h�%�c�ѸA�B:�eE�Yޠ/�݇�g��N�^m�a)��6T���xCZ�ļ�d ���L>t��e�E}:��i#���!��@U�_JD�h���V�K�{����cٳO��!9z�p�M+p��"B����t��8B0��j}�dK���,/���ԛ! ~e�����P���|�bŢ�$�"ז%l)�xcY4���7ݶ�7�`�k�3�R���z,�H�r����G`PJa;Lń�+�U{r� ~�[�O��Χ�������0�_��?�8�d$ŏ4�:�5�W��u ��<hk�)F���)��S�0
�-.�c�M��Sː��I�3y�{���ahb�`o 3;t���#�>�����'R��,��W�p��m���u�黂I��H Rh�j�W�>Ю{y�P�'I����&,At+�bv���?���������x"M��٫plx�%��O����b[�72oV��A�L�k�n��9�#Ǜeh(�_4L�$�P�&��]n�4t_��%�W��wAU��P�R�(���0�"Mx�Y�Q����%NfC�n$@ 7�v1�[��R0�S{Q��+��l��0dJ;��lMM%�`[�=h�q�ОT�_�U�2�����|���+� �� �D;l�O�M4N�Nf�|^�'�)�G|����A���݌�?�(^�#gs�6�w��6v�fβ3� �r��5)!��h�G(�#d�:��.=�xE���&�ߪ�q���w�	@8CL�H�,��ܙ�!��"���%z5LRl���-!z���2x���p2��%�<���ϔf',��'�է�ۢ���L�H?Uz}X9�NM�kվ���PGM�l�%�eF�{��*����K;.��b�QIb��%y�y�*�*X:Ҥ��%�~���:�"�a ;�r�Z�����2��a͌����?� U�Q�CW����cA�JZ��`�F�n#��g��ϯ;�&��M�P�C؄L@��!Y<��W��Yic]��P��L��ކ���cQ={���b�=�%
^k�F�&<�g����_��c���LVu�aS5�ۈ1R8��,9�%����#���!�u�Q�mN��L�J˨�a(��H�Ɉ3�0�T�B��G����H��=z#k�%���W�M����_���hG�y(L̿hH:�z9�7��v�H%�=hh�O�O~���8��v���BK3�o�ѩ\���xldW�?[�;N��pr?3�Rf(7J����tj��;c�k���i�ܴ�APNfũ{K��X��Z��'e̺��`�P���v����B,Y�M�C�\M�)�$y�~tnm�_QӪ9�=�[I���΁������ !�R�"�������)h|��`�v��S����ؓD��!g捙ܗ�VJS����!.��h��-��5�wx�L!���`}����쐌�(d�*�fH5d� �x�WBrAr���{�?U6o�ωx�v���������H��i:$e:�B�;�m�x�XF�yg<��|�xHQëcQ"L��ϱ��f;Հ�L�I\wͥ4��5�Ur̋k,�1N�~j�/�d�)�����^�x�KҚ�n��G%�>���i���ܫ���J|���%���w�P|�����_�/ԗʲ�2cY��n�^P!3y�jA�UFp�,�&��s�y�B���:����ʺ ��c�a\�b��Yr���N �lE��9�_��
�՘���e��0��law�"ip��h��`���7NE�>�c�m���)-�aK�G�sB��w�]�Jm�M%DN�h mm��ML.�d��k;�'�?��
�:��`D�C�yi�#�ީK����[�D�������F�}@�6�#ٯ�>�7� ��|3x ��u�Iu�,�U��u����y�r��4����~r�2��hg�*}$HcmR�Fa�;�7h����7����X\P=�U����k��)}�������,U���&�9-gg���2+<�"Ι�[��rְ��J�(�`n━������u�l(���l�z�Q�&?�j\�}'�;�EI}1��Lݩa4�ǅ�P��+�?����и�L��n������t���`��	_�l&�{1(c��uv�|<͟�{=�]�^ě�:����Xٺ��m�%����fC�DQ�c����'4Cu5���$��#�O�Aj9����7�E+ ��]/�U&�L���	��},pM�3�Y�jc�@h*5A:��(����H�G��Qͭ��Q�%�6����d������
�����X3�Ռ�s��M��p�m��T=�a�p��'| ���[X�R��u�o[A������ �4�ɼpF[��g�.r�f������@d�j�����,��z�a�FJ��PΥ���']DÅ��6^����
H��'g�Ƈ�lڱ���|���-Z䂠��c��G��jC��ͦB�����*Z�p0~[�3��7�D��JJ���pV�I/g>/(`eX<7�s�d1 ʾ/�Kx�n^K}��S[׭ 7l���8/a���ƚ�
��K�g��