��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:��������uA��@��y���<����xDET>��W�����C%�=U����3v���hj��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0� $���ƪ��?��֊��;wJ¯���H�����؎h���DՏV�>j��ˀ^}>=���9�8B��yj%��,�C%  �,��X��TDS���l��2���Ec�1D?6����:�����	�٬�醖��W�*�ڊB�e���.�'F����J��$�$��m�r=I�=����`Ԯ|�Yo4KoSׄ�,�EB��P�j�,T)���?W�wƯ,ȹ�[`����@�����QiG*?��V�A<�*[udrI��H?���zٔ;�;E�����yI$n�d�f��ט��HL�����j��B����`2T�%#�U������ف��?�?�sΓ�&U��YʶK��8�&�Ť�R�����X����7',�'�Z�N�fYX~��u6��w�h�.����&��D�������S�׻��'�����XŨw�%�؍՚�@l����ۮ���I�Ik��Z?�q2Ux��3Sb�"��nX�vbd���s�xd|a&H��?���M����"/���I�ȚVv_�L��AA�+I#V���8?��|P������e��ڂ��`��[\0��\Cm����$Q��9�wh7�.��G����9xMJ�Ժ�?��(y��Z丹���ݫg<���p��8$ή��4b2�Wj%���Ê��&�<���b��=�`�M��G?�ހ��s�)�9�G&�';�E�{��-Ëp{܂�ry#�񙡡研��(�]�-<���Y��������ϭ&W���~��c����s�����s�M¡9�)p�`nݠ�0�w���Bvs@�6�LL.���Z�U/�?��'��V���7�ᅣ1��j�6�#^S�Ҕ`���>O�˫��m�{4(gn2\��U�/m�)�q"�|�0
���wϹ�PL�@p����w�ݤ�A���(���J��[�S�N~!9q&^��z���wg!k�F r�<z�]c�(8G����t���0��b�����{y���3D��)[AG�R�OXz�C, ���]+]" ��:��ɚ�Ǳ�Cc~n]�x6f|\�ʧ��h
4ʼ�T�������b)�J0ϕ��jP)��@H[��ٶ�<�T> ���ÿ�HPf0�u.��e��m#�<�\`�����'�gc<�rE�<T��������g�&� ٴP�_�6qrۡg4�'92!ˤ>n��[�k��sr�Ï����fm�c
�Ƹ���^�.������EE��s�y보�j�"�"�m�@��0��I��,ݕ�IHd��ϐ���'�~�ԡ�blVh�`��%2D���j(��R���Ӛ�V��S��)֡,�Q�X�5Q�����A�R�D�Φ��o�FE`5�H��W�C� 8���D�0�� �w$�F��7��0tM�#��(9W	�,�����<ȍS�4�3�8���Dd�	i	oVˀ��c�*EL�괬I��Y��DFˮ2�Gi�ֽ���-���*Ό2�t+���I����3c�Z�.���h5W������ �іLf�GA`�0<�{��,;����s�g��y[6sf��L����+z	�/����w���H��h���������}����Q% <�nl)i��^�g�h!������*,��m=^z\R~B{�*\~�(�W��u��x��5�RlD��>�nA�i+[�`��1Xg-Y6����X�DZ}t`�����K�1�x�M�X'4P�I�"�x`g��=d5AB�vh��Q��)5�8�?�VG�6�r���XV�إ�Cě��"N+�Qeȋ�1�d�妔�~^�i�;�L�i8���W¯JU!%.p3�O��O�
 e�����ٛ�j�Ij�8����$��9"��8L6O+�����8�K7ga���#N�1��@����O)HVd�%6�����;ͬ��7L7�f��}EHڱ̓O�ִe�K�DN���aV��d�a~÷+1W����2�����͝z�`&k�k�U����P%�I3���KO�uDk�>�q&��D7�.��?!���w���$�e'n��ß�	/^ %�B�����P��������d���N�N�O<n�WIܶA�3�`tp��WM �cbKA��bF��j�J����Z�����.�(��<J��;�{����$C�ݧD侕��sw֭�y�=B�HqyE�Y�/�x��]ƞs�|R��ߐ&��Q����ݍf�0���±ǹJ#�B(dX��Z�=L���?1���L֎���7K�w0"��Z����
� �y0�l�H���n�ȁ2M@������\,\��� 0���ч����oP#E%�T�G��Inol�H/6�5:|�$%�^mp�:.X��*�w����!�C���C�h�T3?m^��wo��F}g�5�<�?^��gKS�>!HP>�{��	�cb[��+�ED��F����L+�����vI�$�U���'e���1@��z0{��o���Ƽ����J�!�%N��
��]U��T�h��f���UY�'��눓u�k�>�Ǫ"X�{�1�1�����8��,N�F�e_.E�]8H���]W=[���L`�m�fN��1E����i~�̣����/���� �4bo�0[Kr~蹩���F��9�(m:@Vw 	b��;¨��P��>P���t�T�x������qmw�+.־=|�S��M{�މ);��KoaQ�F����jsPp;=}�URR#�,�|�6b�=
��&���,�!g�/sڏؖ�(m�q��ɝ_���E�U�*�?/ �@B��� UfO�2P�#�1�C�,,q�zy �4é��6;�>*|��x{i&F*�$)��rk���J�̪7�[�W�t���v�AG��X��i�6���]� ~�/^�u���&��Y"��"D��#�[��c�M��w�o6�}�>@���6����hi8*�3W�A���D�"�(��`QOY�ג'L#C�������A��
]�ʮ&}�Z�>R 9
�s-l��YPtC<�y)�H�y.��Kh;
���&�c��Ԣ������{t�a����u�R~y%�o���l��|u� W �KWbY�Z��'�&h�����L�=����q��h���)����_,.yo�L�u8sL�U�2s�ߪ)U��`�*�2"S��[e��On�O�."�!���M����R�S��H��)B���k[�.K�<'?�XE�(�dĂ�s��c�@˯&0V��ceZ�����<����<Q�� \�pUuWѤ����v�p!�u#N��wʼW/��ӳ�O��KBDE��nw�E��*��p�q��('/��,��,f���_9N�3Hh���Yn�p2����^���R��¨�w�����J>���Y�1���S-��7�7���bV��U�@ܓ��w�&��(%���!����v^������ח7���O&�0�,�kG����ƽ�kѓp�����}� ��~|��ݘ&�!d���=>���ë�4%A��vV�;qb���C��������Ż{_�kϧ��ԁ�qm��J43�1�/Vc����M��c�����g*Y��3�s&��	�kdD|29�X���E��r&�-�4��s+�$�3a� �#ۜdߩ8i�K�"���;ă�%�ؗCI�EI�+��m��'
 �h+��(�ݿ��<J��ނ'�rᵙᄝܖ4�Ǹ�b� ��i���P�����"�U�v�G`���aB���!TY��,�&`�"
`�z�92r��ȽL�ƛ

�	8���dP���h�KJskTd�Z�4�א
*�mhp�=RRs$������� ,�>/��(1Ϥ��
/��r	Tt�2��A�S�_u�p�4�1����+�X��H���lW֡F�-�^є�3k��S��5���}^Ԗ'��TE:C�o]�C��c��~D4��~��W�Z��y~&!�eo+Йԯ��g�(` �;��S�n��m1F��,.2M���t�֞ӫ���3l!�:���^�j�~�E|aH����W���]�<f����C��β6_�^�����f>_x!����pm6��W��.Lk($�V��_Z��Jm��e��q����S��������"8���Q�by� T�sl�hl�����q|������*Y�*#��r:.F��m�4MQz'{��
U�mQ-�"����]�hж�����~������\bC��@5���(� �Z���t�|�����щt��X�N�x��]V��SM��ɋ���^>��D�Z��Џ�`�"h,�tA%n���:;��뽥:�[�2�n��XF�_��b�->/�(�B��,oK^PK�8���#��a�q� jSXSp�6� ������8��>��p���*u}����Y�_���T��Ճ��Ga�ug2��E��Cأ�������������K���8�[d˦Vڊ$��az3}.f.�à�~���O͠ �h�^u�	%�8kҼ1��,���m�����>}��3��Wyψ+����?�\���\O'Y�Z/����5���;Ғ6c����.G���sŽ~��]W"\��h�W��B�8����� ]��Z(�\�_�����E)j-���W����=%/�R���.����k�Dp��\�ǆ"scʭp��cX����1�����������D��I���l�l��_]N-��j�L3�i:>;����~���Z��h�q&���L`�h�eQ���]>=�Ɇ \9ti�����L$��&o�Lrd.7 9�������;R*��߅���f<�L�1�c���m)�@��R��%��v��K,��䍛���/젘��C;�n,=dw;GV������2)-f%'mJ����#o�\A����g�H����Ӊ��!(T2�I�.>A]"��{y2��j)\���,�]"��v���l�B��
ndֺs#���*Ce|��ʓZ�7p���>q (`GP��s(�PL�$�.C�������Q&���z(�R0ϸ�C���Tc�o�)a����*�u���~D֚Ӧ���p���p�bֈZ�f���1�X�Y���@��E�Փ�~/�ܛ35Bм#��@���$�<O�ն�����n3�����?9c�>%�B߮���A+m�D\���p��Xօ��(�WrĠ-���"M������y�E/y�2���0o*0DQ�$�i�Q�ξ�I��7��v�,%�sX ;f�J�>ъh�s Ԇd�SsŲSĮ��cd"���p�i_�aկ%��`�tCY"F�Q��c[G���� /���a��f��R�9L?��Q��r����$>t_4�8m�r� }�V��$H6�eb��#� Zl���=���n,�&W|S�,�~�3�G���㑇���6�n@��u)������}�GՀ�����2���gL��*v7۷�)�'o�U6�%�1�2ރ��2�H����Od��E�>�Ӎ���xi(]���U�hD��3�z�f�\�v��|���L�P��j��%�:IT����^�=$Jl<�=�.��2�K�|	h�A$%�ޯwQ�ǘ�x�{c��[o�P��e �N����f�%�W
��w�g��"ݢ��3ip�o�4Z;�b(��HX����H�٩V��(M�J���D�H��/K�u�:�]��x����Ů�':#r
J���N��)��yz��>9�;g-w?���$W��a�r8��8�.1�ov`�
/�%>��5�(��˱�Vר��g�9��]�C�����Y�[�og�Rx]㸼��1��@li�K�=c��N��d���goz4���o5ao�a���jiG�����K��YyA�̀��=��jx�П���gRܢ�X4����+i;��z��Q���8q�=voW*�+�XP���z��`�YcDT��:rg^
�!��6ZN�[��о�{�%~X$\��EHu,��35�A)� 20�ǒ~�N��x��L�j-*�Ѓ�c���z�p7��݇��^BK��Q�����5C���i�,xLd(�W	8-/�*�f�]`6�7����YC���Y�%�����{R���˳"�-;��}��{�����r�6�ƃ��y��A��o�.����e�T%;]��]ϰ��~�f����12�|\/Բ8���N��^��HN�^XM�