��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������<�R\����nC(4�h�	R���\���?�����qqD[�S/�ȿ+�
F�m7��A��g��W9I���%b\>cAyk7�'�bv�(��mN�0������8=r{<�;5��
h���4��Ʊ�x�f���9XF�(n�� ���¯>J�?��W��U�&�w!�~�;��2�Lkt�1q�"a��|���(�jx��͊&ő-,�^�-�D�>��֣g�*����ݓ0�ӏ8�/��ļ5s	+�f@�j�H�+>*�X�sƼ���p �)њ ;�F���V�������=`�ņ<���7�䐘����	�����al��"v)�>.��R���K8���P&=ۨ��6�,�Vn��k'(`���e� ��μ����8"왗�l\�ŒguD���oi���~d�uu�^vr�TM�zk��,j.M�����o�P��]�����h����i
P�@'0�1"�%dB0(F	t"���A&���ԓoO�����^��%ZJ٠�3�-ԁ,f�W��}�}�'�1��G�K���*nU.u����1���Z����3�6�:�����M��xHP<6&�$ϒ�f��
0�?�0��	K������E�B(�}�&"@������,��7xYfRK�)�ik���М��w�{.�虈�d�-�d��P�B�2d��K_dŹ�[�%�9��"q�	sШ����R�eKe�U�"�. �yx
\ܧ�X�[7���nl��^��x҂m���}��5a��0Dr}��?B,}/��",�#�m� �1�S�����
3�?e?�ix�d~�B|gԤ�D�"
�%K��HH��`YK����i��DΧ{q�	1A7�P�e>�L�U�^;9c�]ߏwӳ<�B�D�R�j3�crI���dZ)�Q�L><C�Z���A���?1
KZɍ�b*F������R3��ϤA��ָ��� ���eS�N��b�@׍n���YPm���z��S��4���:�Gbe�>w��J������]������5���e��&ߵ��_��Du�|
��k~k�7b�n��VO9tJ�� ��K��>��j�-i����giu8��"�%$�t9�<}��J���n�ʏ���z>��+~��#�蔬0^K�g�Z'!���F�������}�-�n����(Vj'�dK���TK-�I�<HL0��	1��FZ���3�v�.Y��׬ �0�t3F�ʆ�F�dK�ڇ�����A��h':fA�{�s�G{=��Uq ^�}ߘ\1t6�U��W4���lk�!����̞�����,�.�g���Gd#L����yCQqrF�U����D��H�� ���I���W{�{Go��b�A�����s#��NW�ɈY�8��<���\yst0_�,����kꮎw�V����U*�NE/܁.[��n�бW�8�=�_�=E����Nƹ�ʻ#Mh^��@`�h �Q4��CN�x�#�N�����@݅2����E�ּTbð��x����G���H�B��%����E��`F׶�}�$����Ev�t�m�Kk��e��U�6ɨ�5L�t$g�|xR�F�*6j��-���FB+I�[�#�Je1�2��}|��\ɘv��;��Dl���Tƒ�������^�����ɪҶߝ'ůוbt�7�;%28�5�*M�h��Q���k��[}G� ��Ԡ�����f�݋p�o8�A��67=��+0�aG��ᓝg��]��4�؎�X����
��o�|�ئ��p�4ẚ�8�G:�)��d�O�h��.��� )�v�.��r�4ޱ�e���?8A���mc�p�~���5'�֍^��h<��R���yd�\*2�G$���sH����/1���X�:yA8��-�_{������D9�O%�m��oƄL�È#aA�+�xz�T�P��I�7�Aݤo4AN��{�{K�I�rVz̔xL�4cpQA"��\x.6~����G�ʡ���sַs�"�ix����HC��
N/\C7?�Vm�c�6y3\5�Oԕ1Τd|	����í�ٺ�T$���x��_h��&�9_|FB�\���_a�
=A=�/K�Yo!��2̩�bְ�ǐ�E�t�䞎�ڟ�Ⱥ+��v��~��a�=����"an��3�K��D��+��H<��2ILԩ~<�!@�m�V2�h�8R$��� FS΄�f��v~��P�Wڽ~��-
�8�.�	���*�E�.&�"� �0�|�N�q���j��G"�������_����{>������/0s���r `0E��3Uhmgom��AS9ׅ:|�:l^9���Ork�,U
[l  �����ob�8F���3��5��P���g�C F�&h%��H@B�ƕ0��*��W�'���տ{�&MYq=�6o���u�����$���E�Z1�K��%l��ՠw��|�K�`v�ͯ=L}i5F%��e�a��J1*����z����i�|$"�H}=MRŲ� M�	����~���8���ş� ��V�< @p��Qn�#�Q�R����	��E��ie�R��/! nڴ{w'c�O��9i=�o���fB;]���d�~�`��{uX���QF�����(N,���@S��algx���,Ӫ!}�6�!ѱ� ��~���Q'}���Ju�P��`g��>�DB&N�JQ��v��x���f����\�����B��u(g�+�?{�kzSs�*$ �;��/�ީ��O���6T߰����f�_m��]��T�t�I���(���@�P�䠡��g�n��"1X�Ot%9S�w�)���ӏ~C�e05kŻW��6A$ ���|yLH�2PG�����<;5t5�&�R=��]aj}�Rj+G��׼<ٰ���������bDck�0�?��/R��fn4Ֆ��Y�����A^�U"�R��-̡��=�;��_��ț��u5ۉ�l�=��ںG�w3���O��HZDb�}J��{��Xܳn��s{��S�F����G��b*GꗛE���M��ug����c�V,�-��X<>r%��������mt��m
dP{3�x�:`��6�4�����>�Wk��Hg�(P2��~Ay�1���z����bG~��nU�R~O\Y؊X��X��9o��2K)�!9�0\w$�:�B9̕fDb��#|'�W0�3ր�=�����óSg��($�laY6��e��Z,>���3����<o�$EJu��ۈt�"N��������z�q�����pT��Z2:���߃���^�[^<��9Q�@��4��Ũ�:��v6�Dlu�f�9�t���~���� 7���IKl��눥��+����J��s^���o�cQC�E�൸��p/e��(��[���<�KT!�L��^p"i��8�DyJ�V�N�ᶰ�qX[at9�,e]��{Q�v�����WvB#��n_
K��L��5F�K��IsJ�ōh�ݮ��B�/\�Y�m�E����AB-���NG �\QL������4 �����r�D����d�(F� [dPr�6���rlAn��S��f�����T��s�����ˣɹ�(���_UȐpj��RE}M�7v�M&orb�gd	�ܹ;���t|�Z�o������!NaEj�wC�H�5���p4��S#8T7���g �ц)��7B��-�}���N�o���^�勊P9�^<��Ԣ�n�c�҇���:?�xwlB��(�c�H���IJ[�LD LK c�z��K�7~�YV�0�\hPIX� ��#=\�����]fO��'��*W�sw\*9eu��"��ԍ�bG��n>���B��a�m:gK2~�ac��7�KP�Wl�K��\n0�vwG�d���qr�1�e[�$����o$��a��-FȀWV=��0�un�HF�k'=H ˢ⨸�^�Wۍ+�!�X���1٧K�_���+^��dx�~�8�d��T�+�������a���7*!��ޏI ���0��l��(��<9\�uS!��W��D�&�5��**���wv��R�R���a���������0R���:�ONU���W�:���V+�0�}2Ma:����,Z
�%T�M�G*���4�ɼ��:�I��C�6����[�Q'����DS�>�'m�C]�_�P��c��A���P0�Z�0h���s��B�v�<�0������R�﮸;l*���	���|�O:+(~��>v�6h�y����	�ꌉy��QA3��Ju�?��p�q��CZ*�aO��Ȏ�O�i��Bd�Ʀ� �XD|������ 1�=6:vJj9�4*��x���:�}�u
k���ň*��LYB�ӱ�F ��/ ��/x�`�T���N4�:�o�y'�|�1] ������V��|����F��M�ඨݐ��Ǚ�M�	$L��U�Ϲ��ޫ,��E���h~
t�j�ч�]�y�p���9���R���!M懴^��:�w�P�ml03,�x3�_�b-�I�&���W>Á��3�%�I�#@����*��A��yLoV�~5���-��wv���<{�1r�J�{�J��r\UZ��i�����)?I=a�U�b������\��O���U:�Ǻ�6�����a(*U���w&�=��?��2H�P��Ǉ�kJ�A�7u���.���:D�akA]�qV��N~c6��Ӏ+m��}�M飇�h|��"U��ۥ�C���j�z<�͓���f�t�s�u����h���I��p�Ie݇�v`�R`��u�RR8�l\��W���𤱛f��G]��yj���`�}��Dϸ�C` ����}"��n�v��b �TLf�\n\�2�x���g��Կ�fC^8@$�N0 ��+�.&���4GJJ�2�_���
�[�����'�ow�#�,J�f���S���ϼ�h���yq6��+�&��6Z�򾮲x��>���V@���T$-p2�@I���4�����:�#k����5�| U�y�q�!> Eq3�TN��.���z.�z�UZ�Q3L�� (�C�Q6�~q�5�M�|IH.~;��!��c�G�O�帎�2�<�>&�u8GLDY��dA���������<YP-@2X ێw`=(OPp���=VM�8@#k�
���h ��`%���t����j5���tr������gY�P��J��5������l��,�:���vt�H[;��D:��F"�sO/�"���`�bRǳo��+�u�(����bcX�M�s������E͎�B?�`X��J=�����z�^SlI��L���4V�)�hahίP����'%���Y=�~t�r�RpfJcD�r��/;8W����j�"�` ��VF~��S��N��ns�YT3����#j�G��#�yU�Y(���s�W����J�41a����P���uq�C��V�����w^xb�_�(h��5���Z<D�j�j#T�ŕ�O��s�`.D��$PJ��Ad2��|D�I�O��A��$�ؙ{[�b_%�m#>_�p�������}��vrPG��v羂��4��X���zQ�y�~�8\%���:/��s�T�96p]T��p�#T��S0O�G�8�����<2�7�]v��Id��J\�J2KZєވx����`ƉKqK�P�T����+r4F��Qw|ޟ�ĞK}�2V��"�n$�G�@� �;,t0��q�DfI�RPk���K�]hXfV�mf��@;+��C�a�����Fh4:|W8�O�	��]��s��y��ΰ���/)�&��^�O�-�E�R.�s/ڋ�C�n3���b6�B�	���}3-�
vp�}.k�e4��4Xm^���g=ҵ?���c�i���)�
h�'=��j/;-j`ʤzH&%�6F�K��j�Bt�p�f"����e���s=å|����X��ؓ���IW�ThR�͂� ɲ�T^kf�0���v�/ԧ��m�	<����O*^Uj��#���cu�+����lU�h#���k��9���YC�*
a�Xa��@������ơLw����"��,�3u�����ӷW1�ώr���	��h*'�BE#5�yH��݋ �w+�1�����S=�>bԐ]P����G��� ����<⠺�b�����n\�O��L���nބiw���x���S�P�6V���d͏`J^Z�����ZnZ \�M��g�!����HkN��,�k1lW)����X�����4�׮��̄��a��"M˖ڈ;��*����yb��2�``^h/�㌆m˂rD�Ab�H9vNp6��_�9����[�a�T�hs�=1��JB���:4��կ�'J{k��\S�[�����6���$�QnZ�т��ūp��.N�?�F�V��Ӊ��%��`	i��t����^��I�K�f��<���m�y�&�4�Y�����TS:���EP�]
����jK���ـ�J����ە�IG���޴��Y��%�V�x�Z��V������7�%3��x�a�i�-J)��\�7.���UZU�8�{$sn�	a\�r�b�Ұཱ[/_�TW����}�p4�bGOz���� �fB|B{dH`�$�0��.f>#cF:���e���e_F�ѽUU-���s�?P�P��?˦;#.k�d *���j!7�]J��iDz6��Q��0�_������q��a�>�,�>��I�,����~jH��V��Z�ë�T�W�v��{j��㝗^k�ȅ�U���aԮ�:d�uF��~W����g+
��PN�j!�Y}-Z�<�2�9�+i���*����#����Z�߉�xf����l|<
P�2���+G�J�ɼT�	9;Z H>�PH�0�i0�e]�WݳKa�DDa��/��QQ���K���վ�P�gn� �x2��f��Ӻ����e=��f��'pS�tq��đ�'����k�EDK�J͵# ���>��2�^}��7��V3rd����=����_���a�e�(��g������R��)��8\����3y�;B�9<���߿���{VՍ��ikG�x#Oǹ�vԋ��Ɯ�앧lck	�n9J�2z�};��|�0F�S/	�Y�=I#^~��9K����5٘�Pնa��j�6��$���R�D1��{d�ߺ]���A���yY�6�Z� �8���.Π�?�P"�>��x��{�b����_�	�V���GH��i�.���Ujӥ�ń��{���[�%A����$�������7�J�#D��Η�6,;*�]��<*0�?0ytޙ���ԻB$�EwA�˳����ȗOƖ�����$��k�`5�f���(�*���uؗ�T@i�[K��E��F�۶�o�ҫSO0 ��I�<����{��T_4�����Ѡ���bZn���V萌G���á���UwCX�A^w�>����+���,���A�������`��-��; ea��]߱Цo�MKK�W$�_uO\�������b��vb��2�£"�z�q��H	#�}?�5�̭p{U�³qp�_;&B:!���2��ǻM��Q�_���s4�4.�U��3h�h��}��MWvR�Vii~M(I4��	�AX���L�=j8U�AHQ`�-��b�7EN��~P3vm�R�J��<�w� �n5��/�-�>	|���34ȖȜ&�{�-q�R\��ޗ<Q&T�_a��?=.�o�p�mV�u �v�p`���>�z#�o��Y�qJ��=���2�ݘ���E�	�z��NFEtB�_�	�,b��/�F+��}���̱��{�&� �6O��EC[���a�C�nhal_�;�T_�p�\Q��{�JǱ��o��n]����@��~���D1~��Dd ��pt�+9[Z��gk�Ԃ��y,��s�BlQ�����j� ]kU+x;ҬQ��-Y��HrҀ:B"C�{),_Np�tV+�7�G
���4h���{x�^��i��Ƭ^��	�Qr�,0��?u})of/���gfb�gO+�O�+�$����`���F���؋��#W�(VK@���9p߮��@6����u~h������?����d������8xU��{��{.j�vFo]�;�%	����D�} �Z�k��s�!WRRٺ��J�®-�+̀�.��I�B)���<��=:��>W#�h�E��^F��".n7�1�> m�����q�$�a��%K?4 "�J�.ڴGg��+��>���&��븑�.x�!�KQ����|�$u ����HH1����"~O�pj?��������׆�t�7��F�q\7��_�W�.c՝�A>���ޘ|k�*u���f��gP?nH�Qb�o[��Bf���j
��ي��՘�h�	��K�[�f�F

��v �K�I���ʰK��!����<j>�3@\a6[�fb-�SjQ�7E%3S[z�#�X�+9�uM�Cg+��f��_-&����ק�S���)�d �0$$�w���Ӎ��:i�G|�3x�	g�{�6r%p�u��2�nUpD�U����r����S��T�Azr��\59UG��1���m�U>�#o�o��3�o�D�"�T,�a3%x�Xn��7A���6}W�����=�t-֝C'u{���aOe���!�9��5yh���A�iK,�04�2BL����%���N� 񏁩ѱ��.��O���hv� f��}�)_��Dg���Po+����HQ�4��2����)��2����cV	�1wل�Xbew��a�<[�OQm�4���j�h�d�@CE��إp����'�Z�8
<��yB�qc�.d@�Y`�"� �9��oh�̝-�Yj�����y�&x�E�ݶ���O~�B����1Hx�dz�CV��;�<���Whc��y Fwa��1X���-T�:?\����ε:��L��!R�zg+�w���B�S�H���N8[�>L�]�^\�v���9]*fch;�*��u�$��OU���ccFt��!q ��4d��^�꽴>�+B�h�%�֬j=/=ߴ�a�x�ilƼ��ѯ��I��9x��2!o�랉�K��v Q�WvH�EP�q�'9�uI�m[�P�g��wl�^*��1�oj�s�K�ȟK@�bK��Yr)�[��A��T~��E��U���U��F,n .:;ͬ�.����J�@*���������P���뚂��ج��(�Se�z`���^?+u�
�w�wb�y%ԋ_\��P
>}�1�~�(G��zi���)�ӤI:�+2��4��"��;��H|!�'M��ҧ���D�_p���A~fJ��T�ؤ���g����a~�ӘT�����Ͷ��$���R΃=z-�"*���.����l���|����O�d��CB�;����;/%�Qd��0���˙y5G��m�7��B�L�!�3�CHL.�9�.�L4:�C4��B��%�l��ؔ_�,��B�H�2ILZ�TJ݃簲|�N��KIq[���<�l=uwטVU�]��:�A�C�_v����.�7��\3�0�Ľ)ܦ|o�uNz-"7�o�R"���]v��>�z��m�\Jt�?:�g5{r�|���>�'��pg0����(Զ[�'��Y(Ց�{v�����SK����<s;��D���#vH /c
IT��)���8� ����a�1!�b�]$�~���L>7����,lC8`mcbw�`x�NT��WH� dٺ=S�M�*ǋq��Z�
F%�g�*�Mw�Ω�6�v qZ*�(
��3��X��a�-
J��yᆽ�ǐ����{�3f"�.]�2���y�y.ڜM~�{����u�z0��l	l�z?�����F-�R�`�%v|�+O����V)�3j7�_�����|CY���(ӏp�a�+i���(�*kW` �fa�7z�4{��r�0�&::���Ĝ���l��Q�`���)W$Hڪ#�O��K>ل�nu.W=/�H|�Pi�K'��DA�D���)�a�[!/�m�5���g��@o�㩂�)�!f|`^��*�m�^�3���`��!lx����#���n���4�l��s�[��t�C�a� .9P5�۟�:޼и��0�HU�����'fP]�8bH�Ӯq�4� P����j��b�����w�3���i�����m�i���-,�,�#����=zA6�BS|��s|���4{�{��̀S.t�8���~aN�T���[9�a�]^�ad�F+`�����y�C�����Ƨ@ ZF���d�_ϸ�����@l����p,������#���&�EҢ��W�}��!*/���֬{H]��]r:�[6;�%r�Qx�� ����IԿ�
�sN{�eqzT����C*5�Uw�sl��Qƙ)��N���ЮnUm_�$�Ҩ?�i48����Հ~��6��WqF��� K�h�������wgO�C��=b�� Cf H��0&�<�/%��i��y�����6�l�Ҕ>�V'8YО�#�42x���߰eH�Fwޯ$
4�-�ȅ�ƽ߼&�܇TR��E=)������3؎rқ��ƹ���ʙ_�$*e9Ͽ�Ch���A\��#����~��L�Qg	>�����/���E�m�' F�@3�p��qpx�*�o��V��b�	�x� KU��9���~U��Fs�w�0��X����bO����m+7m��I�̧x�q��<6�-i���F���_�]�CNe8e�!V-Rs{,1V v���=oPF��-�zp���waS�J[��6j�����7�Tx4��E�+���I�7��@ �gq�Ho��T�x�9����}LJ�-�!���s�0��ց��A\�G�Vη&"��K���ѐf)R ��s�m&*yX�t�'L0A�,��u)�9�;�`I��cr�P����URc}�p'�n�e(t�Pk)�Nؾϸ���I� @���5�:�f� ���+�jb��ɋ���-a���AL"~B�ۏ���bf׈Eʐ2���ȷ�G8	��o�!I��o&M�ڼ�����xhgc���[�~��-��'JN�X�8��;}�PzG�V�CM��<�c��&��װ
�+��bʿR	�J�J'��	!�i�/A�M=��� 8�1R��f�x:߾���r�B�).�8���v�~!$r�[������i��Wl҆��Ea��@��g�(K[�&�.Z���UeԪŇ��RQ�)Sc,�?��]�yT&GU(��r��%)s3���g"��T�%���+���p���B0�1_r�eeC�>���6�;!�"�)�#S�s�b�=x�4��|���4f�j�}�#0�~�"N��Q��xw��xU-���qV+�
;�sR["�]�Ϟ�y'��)�%��!H��i
�M%/u%g�,/eM�����̽����e��(�.=r���9�M���A�2�l�<C��������+�#&o�ṓ8���ܽ�yWU6��5EK�Q�Z�d�L8p���?e�UƆ��e��:�
8
%G��+�j�~�a�dE�1�YMC�������[q�S�[�/4��!��1�jI ����h�CQ���W���c�ײ�j�h0�F=yx�!,��+��֓�a3�׍=�o���(�9�I2U��y"�i��;Z�3�/�m\#cۘ�U���dѶ�j|uX<�,���Ql�:_/�g#
�m�;�]�hb�VZ{DB@�L�#�v(��jK�� g=��ز�Y�`�RKh�1��;�r���P��>gb���*88��6��1�SQ�B�ڈf�U���{���|mQ̳M�-p��$a�0KmO���o�ո��n���j� ���f݃��1�=���x��n���_U�}io���$���F5{a���\b'�X¬�8C\D�u�=�~�j(X�*ckg�"\�4�d�Y���=#n�"ٵ<G�Aiqoc���l�Y���֤�%"�W�G��1�m��R�o�#`y��\gJ��
츊F�;��(�����;��N����;��,���&z7#��A�D����&Ԓ��N¸9BI̳" �Ս�bx�%��U!���;�)i����'E�nh�Y1j& qk����_G�!�X���������=��KC��2\�Y؟8�D4���Q�'�����c$��������1��Dv3��F~�I386����[�j���j�AM��v�w���gic
3P�w����#պ3��E�}W�G�L��
Lb���q�UI����U6\_�m��	ܗ�n��r���V-O� ��0����}��v];R����<�9�pUj�G�,'ـ�[�[���7XMȡ:���Mcx6}��^��N�irb�h��˭��Q8�}���Xw��r��
��ü�/��w��Q�ƃ}Mɾ[z{1^&}�Cbx��Ĉ*[���D�!����E�0�:�4�S:�HO �|������"/![�h X1��?��[ح�E��q���%<���QF;v|��Q�YУd�n�Ѯ�(��M��^-c���G� v��ҧ��#��N˚�k��C'����_>(��Ί��R��"����if��V�H~�g9���s�#u�5N~��z��F�	0RT�R9���W&��sȏ��?��Ҝ�ed :5=����`C-Q��2�״'��F��k�)���'Ȇ�`d
ڮ�0��F@��6࿱M���g}{�:�Z�N���.0���!�B�M萇x�%���`�|u�n��2G��.��mt>��Y|�T�8x�~<B�L�ΕaM9/��A��@���Ό`'�94�Z���*c��VL��ҏ;L�|�������I�(���k��GV��F��:�!�I�W6���:<�KJ��d��M9ߛ��ߣC�J�4���&�E� �ք�eN~�o�����W�ǛU%��j�q=$/�n��BT��
߹Q�zNW��p�~Z|�ퟋ\'X4S첮�us��)��`�{��U�R�e
S�h�}&/~>�~����{�*�:z	�"�ŭ#)tڡ��q�K�L��x�p��J�nu%nC~���T��%�#��,�����k¾7��'���{˴�l.p��:ӫ�tWGΛPզ��ͳo����M6Ɩ�κ�Ur�{�"ɔ�ʇD,�6�+�.���`�|0Y!d���ǒD��ۧV!}��~e,�/ɰm��#�"��,z�.}���Dإő���|�
��i���V_a�;��&泻U�U�`��Vr�Y��������iF%%��B�ʳ�_Y�B�*U�{�R��5b�?� Qk���h�懦�١w�BJ�SC\lh�1�J>����� ���Uc�k�%�G�H9e���[Aڻ���Z��C��8�	G�rQ��;P�O��)J�������ab$�C��81:A���m��6*�BR nA���?�y�==�I
{���3��#������Qi1�tQ��c�J�(�G_��	��ӭ��L+u꼌H��-���Nb�GԦ�=��{Ǿ]Z�����!�&�+�!C�F��R0�km�O�(��t��}�Q��S�w������3i��Zvq��O��"�?K��}=۵�
�s0��W����9��iw�WR���(t�A���":.�!<i��.����,����˷��aF�ED�'˩�~
`��������1��k�3t����p�om ��m3�,d/b=��Ԫ ��A��%��#�z��X�k���۟��� K�^�kH��t�o�6�&BO��N���Ja�P��x�����o;�չ���!�>��� ب�=�`��'�]U/rϬr�	�@c�fkx��?^nU;"Ltm�V6�3uc�w+7��4?;�&��*���
�&*vf؀+u���X��mx�qs�X����!�q�:�� #lF�^5[=[KO
܀Z�O����3���=���x�� :#���@^&P�n��F��p%W�>Z�2hT?�%]#�B�r�1Ȣ��+�YG$#_�������yx2�R
`���������L�_Ӓ�@�?%�>{��l�pŀ��[��RY/�1��~�2jA �������� ��QD�$*�i���hY 6�(�z��Nj7�dN�����L��5��@1"]��e}�۞N(�Е�ǧ��f��}��%f�r
��[OLPd��e��Y�<aW~�]t�K �"����Ǔ�K���}��f\Yi�G��dnbq�h�j�jj���:�>>#dS��*:�/[:���y�-�b�.xYpR2/}��w�>�t��L"�&j�"g\N��a������D߄�����WE>�v|:+u��=�&ܿ�E�*ޞ�E�� ~���y�(��<A��`�����"Z��'��q>�Gq�ӫ�.����\'�l�_�7A\��m�UuOx~�x ��B�����r}�y>�QDh:w�[�Iٷ�6L�o��L��!�����F��撥�v��rsl��'�a�}����-���w���8�o�)�δc��*Ajh�v��T0iP�WoG��Q�W�e�̌��}^
Y��MJHSb�Ǐ��z�*&� w^A�&V�$
�I�a���gｉ�m<�E\����r��,�I	��]3����J�ő'����̗qkP�ې��-�;	�,�s�f{ҋ��G���A:�Ԕ��Zm�Ӱ_��Ռ낄�48₃�1�p�z�{�^`��3_���r�Q��a�Stڒ���������_(lL(ф�4�:���?�Z�>�S/e�b
�g�#��i�@�� �lr�8�OK��t����6�R4U�d#��I����½37ɨD'��C�&��'���~�A.Z���TRJ��ԎY�ft�y������f����#-;��#bi}�ۂGo��&�y�(�\�q%N�7	��_�cY+ ���9R1=�/'q�rZ*2C�ɭF7)�b1���D���h~�?a缈�Ũ_��*��}v���K�|+�:�2CX��˽�E>w���ڤ.(>��c�6�a*��o�֘vc�=byɌ��������"!�,z��z�L�Sp���S�|�7�ҟ�=�p9VW۞��D%oO�#X�oՙ:�XrȞ9r�4,��cK�?Fl9�2��7�
3{���+���1�l�,��G4 (҈M���B��{V�׍P�����:��)Hq��!�)�MY� �vh�L6�qS ��̌v��e��3T��I����5��%�V�A;J ��>>3r�RMy�r�"p0�n�U��~2a�(��U6:l�wUF߉��8<�0eg#$�K�@��x9��q{��<�m�Ϣ���*��D��zͨ��_�X�3�.Z*�HTe���0�R��5ҧ�5���6����-;�|5T7?{�3`�]���%�kW�f�,��X7&�1���?��~�y�2ɮ��˓��:�/�k�<o��ϸaM�!C/�����:�Q^�0ZW��aB���L��,�k��@���dM�)��<@�Yh�Cx�������^��'.�{?rD��>B�>$:�]j�_�F%F #�ԡ:��K�89x�ѐ�T�G>*p`���0�5�r���[I,�YE�'�ʍV=�堧�m�a������'n�nX��"��
�xG�����_@.@tͅ���i</�� �[5�-?�e�\�~�81z�eX���ES����BJ��9�dh�p����.$�ѯ��.�G6&����>�F�y;-�, `KGc`����q��! �*3K�FY?�;���V�"�l���|�|�����-��,�)1`�5f���%���W�س�����߼$6��'��-���g�� ��Wˎ���Z�k�5MQ+�d��y)U��S��nY*�p�� ��f�
�!kO��u�J���AkZk3,[����U"�\hR���LrcM�VC/�-���%�� 9���H�#���z;��:|G�8+Ȫ>�v�.�j�|��أ�a�*
^N	��VsX��2�F,[6`m�+'oI9��v�u�]��}�9�m2��
���B�h	�]{�C�����IҌ]�?���׽�vyO3;<DAO�Ķ���OWx��cR?�~R�S_���	��^��/w��9����闰�	|E�]��&-U	
7	r�B�è���h���Ps�7��eҨ*!>
17i��K�s��}6��A�=0�[�Oя=�X0c����kr�|�;f9aɜ�'���FB啬�d H	u�^��+�r7����^5�����r���\��uRh�G5FK5�x����x�c�,�8��q��Ie@��-�|�e`g�l7b��_g��f!?B���e���ͤ�v�� ���鎰�-�p'+:�}�q՞"N(��ڙ֔�H���m����G'���an*j��U
��K��|��%Z����#�2eW}��+��mܬ�x)4���,�:
<pZ��_�ۚ6�ܲ{`=����>#:BD�0����Z�o�v#a2D.���X\� a�r�,{-�ڨ��5�k���11{Q�W�.ut���o���66�7����� z~��Bq����ǔ]�G8YϠ4 �Ca+G���-�����Z���b`L� Ut1�x|��	�SΪ��f�]>���J� �Ҽ\E��n�6����E��t�uD&��ꧬ�Ěn��F��qۀ[�{�����dyv/c��Y�S�7����[���5��h��O�iP�M9M'�y�����s%�H�$1���A��SL����Ll�QXh�!���ў17��E�/�S��KF2�ho勄�'�C�*�ψ����eu��$7e�S?#B��r����
��t�����
�_=~�LP�lP�7l"#F�G�C�0z����k�n���2��x�"/ �C�h���teF�I�*�\�8'�D��
W�'��F'Hﱭ���uY���e��h��{Yd{~s$��B�MT�[x�7yo��Iֱ�M~�0�m��A*`*��^�n��H	���"�z�మ��K�cWe£RJ��:ā�W�Y_�D������Ҕ��|ߜ��W�xI{��� ��D���@`�u d�wV���M7�5g(�>+i�/��@D�/�~�cd1���
c��������_�i�^_�~Y��p�j!?�BԼy�F3� FC*��׫w/�I��]��7Fn�n� 9�X/�@f����Y낧��� ��������'N�bǊ-���E��äͼ�]� P�����r��c|�/B�H��R6����u�֕�E��� 6ħ�7�$4�7zd��HD����&@�M1=�)����d�p���<L���vLO��W�w��g����Un2���q������WS`�|����]�a�x��7/D%�>Uڿ�*R�{��51�5	bi�.&��sd�n��O��nЭ�2��-LC �5Kq?�tr����GnҜ�*�Şj��m�����G�ڂ<�@b>����X�\�ę�A��$3Iѫo��_,�a�o����F� ��/�Ɏ,ۖ��'-��_H�����r�?���	����ɗ�zedS�A��Ig�#��n�|CQ�y��_�LE�+P$7��?��5���x	��-�8��Qg�>���p�5JWDP�x��k�+'幽^��T���6�����1v_�M3\��\�w�������'2��3��/쒛��<�_:�Ff��im�.�ۤ��p��<+�ŅL;��z��ë/	��������×�mFX��{?�W_����+ۥO�<c��ŅRs'��S����)�n4�^�"��2P��HC��O	bQ���F�?����Jd$�
	�a���Βė>�Q�'�[--����o��yZ�
���(tep�A.��)U¬�H�U�۷>6�{��
�{V"+i��5�A�*.���z8�w)A���%��6.�N���0Nw�0�0�W]�,V���G�eH�n��)��I��+n6��K\�X���0��$����/�E('��Z"p�" 6�uJӄ���+����"j`��S+��T���[�Sə��ʐ�J�?|��2��.�����J:��))�$䈶ꨐ.���7��n�"2	�)�*��:E�YWf.�w��i����^QКIԘ����N�఻�V����y�v���%���/y��7&G:����������qz�P�*��u��&$b���;ɩ~�+BXZ��ʢ"Y�dQe/�`SR���ܟ�,����9���O^�0e$Wh�J׈K��i|�9L-��=��<C���~�r2~���±G����[k�r��_����nEīP��*��	�`����Y���qm�p�^�B �߯^B���/Ğg�#��ސt0�Ì��7��k]S'_,gc���p��1D��ً�1;	��-�H%IT���kĂ(Ҧ2^��)��D8<����kG�Y՝��k����38��d>�Ӑ-{��3��fn~M��{NXG!d��!���;�"�jeLC��,���$��2��
@%k����T�k���j�"6^1w���[�%��) )�!Jc�*̉��<��I]+%B³2��g�sx^#������>C��Sv��/�f�e�Zgw��ӆ�AXsҐ�3�Q(��O����B�,������h�b��񑳦0���R+j�c�˝�n�0�]^�����a��� ���tݑ���}̫�)O��K�A�X�1&v����D�ee9A;k����Z#��c���?l��V~	h�V�XTNRu��Q�ʚ�~E�����O�Y�A��˼�_Z�R��*<x?�$)�E��[)K�c;�qۀǤ�3m�w���66�׌H���-G߅�2�m��_��_�rF��B����!�z��J�wԬ�Ҕ���Vy	�]�����r��
M��C*���dHȯd�x���gչ�T���x�t���7V�rז�x��0����
�L��'m�Z�C�����~��`���
�����e��~K�[���B�)���,��`�#o7#ڞj��Kxh�7���	�-���,*����S�f}��H����w��Z(�7�9�·�K�<;�=��W7����L�Z�S1�c�n�&F��@I�2��f��$���U�)X��dѥ�5���N+��_�d�%L@ ���^���͔�O�Ҳ"����1��)�T��*Z�2D/�6�kLW@OUF�����{��M@AP��D���R3��!y���]���x(�v�j��Q����d��a��8qQ�Z���3���;F��G�>����#_����rx����s�	9�'!���C�0)e�h05��B�6�H�B���S��k&��L {������c�㬭�4���qc���I�ۊ�F?�b�!�Q���aV�0Ώ󅸤��gb�������v9۩Y�yx�$G��0;���n���m�e>Yjd������UlL�@%�2�(����>;��lړ�ӓ/�H�[&��2�d�VB�0)6V:õ�f�9M(�-1;2)_���`:���xd��X��'���;�̙%��0�iȄi}�B����s�f��U������ܦ����tZM���̽F��I�����Q짗���K�����j��¡ 0�8�q%ǩ&1����*��/c��D�<�ȧk~�lQ3X�Rʰ]lvY<����;��Vz7��7Ԏ,���$Ԯ��5��#�����F��QdZ�eק���cT���U�J��ݹZ#��	a�������&�[����C9��k�ߣ{I.��0�m�"��Ds��Y���xI�L�E>����̌�)cpG[]h���:B�3Sd�R�쨜uC�d_9(�c[�+Ԭ��;�\��+��H�ѿ=�|S��U��PH�Z$ÖD!�o�l&�4Ł��|x8f�BcP��<7u��lFF3N���&���%o\������0o�]8���C�iش��<���y�\P*��D$N�p����y�3	��^���i��R1ddqxdbY���ʭ�x� ���%�'��vF�¢���.��\��'�z�avT�dЄ�Kl���>�5zF %���X�su��_tC�����n^�� ���C�K<�w��_�A?��_{k��>q�]5� }i�<IV,$���(t��+
zU^3�ȦL�Gtf���	���t~S�N��b���1MsW�{�}��R��g{�Ae"�5�0��'d!�͍��Y ��-������Y5�oM�Xr%2�ۀ5b��2�e, ����%Rq�C�cL�?�1�͙m�vl�S���ټ�$��c��:��
풨���g%��G6k95�-�������A[���ݭ�$����Vs��pzI$/����%�'��vG�p�a�~��mUn��h~�V!,�{^2��.,zh�4��0���wq�%�)�m=�T�@�/k��>lvI=wY%�[
�9LӳUr��5���������PL��O%�D�c�ٗ�r)���� �@�f�/�_z�H���Mx\��nfW%93� ���\�c��́bXk�C'�m"9�
o�>��Nf��|���=�h�`*@�u[ˢ��T��g�2��#Yt���C3L,~����n���?ұ���`Ya�_$��5�il�M|,�����Y�
$'flY�#@X��&�.`�!��{��h���#i&ӽ�#�W'?���5��X�π����dZ��eWvd3�2���D��_=ъ������ck�Έ��O��1V^N�ת�Ո� �����ɀ��Uů#tݰ�|��n(�3�Y�{�v� �"*����d_����|�+������sb�g�G:�.2+�a� T)>qfԼ�\�$�U��J���wNw��2r�]5{�u�l!fn��*�D\�?����{֫Y�E�zG�|�)�U�L�=dkъ��/M@���d%f�U�Bm�E�&��x�#���\��w,l�XXĆ�?�;n��ԅ^i�����p�+��j�fV��ߜ�}�� �9�π�[���u�>�dҿ';Ed�У(N&��"�M �} M�g;&�t.=r���f�[;>/R�c�<f�^5A�D�/�9J�p2�CU*-Ы��4�z�y�O?]�$�t�q
j���X��Z�2�X�En�J�}q}=�d#��/��{��qK�v"XB�6�at�J�]50�y�b��`s�Š�
W��H3�59��F��.9��r�0\X��w�9��Դ��15:�tGח�%����!e�S;_Դ>�W!���8�ԁ*O+�% �e�G�2Ҳ�ԫU�J�"S��͐'?9���x�.��͍���(��N�%�}�K'���4���17�	�����^����
��C֬�α��IP6�˰� �yR���(�W�y$<���+}�9\,Pc� {��i�ϔ�"��?bsB��]ߑ^��*� 4��^���&�d �Ō�I$� `6�0;�Hs�����j����9r]T��q�҈>�ni�Y��O�&+��P���sѺp��h�$l�j=�cBM>�lܸC-����XN�1pɗNj��o�����L~�L]w�<�Sp]�j���W6�wk���/�)N�g�k��ד�Q!��@�N���B�u�R����CO�����	A���z$��0^���*$xY[�sy�)p���8�1ܮF�z��nSi9ꐛ��w�hyO��QR`�Br�b�O��k�Xl���"ĭ1?F���j�'�/���g�T�����Q߷�[����Yߗ���8���'�sg�Ȁ���x6��a��kN!.����\`s��~Rc.g�8Pm{�A��!y,G��o턨5�z6.�>�0W�����@"7��uܵM!�V����*}RJUD����I��G]���M�M��ժ��:��/(fi�5����$F���"pO�5B����B� �W����u�%T���q��5dV����?�!H�d/,�Mul��ȴiA���S�{X"ǜ���Zc�5��I\�cY
$7a�T����.q�!"��+��3��0���b������2u��_�OC��&q3�懐G�\{�B؃96��m�c39mq�!Y����W/p�����F�&���P�
�a��'C���:��� H��6p�*������D�Ta��MʐP2�;>�����WVd��w[ �7�]�-��Q7F�`DR�s�=A�J:p��5,�D�0��䠠��pV,zD~�K�����V ��h�B� ��;@͔�+3p��d���0;���=dT�Q��r�P~�YVu��i���8�t1�iS�f���#�m�a�ȴl'�h"�}�<����+�:�GQyV	�F##�`�$��ҥ��j�3#���~yGސ��;g�v���d��imK=��o�jC71�ı��Wx1�gY�;首R�����_{��ZL�=5�%���Ϝ��9@`O ���72�it�{����5t���$9��H����yl��/;��������[~�i��7�,er*0b ���
����mnqW|g(T���Xs�9]�_c!_�2ʎ	�w4.,L�ä����3�}r+d��:ɞV�7���֋�&�*�����t�s���])���ICkml,�)Yrb� h�0k�̪���_����2����[��5A�1����@ٮ��흅'�S���g��V>����T]w��DK�d��UF��k�@��uD%Q��L_s�ձ5&p�ե[��%V�sU�н˞�ߞ?��u�U%�]{�+�70E�?����Q'o��j{2��o�R��:�I��v�u�ޘ ��9!H�3� ǝ�֘"��V�c��?L��Ȍ��Ҫ�J�A��TT���3��@����C2
5d�3���N�i�p�1*O��N?.s70X\�b��v%�`.�g�#g�l�p9>aH�����^�>�9�����j��w��m4�c�C)C���I���E��$��e�U�9�"�m�j��l
C1���̈́v����!��vX�G��<�����R��&��2�/R?6��N���V���o_=s�,�cRÄ�W[�>9�V�o{B,�ȧ,�!V������i�=2"�T���ãoװ!m:xF���4V�����S-u�{|�(v��3�/L�1�Е�)T;C��J�6���r�WV��"7���4k��Pz� �M�/kZF��r{e��A9."����##8�����*��Q�)��bA��?w�b��(����_(�lb�g�|&��u��c�#cA/,ݒ(8ͦ��
|�2)�v�C�}f`V�B���������ux:? ��F�eXU*�.͢�ב��i�I$�i	��X�
k�{�9q��Y$h�ܰ$K\|ٸ͔�X���w�=ƨ�q���Μ�p�����^A��E��R��;T~J�u�Bp�m���~|�b�⸲���R�� /��tL�
4q�Q(�7#�;���.CؘT�E����A���\?��=�:�q�*�U�m�D<5���d�ۤ2�����vO#
���<�������}���<T�-��k#?�<��?B69���9���hˀ�~M�>rJ�nWS50=)w�VԦu\Oy��ai���T4=È:�j��&74Ӝ���;��y��󼀖�pT�b��?�}���2�0��Ψ�7�
��^ڄ� ��f�t�"����M�ɲ	�Rm��3:IMu��(?o3kF����[+v��ɆK�)�}�ˋ7�q�铇{��$'~��'?��]C�,�Y3 �fCm�&��#��+����1�u�22��S�bq�V��"�ޖ��F�� �;9�6UE�X�7��ަ�"so�f�]"큑���W9�s\�7_�z��_h��ղ��ҌЃ�	=��@d0Ƌ�}Hi�%O�	*��J���ɡ�k��Y
w54��j�Ie��m@f��݃Ͱ�(�锫�3:k�K����1����i8ZJy�#�v-ѱ �<���3��	V�[m�5Z���c�p'�����\q0��q�����3y���!�L�}����N������ba~�	���)�x� b�A���Q����_$�Q�1�}K[,!AeC��C�z���yܞr��<����߭�߸O�Qw��d�S��R1v%�����Ò����:�+z[��p(�y�29�ԾJ2RdzӺd5E�69��U�/+��%��S�w�{w%r*ju�|�Z�N�?�R*�s1�J��j��@���n�I��T��$C.	EyT`r�a�HAu�������Ys0$Jc��(%�0Ħ���r$M=P���n�`c���F�W=<�p���b��4��m��.W0#�k��6CR�=���_eI����,\i�'�Jm�ZêN�^J�JK�D?�Z�ډ;���ŕ���úU��eeO����|��J���#a�"�0' ���" �.ijݲG������cӦ�eMM����A�rk G��ݚ�?Cu8�%i6��G�t"�Ky�cv}���)BX3�e�҄NJ��f����<��pռ�Q��X}�o1��w�B�G1\�8ag�A�\�o�\�7�[�5O��7:"mD�]��˶/@~����OP
�2/���h�Q�$y����|���s��E׻�۳������<���P������+�넭-1TM�-���uX�ϰ���x��V�>���Ϝ㘔o�v�Sk�d
���}�j�Ah�Ë�JD�4�������؊�f:t���nr��D9���X�̋�|��5^�А���Ł��@P�-���=�o<wu�����Ɣ9�l#`[����2%w�W"�r7�բbGFǓ.a��
�;��u����s�z;t�&>�_}�E&HI�f#�X��Rk`U��XI��x��2l�9ƈ�5*�����ԡ+49��'�<sd��yʬ���J3�מ��Y�� �,�e�W�p~#F����ɩ���?vK�(WNV�ZA�,����uꛅ��|օ|��=o o��f��Q/�9#?����W�A�j	8ޣ2�;�e��	�@�GA/����id+7�H_�����/�P��!�� ,?�]����w��U���B�f�e�h�"0#�����@X��#_Sb�=2hV�Z\�4����uf'��K���x�����-!�DNJ�f�%��`�3N���I��f5���#���_8�)��bqb@l]*�(eSٵ{���6�Оc��؜�r���8~�z��Rr�&/�8��'��ƫ �)�EFsS�ݍ���F��ڈOQ�@xz��|xJn�=��|/�$�.�]j\T|�"��.?<�Z�n�^�
`�����b#)QpU�b�I n��ܻ�,�0����.N��J��l��ʖ����Ǣ�sI.��>!�gv�,=���i�6]�5h$a�b�\Q)ٝ��'��������s���	5 ���D�.�Ǜ��@�o_'y����ZK1���#S�|GK��4��4f|��-�
�p@q�pI�ϼ�B#�k2F�V�aQ}�2�	�g��q�5���ų���N�o�_�I�%�z�9��b�	�|����ܞ��~�C����<R��m����OcR�67^�Xt�ZR?�r�d�}">O���u���?3�����Jb��q>>��پ$���{*�5KEwN}MNAvA`s������|/��M�~������o�Un5�]<m)w��l{�����u�;x�T}���J[���DK�L_Ҫ��c���<�!z+:����7���rI�H�^�Jz^�x�0�_��)�2V�8�4}n���=���毄��I�"��:32}όy������H��.�0�C\?�+�cX�;�avt��?�P�x��k�&��'iJ�J@Ҙ�?���͸�]9�թ����j~^N3M!�2��ة +���ll�d�t�.9���އA�]��3��R]!S'�����3�a�:��Q��49�M|C�}�[p���'� ZLh�D@xY��Sj�lY��H�����E�����U@� ����Wn<�8[]��(����J���K/�B.A�x����7 ��|$+� o�����f*��~���>R*���\"������=���B�bG�)��k9�R��A�B:��*HV� ��<	��F�(*�4�$��ló�
�9�A���3{���4��/�B%6���Rs�dɀ�z�k"/��&H]���`��N~P��4���o����6��хsR����;B)���bY>'8�Dz���&�W��Jh���П�t�]^��m�����`�͊TC�2�M��(`��6UJ8C/9?�ve:�*��>,��Dn}砆�� �(-�=0LD�b�%�R3����#��.r���%sWxJ3|⿯nhH(��������+uLk����zot���)�C�iw�����!�E��v�,a�����)-��cy6�D"�+ �s�Y�]I�W]1��rF���Ȋ�r}�"ph4F2�H9�'A<����}6�^�^ \.���c�A#��vǜ��k����V)S3����&��r���|l�j��qȡ<��O��g�N/�{¾ N���J��Oˆ�i �¾�T�C�YV^��?	�!h��V�([��mM�Qr��*<�g�ȇ��q�?AXP�j�k��|_A���,���"j���8�x}e�Kdr]"t��7����4mí! �|4N��å��,���sy���M�Y�kE�ΐ����4�e�l�+h��%���˳���'�Ng=fKYs���N���c����(\d��I &{a�b5��zM�|�NTLe��A7�)Nh ����i�F�K��ϩ��+�"��_��,�cc�w܋eܘBq"<neĕ5�%6���މ)v�C�Sa�X#�<��Z"_U�q@Ӏ��� �hts�_��sɡ�Yh�����>/:ٷ�!p�ǜ3a�}@��h:�79Щn숁�$�F�:m�٘���%C?�n$�J q�?�!�C������I���{kQ]\!��<ڡ����7�|0H�I!��Z�����4��[�s��K3��_Yb�(2���8=g�=Xԝ�#����up
��D��L��_k�ŝ�\��@�r������
�h}�D�ߚ]�*ԋ�������s��#i�O8���XS�'R���[����Q��2�,�MMȖ�O�9�a��TL,Oy�C��;&�xtx8�3[;�|��H�fYF���b��O0�x�h�!d��/�����եTD�lޟ�a������v�Z���g��D1�M��X
���4�V�)io)t���j���Y���7n����{u�	��tC,L�Vd�������rf�u�F��ܗ{��yQ�W�5}?؅���cڻ�G�ʞ����J�#���]�[����g��FZ/�W݀�C����*�[��������zo�s�&�u�sR���&�Y0`���E�`BA�`2<ͲDI
�u0���[�&��J��ѷ�q���.}[L6�o܍�R�!��d8I]������� S�n>�N��X,�e�6��HL�M��Ői>"�,K,2�N�j����LΒ#f���|6��i�YB^���ٰ�p��1�!a7�sAd晛K�@A�j�4m�C̅��~�T9*6G�46�݆��C���פ�uHX