��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+�7;���I8������b�bM�D�czC%3��B{;�德(�����z1V�`Z(�+� ]�{9�+�:p(Ve�B.vvO�*���ߒF�q�I+a2�jV{�*�����V�T3|4p��,s�T�-��6T�[�$��ۇ�p;�~,�#���9��^��ahw��N^f�$����t���`^q:�)8�2++g q�`�X��|I|�*���f��*6a}�p'���и\�����d-mȖ������H/��`���g_e^d�Ƭ֝�MJ�P�Vq�[!U8�^޺�����΋R�p���;d:$�� �1f;Gď�H�8�l����a����s�&��h����u��MG�����2�2��>t�T&X��w����Q�������l��r�n �L���wWm��Z"�l�,��L!/bcG��v�ޥ��I,��լ����V�di�t�C�"|�U�L׍u���=�|�V�m��v��{߸� $����|����$�\/8�m�$�~ �*�T}�y���=l`e1g3�D@�.��X6Q9~��
��N�|Tؖ������݅H�5�
l��B�;�J�)�l���R�iDa�A<�Y˂c����~K,zá:�J:�8��j���93�����[�_�2�'�S��Ё�QA 4 "�����6�a�ۻ���0h�!��V;��RCq���BЧ����a~�g \�<0��T�Eԍ-�"�K�o<�03�+�����=��ܻ��{����Y�-?���x�$S���>��ᨮ��k��q�0�Or�s^l�G/R�<Jm�y	�F[�����5����MDxϮA�@n�}{!y�?t�C9��Mx*�a ����∉�qd���%�~W�},�91eH	ܝ�Z=F�����	��w+������S���ܽ6��h�?q���
���^Rj�n�F��!�,Df�v�)Dh(.�=ο�!�_��idz8rݏ��vf�S[J��^����6B�
۩3��ڷ��{=�����G9�VE�����'&�x�A-�Vi�#`o�u]�{p�̵ߚ���qaŢ���?'�^�UG'@���	
����S/������݆��*\�. ��}��-7�!����h�ʆq6�(

S�������v:�h�OM����i!$c�]_��*��23��F�VnȽ56.�S�<���S]FD��}�&S�X^�d�����P���!\��|�("�/���3��$l���O�6�w��?���4$�bu��i��0�_�$;��\얂��y��4v��T�RR`�u���'TIre��>X��4p��٣�����������b������..l$�||S�׵InDɋ7 ��a;.xxM"��K[�����a��J)ۀ���9t�b���k.,ɋ�+�-��H��R�x����ry�h���Rсm��31x�ӹ,�}��4?�5fi�	p�*��%����V�3���;}vT��?+P��G�����{���������F��*�vO}��S��6��g/��=�5xy4����Q�����"�����{׈ˑF����.�7�~k�����D�ڈډկ�'Ca���y���5�N	㷱C���V�ݙ��N���دi�*��ċ
�� ����}3w.w,��N4�cwL���T��E�ʆ�s,z;�J"\k��M�g��& �[5c^Z�Ju�mRd�� ����5Ǥq�(u �ת�����e<T�����+��	���X"�-l��B�OO��4�����l�1[:?�����䰘�hps��J���r�pV�Cс��~G�t��/���U1)_�̿�
��U�w���hѧ�r	�
�Fy�وr�0�;��Àv��!�Y�INS3�΂qO}z�~<���R>9��@�t��aP(�S7�C��{�9��;8��8*�ԔM�g�T7o@pp�^��n��p&�O*I���3���߁�`�]�6�X�Fwt@����8�Iwq��k !iδ��i���8;����vU#{8�s<���m���\� ��J���(]m�B�y�.876���u�$��~�Qp�&p%��3�J�X�S�
r�y�`b���(���v�څ�Ѽ=��?�g+A�b�c4��YQ��(��i�Z4��� D�?�=2d�8MV���ޛ����A��N#:	�ļ�O����X�ܭ�q@�Mr[P!�`T�&��}��I�a;C�wߨ�& ���K�It�/��)8�dg<ߕ�J�#b�_q֮Cm`t9�˜�2%�qR1"�=/I��J��7n�t�n`��mB��J��4z�9����"��ǎ Ǟp1T��p�^�T�l-������<����a�}7��և�;#.{XNRrm��-���u���9���E �K�7~�^b�P~�U�`Y���gc2���-2|�t`͋���^Q�D�pBP��m�i�㙩�!�>�ʹ/+��n[��A���7�ɩ�|�W�b-��i���V�BD�H��Kk�O:o��&P�
�;�:��m�(q�������p!�/�@$h�Q\N�N�odI#�����C]����"8�@� ����L�7n�s�R��P�U|)!�k������*4W�Z�y����l��<K��.sm4ٛ���?T8�`�4�@
΢���M�����KG�>���=�:0"x�$���;{��d� �9ag������k8�k#��r�1��#2�Nv�b�Ӆ*�����+�ؔ�U�ٲn'��2�4F�g��`2�<��o�G�o�