��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�������֦�P��g1�4�q\�v
�`��r�T��E�����˒�a��g�0��nYO#,S$��nd��U����%�������C^⧰��s�z��`���kX]$"�aUs>��E� ��I rP�%Ϫ����+s4���%З�P�ەKx����nyxyHrO~�-|GI�@�f�"ڎ;��i��ca��f��E��h����X#�=�a?>���mK="9�'�qZWC��>�T*��M��c�F�d�A��j�M$�Ĥ5W���Xb��;�\^.����b޳�C�cӈ�����}��;�;� (R#����.G�*y6����{2Q)����
CGAX����p;M��v|�?��b�0��ز��,W�js����N���)��Bc9c�X�R�A���d?`��`�������	gC6w����ci@˘qġ�X��߬S�s�O�a ��x�e��(؆�'
6�p܀�a��v��r����f����5�)ޛ�Z����4ҷ�v}��m�O��:h�7��	�I�Go}�O��c�8��W6�6n3uȾ�q+�y�@���IN���7�H��S**���·���å�%H�W�j]N��M($.ݦ��&[(��@j���ʏ��;�Ĳ)U��.ֿ��5�+b iD�q����@<Ȱt�>[���l|��Xx"�;F�d�/�T1���
�.o�z�D^d�$�*+po�xs�{k����| Vzx2�8�J�r�ڥ&3&�<MKiI:�c�߫�����~x��M7�8�'f���7����M�=�B��8����q�#��6�Y��o�V�C#ub��"=���,t��?���	3�m��gYĒʑ�%��8�ɘ^�ߥ�M(ӻ&���9�qq�(�P.W]RE������Lw���l���54K��̤��ہ��R�蠆�ln�������er�~�
7���]�6�8�lۆ�inE���!�8f�
^ ��r5� ��@��5��ܟa����Wyv���]�����u�%��	���$��##�/dL�e5yD��Bf-X��*���Ͳ�>��3��/�ʉ��5Bz+uw�("jD%�s�nj���`��30�c�C�R*{j��d�2�/g�~'F�����nN�Hȼ�Պy�|g�0,�P�D¾��eVl̃��@r^+�P�/�+�ʡxǐ�b�b���6����)���/挡���S �
��uެKr�z���}�*4`�-� @�=��R��G�^�� ���"�c�,�D�=$t�m$�_c��_�au��
c��.٭�=�����t�[؊��[?�L��5���P_!��w�/��Z���&hIڌ^~l�7���������nO����r9�[�NWs�A��0?�� �{��/V�h�҉�nu��B��*�0{y<h7w)�)�t^�����5��g��	��[Vݰ��5�0@�s�k�]���B@g���!nA!�&�5_����#�(��+m���o+�q�$�rh�ڦ��}����\�<�*A��S��/�
 �f�{����2��,MJ;I��"(�_aȪ�W�A�ϰh�[�K{�^~Ax�s?��F�g2
!=��;9h��e�a���A����g���b�HX$f;��s+N����͞j�ܩ����1Pa1X�=ٚ�\���{)B���m�A��������1�.�L�#Le�xw�i��5��*A<��<'g�U��\s ���]P�v^�^�X��I�������\!���#�P�܂L���Kv�H$�`qɬ���Zy�pDa�f����P61(>��k��}�ĔW֎P��j��Ê[9�?�f��C���+}{���A��|b�	����=���t�ܭ&"rX�B��1Ñ����N��y�Al@�tzs0��O�f�]��Q�zR�Tj�6���*�mP�S�Y��սͫsD�����&"d�7
 :db?�'�{J��M`t:ޝ�tZ�;��qtuk@�$�:̚�#'k��T�2ㄥD���jo��9j��^l��������RPb���ʊA93Y�q�Z*��j��T���)򡧇� �� �$�KʯZ�~:���ܦ��k�����d}px�Fq�0*y�ZTq���#4��j��<�~D� Y�x�R{d?�m�� <�m���R�!�!D���,ɉ��9v9��G�ͯ���ߔ��R��;zVB�r-N�B}�k1m��k�D�p?��c�WL�]��k����&(�y�,����`�4a4>N��J�ӯ�����C��g*�Lkg�1���y�p�P��L�E;a�ȏ�˻��TN{"�|��Bz�!H���*��|�A��MD�D'���p�j;mڬ?MZjMz2d���V��q��Av�0Y9��l���/������0*�t=k[BzS�2{b<�KlǗF��%����$��T�!O+�A��4���`��4n~���#��K�m�<��#'n�P��ㅪu�'N�p
D��n_#�a$�ɜ�V.�'���x�@�O�6`V�4��JSQ��N�ts<��#ߧ�]�9�(l���2�>a��J��W�����4�e�| RTߜ[�ߎ:��1P	z&:��-���z~�j��wP���7k�k�����5�����I�Kx��n��\D�|36�mrgY4�fڥc�כe�]��?���q0�.Mt����|43�I�/��Kñ��N����\��o�`%E�ϫ�M0٣l!����W�j�����B=�R5/�k<���}�P;�R�����m������i�g
hܥ���ƚ���2{����� &)�E���Ն���ݧ̭�+\��̄�d��v�\���XFn��%��[���j���cܣ���m�С�Ů�Y�
���s	��I��Ɠ޴#��zùm�O���bTz�|�w�0����������r�C|YQ����x��S�I�~��p](�=�K ��q�~��L�U�"��QFHE�D����A������<~�8K5]�:0�ojҒNd�#p�;I]�R���A��iZxq��_3r�g�j��;-�d�6����{4ӏ��Q��Ά}��%Ғe�Sa,�z�)w^F�s����usn(�ySĵ���=�Ȭ׀�|���=�3^�T� ���Z"Lh�U	����L�6:����ye�|� ���i|��:X⪻��	K �{�N�RN��誼�;��`�$Zk�<�Q֔`)*�IB@,�v�WW��e:+/`1�-�K�@LQ�zR�W
|`K��Ǖ.(��7���$��:IR,���wo�j�����i�ʪB�c�@)�,/X�c�@i0a/���?|���&����H�剰�ډ��85>�nK�mDA�W��֭'i�^��V�p��\�g�
�����5DڷYN`�%tb�e�?�Ǝ0V���N#�'���S5��|}�{��^�y֮��S��[����t?��hb�t
��Z����!��U�rTB�L�lT4����X��N�'�MT<��A�7H7?��+O0�l�C0���~�,����c��-� j�
?���t���T�4�t	�툶A���>SMyZ#|+��������)i. ؠ��r@'����d���Y��YmE�A�K���*��t����ƒ���)�I�����G�V�����DDM�'�g�߰���o����T���jX�%]���v����%QN�q�Jai��C��Ҋ/vn.P�.Hs����"Q8ɟ�#��4pPp� >+C��)�,����	#[PO�ÉU�ͯ�m(aM���l|��0����|�,��qk��/��^��� o���n��1xBҒm'A�3�&�k�`����`yr}��_x./����Ơ�onׂ�⁷�����s���u9���2#jv+jEޮ/�ի����ƭ�&F��n�w�$)���BZ�+��`h�R4�]
�#ؓB #���8]o��5/���*�\W��p����#h�,EK��mr&��iNJ�Z�����=�H��}Wx��O�:c΂=�Zk���[�d��.ͻ3M�j:[�w��'Ξ	";��ǂ@XXu~�z,>E=��14�x�f�+��]�YE� �L�uEg�H�S��s�j�Z�B�4u��cz�.���i0YJ<�6A�;K�N2�""�k;�����-Ie����X��M4^���w4T`�����,�M+^z��b����WF�r7�Ue?U��@3���a�7�"<?Wֺ����>w� z����2�J�%H�b\F��XW����'�V�Moi �ݴ@=�P4e����X-[%�A���:�f��}�#��-~�#B���_2�-|K�9-�Q٩Wd��$�kHy?1��Y��!�6�Bpp����,�%v��\p����d��{}�M��YM<m��b0�\���S�{�h�#lν�yc���7,���u�F���G�==�Rk���m՘;n@�o!���Ƴ:��A�'��!�������:�P�V�,���J�W�"� c���
��3M=!��/������n|���*�{��'`�ͦ���=]�%~�;6A�蛙�V��^3إg-�`��Z��(r	TCUK�\zR���,�y�=�q�x���ې*��0�k��ʋ���)��I���O�\d'U11���*��"���dn�I�xz�0u������]O��� +P����;����/��wn�6ե�9�	��|��
Ku��f� ��=RV77.|��e��ST>L`dF�E�,�l)w4����@Q2�{��������̢q�Qx=�4�n	�@�@�w���s�bݣ���w�� �bck_ؗ�h�煾M4�mU\X@W��m�SX�
X���g���0�����ס�xg�P
5�.s�^
��ɒ8X*���/�k�|�"����F@����8캑 ��ec<L�*6�D� �BS>�Ѷ�`�l��z9r�g�h)�7ӽ�(�&���q�嘬��HU{c+va�[��>�R6_:ŉ�>��t� a��X?�9���k�E}1e� QH��)�{#r��ŀ["�����e�#��M.�����H�S	�JE���&�[eu����%"��>����f��b�w�[I�2@w�$y�G�N��|���m�~�h��Z��Y�v�k-��v��}XSH�|N�(?�
!����S	h�FW��H�'�-P} @0���y=) |�=0l�>]�2Z��G�^���z�s�8�^�5�}�
86��a}!��4�f�g�dﴪ��̨u�
�z�7�$F�)3��j8��֠ �ma���MH8ɲ�xZ�K�Y{vÀ�1��m豿S[�_[.K�o�;��!�oB!�3�I{�ȕ�d���E�E|�HhP��>*�,�J?|j{F 7��gp�6��8�:�b4ߥ���I��PB�E�F�NA�d�[����o��/�=�W[�Of�z�]�Y�w��mk[����GM���c��1�e>r�k;&�d�_��1T؛C/����}�׺�P���ne�g:�">j'0���K���Ģ�υ�z(5�w@w��-�n�UD`A0�ͻJZȣ���V�t��*��$i�R�>AB�8*R��>4��VX�'$�\J��,�+DM���ԏ��a5;X)"��|H�����JC�q����9O$����PE���I���6)����H�GblmM�Q�,�b%��{'!H2	B��.g����qW���u�j\�q Z��x2/Û�X+��w�-?8��r����7VKm^X���[-#ׯ�0�������b!�b��0yg$W`���	o���`���S.�$\��j�݁������a��8sZ~���h�+7T�%X֙��ڎ��N��)�� �C7t�o����yt]e��#怪��+�M�=Ύ��6��86�H�r�_��f��2��/3}����K�u�j5Y���Ю�!�$���;�M��zW;-јR̎��JD���GË��<�S%�Q �2]8��U8!J�&^���u=�&�M8��<�����p�q�|S��<����)�a�0Q��t�I�Yـ���n@��p��>a�>�(�¯b�_��A��F8��7�3�1�!H2VZ�9w�w�1j�u枓a�Z�}�Nm�}���f����K�j&b�y_TӰ�'p�Er�CO	E��	v��~����>�g��t$l���C�8�����,i�C��b�&d����a�2�������^�|aN�R��46;��%x/]
z�b�>�SW�"��¹�'p�f���@*�^���2C3�!�r��x�T�����	���	�����A���a��r�ELߵ��ķ?�G}��zXEۓ��h;�~OՈt��r�9��]�N�:v~�.��������>2�2,N E�֐t���T\�|3!~��� ���ȈJW�6�+,�6���~���Wa�[����o�F���]�$��S!��h�9/Ʈ �W�h���0Xq7�ޢW��[���D�}�6.�'��柽a������`*a�Q��i �4����l	�0q@�rxB���Ϣi�S�ήTK���!id�8uʱ~X��E��Q4�?ɴ�?�8<�$Qtf����z3A�2�o*�pʊ��ݡ���!q�4���)/yT�k`J��AXrCr&j��⟧2J��6H�5�~��������Kf^��`�Y�!HEy�#�Ӟ�v�zA�l��}�nfl��zBf�5����Eg�*��� 8/�D!�������k-�
���������&J"+�����0��Z�����amAvӓ�&������������͙��k�؄^=O�Z����
닶�U
�t����q�8�i^��5bU�pw�d��d�T��g�IIg��w�tM.`��x�KJ]Q�P��|�u��_���IZ�=J��"�����f9�`:��8��+���q���Н4e��A��P+Ț&���'�x�h�+�wo.I�3
�W�kC�վ�6�k_�*�.xO�;
=��STЮs�Y�ޥ<'ƀ@7�;�ëD=u�V��#�gD� �+��%�õ[�׵H��-ƫ�Z7K���S���w㏳ґ��������c��u�q�m�J�AW��8�	�	z�����hF�\�Z��.�~˸�:
b(�3���ɦ�[a�~pA�#m��9��P�B��[�)�ћ����(�v�0��߬ h�.Zqp[���l^*H�:vPsjk� OŞ�-��>�SB��j @��S^�w�ڴ-�>�Ӽ�M��#���T�b�Ρ��K/�/^���E�k0w*F?L��+�dK�U����X��{ޱ	�dѝ@�[�^��u�oS���|�w��/e���í�+��NgT�3����N��hd�=`��.��&�6F��:��"�*���J0�|}�<n��6��ªQ��Q�������/tp��[��!��'uy�ܢ&|΄]w@%z]����鑹�N��Ur��3-�7���{4/6NH8�(�62Ѷ?	�����a��LO�H��Ƕ��6Ƃh"�o�%�oAK����n�[9�J���*�. i��$�l�ϰ�lv7���ض~RDo�S�:�xu;N������Ѱ絊2A'd�G�\J�q����
7dij�J��pkc��A���E���ۏ)�~�h�R�E­u�2ָG��.���Wv�.�F��V��5�(>B����l.�?Zs�A]�Y�V��n���P4�A�7�||B׭YO�����L��'��kj��D>4:�F�@7,�"{���)̋��u��"�l萈���}>���Ve;l��;��o���
��%��*�\������ޗ!�ަ����!א¨,&�����Y#���S>�J,� �s�����4d�u_a��Q����������TK����5h7f^�RZ�̈�ґ&���|c�m6�����P�l���tO�����2D�D�>�K�U����3�:��l�KW�u�����Ce�e�eox���(s��.K�`�36v�˶�O��É����3�7�6��t���4KI,�6�H���,��W8�f��9Zw`� ����!��mu�]	i�)��K�im�뒊ӈ���4]���\B��X%S��Z����3+=]�˖�{cV-�����E�n%� ��SHK�|�8�6�+!]@�Lc��eB�y�B��lW��1��	NNeO|dJ&��J���y�%#?��l���~+����g�901=Q>4�$�괳Im���/��M�#�{����疍X�[$��z8�"�Νe�Ș�S8���́4�8jJ֦�c�R�}纵��q�5���.�+�/��Ǡ��ɇ1��w-xjC�<��E(��^���q8�R!ĨO�M���C���.�F���SR���U#����M5ϟ�,�N��ZQ��n��8�f�9^�Ќ�%�gd�}�:��<'�>�8�A氞|R+�{�: �qә��6�X�[��p�A��"��/���Z�Ϗ�d�efHn�Y��q�H���IGk���1T�!�dt�N��a���N(��q�z�v�jf7���~��Zٸ60�`���/�X�ڌ�tp��0�<@��������d�������m��h!*��E�leSH\m�^�:���5y��/��rtX������KCw�m"���AiX��B��R���L� r�z����
�����@LP�HaXf�3+�Qb����������a2~�ቚ�"���}��Fy�m,e6����Gѽ��Z����ۡwO ��_RZ�Rא�|�.n�G�+�R�:.}xF� X�#W~y��h�8lZ��*�ț����W����r���er�@���u8?@�����.W�7�T���f]�G�-��(� '�_{D��@
��ۡ�-�� ��<��p�t�~�D
��0®SWs̓��}�8�v���3�/��]_��Y���L/
��b