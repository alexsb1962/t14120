��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������U�#R��D�L��G'ȡb���-��XR%���[�!
k��r�U��7�I�{�5�|� o"͍�g搔�v�{����Y�6�""L�o-m��]#�;�4mߝ��Z?�� �R��ː��^���-?�Ȁ1��/�)-��,����<�R��)���J�\%La����v��{Y�����p�p^�^���ہӀDY������
���/〶����ny�O���O��Q�m���W��B���u��r�Yd�oh��	���Z>�<R^�Ͳ1��޺�z�[��V��L$4��K�ͳ�S����nmx��=p$�s<��8��׈��6�%ϔ��|����o��?��DP&�P�>ۜ�8�g�]P��N-n�y%�k�	���,s�+�Y�)X Ե����x�iz�r�K��/+�*�Fo�0����4��D^>!R��.�Kwt�C?C��J¦������${���MR����y�-�j��t�&��s3lV�)h���Ek��
��i c�*�c��Z�ZS��KYd�a�ûh
Х��VQ|��#J6#�]>�=����nV2���$Ҩ�)��5���.���"R�{�|���+N��^À f�ǈ�]/QG�hƿn �S���	+�a�e�Wl��7/�2��"Ԟ�ϧNt,l	�e��x�RYM+�կ�^��]��Dњ�oT*�U��y꠾&�P��B|)O�G�
A�"�� GYD�,؃%3�x��%
"jOEO�y��k�FT�}Y�Pl2�ylE[�~3��a���}T|炙S!_��BB�H�w��.(�����3Xq�ץkC��-��9�	�쓻ZB��M+]����[��:�Z������i��{ ]�L|;T���c�����)I��Ó��:3�b\����0*��P� U,�wm�V9ĥ�16(��V)��8W�4��jJi�$���7�����a�TXCV�r�_@�&�;��-�	s
:����<"&��R��'=��󴥋ۻD�TN�x�C�v׎U;���]�&���	�J��^�+���(jw]��9ȉ�`���v�+ۈ�K�ί���W�AF���3������j��^ڟ���6��,�h���Y�X�(��ڵ�wĦW\�y4�����S� �rN�F�_��e�����텛�	�#�J	V�R���\(�o��X5YWVCE�R�si�T��3�EYo�"~�1����j~l/(�a'#)�=P{����S���O\�\SC?�F�iZ1޳ë�s~�v��q�@:���;�o�R��9�f�d�[%J������Ce	��r�p��0�`��t�m���t�->l�#���C�bq��g&�L͇��~*zu1 a��{.oй䚪��������-���5:����)EH�b�H�����5C��#h%W��a���h8�(���q�B�6�)�;]�]���Ymw�wQ�؋/�2NV�v��(i�hS�5�c�SE�.F$@��p�U�p�4v�gL�Ӵ
�Bx���Re���}`��,�y�:�@�4�>I ��aГ%�?�����/_l�6�T[���hoZ5��N�N֟�"R��/�Ǝ���:ag?S\Vc+>f��EQ�y���R���^�)8|��Ֆ�y�a8
�g߅~(���_��_9}*��	U�*�G��F%a�0�ajoJ�^���PE���Z��}��>��T�r�l1~���~�^�Sy���4��|�4*�9�iX�ƹgJ�S�����J]hBc<���ތ�fMJ��;�0U�\t�W\�ha�v���/X܁�!LQ_j��<;�k�	3o�N��!_[��H>2�r)"c3��f�xͰ��aKCW@&�7:��Mk2e$�o
ء��w~��
�-��?W�����.^�i��<��H��iۄ=��a�Oo�%�րS��i��NZW���z�^�y�L�Et��&�_9�8�^ �c���?�ĳr1B���k�䟙#T��`/�s�~���2wo�[��h,�,�Y)���vݕz�]����v%��x���+���7�m�}g
��$�%���F��O}^#a�ʵ�ͱ�_r�.QM|��du���
5[�%�HA&"�8S8�j*� ��@6����V��%�C��9�@�M�ܴ�ԚV��:r�G8^�@	��jYD�j8b�lm����p>��E��0FE�D�ɬ܊.՞ddc~��=<�r	+�-���6�h(�R>e��66���(���ڒ���x9��8:͜R�cM~�ߜsϙs�lk'?��_�=�`�2��/�_��O��!5y
��ʂ-G������[����&�՘5��@2P!r��{�������yj;�I�6O�+6�-�
g×�%Lﯢ	�|䳩��IZ>w�=Lޯ��]M�Z��lEy.UT� ������as1mG!�];#��{E#��!�>����k���z��63��uvU�|n����%[��C�Ig�Z��#��5i�
�;��G�=_Z)��5�&���A(%�������tw�:R�͞��<�q0�$��pL\�w�z�U7��`|G̓- ���H|[1���I�2&�PIյ�3�E��7�
w�6����~%Y����ߒѸ�*�Fa�탈�+�̅\�~	��������Ů���u-��9)ȵ�I-�0���K#O�}~T����m���˽s�L��dS"Ӻs���BƷ����~�4��ظ>��=� �Sjh�9L��k�WfY(\ƒ�>��2*{�d��o�*W%���c�6D¯B����쓔�v@X#���{#��ʓ���|j����I20Zt�ɶ�%������f
���-���	Cm��~��ǳգ��ծ :�W�V[�y�8���_�Z�T:�Y1��	�#�}�\C)�su�V��,�#ј��3~��܈1q
�?'mx��6��۷����p��Z�W��ڏ1��{KW�@�`M���X��-�ď�Cni(M�Y�M�'[r���[q?}$|�U5R_��������0���v���*�pދ��Ә#(z��)�Ʈ9F�������ë�2�|��� ���?��"���~$b���9^�c�h�,%�����q�;R��k@��)����R���r�?S�ы��.3���Qi�a��(���6�x���$l屖1�$��}g&�����+�Ȕ:��FJi�
��n^���Qu-�r�GjdM�Ar��ݫ�V&v��"�����RA`)��S R6�>e_�&a�(���J_@h��hv� ؤ��)�?�ho	 �HX`�L.���#0�'C;���a5�d��T�I��e����\O�O��Q�8ׂ�٪����T_m��i�l� 
�T�R�_Ե>4T�nC�oۀ&���F����9�A2�0�1�i98�X��Fي8�1��1 �|�J=���0�b|3��m��n��z~��<G�Yv݁��A@�q-y�&��h��G�c[f��Of~�r���|O6�A��a�2~�ѓG��	��Oͥ�4!�%|������=�LAbW��ߓjc�6��!L�ݘp�$9\����/Fbi�?��]�z�wE��. bË����ct�hX -6�j�R�O�\~+�u�eIymyu��A�����C^�+]�I	��~�yI�K���+g�=4���E��$�>�K�3�P�0�%�����B!�_���!NGqv���CDV���y��l��C/?�q�S�DPܳ	1���g���J>�9��{v9{�%\@��[ ���B#��{��B�t�l�äs�_�cɂi#����ޥ@�r,,�R0��a����n6�:��1^���q7F������gϬ�;1^O|e����j{0-1S:��l������[��C��tL!���X���u�*���C�>����K��~���9´M����V�*�_h���P�
c��s��P=��Ԁ����3H;ی��I���7|���ޔ�MC���G�V3�^�K���~�� �Y2�����?Ӳ����JF p���uu��jr�W�FHݾ�O���;��&s��w���ͦ�{w��7k���҃�H�&����=�~`c�?�,6~�U�u��w���v�X�k��U.q1�����-`[�L�R 8H�\]�������蹍m�W*�́�BZ��=4��6i6D���<�'�9F.�a[�Y|>��5Bô�����J0H'�:<ӯ��0�_�ia�b���34��ƪV<z�ĉ�'QW5����z�4f_���"'Ys���?�yj'^���g<#���T���ؓ1��΂2��Z�yC͞?��1��y�Q���.Z���O�����_�����J�Pk;����ji��t:2��(��P.}J���񜅴��8�cBg����ᱩ�j%�s��v��h�[�U!�M��dTW�<k��aa����tJ_�8]¦Y�YϋG�7vc��2[������K��v~֯�0��Ce����]3�%T3���?�'ܼ#4�U��l�kA���Gp�	����qIQ�?���l���4�����I�c��Y�UinŘҸ�n��pV���6����Y���)O�%*�CbbTj����z�2�������S�( ������_tI�tr[V����Pi�b��0fr�?