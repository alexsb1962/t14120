��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~%���4���Bܯ�&�	�������>��C���F��N�6��r,�_ʝ��lq�����L�;.r5��|Pq翄�$����Lq1y���b�� Zk���PIcJ��ɟ#�#�ܘ��A��P@�`����5�,��H���q���0P>#�C�v����U48+��i�@��U���Q�r7<�����-��p�T�w�㋤�6V�UY�"�����y8��N��I(h��@��I;��b����xf���Y��4t�1���q�w��F�'���?0S:�%��UU<�-'�uMcL`�@(4�h��" vvm�p�iL�O��c�GŪ�����R9�䅞��u��j^��I�V��(w�
���ʹ�]/E�׌ay�P_h�n��ZAT�*b�N��0�ӱ���8��Q�����5�8�<��g� .u�\�Uı%��P
��^�ԹN/��Qv+��+��S�|Ð����tYr��H���\a{ʑ�(mH�	�|�Q8[˄:D���:W��(eӰ���ﲥ�C���@7](/���~�E�[���%�����3�WD����.��e?0C��-F�M�2���P]���$���)!�d��}к)���n�MeY��1O���y#~�k8Q`�҂�ěG)Հ ����_�m>M񧒷u,z�:�8��
�I��
�Ͻ��*�f@eTŬ��I���?�����r!�H��M/
<f_���^3M]��d/_��q����	ݭX��PA7eF"���x������W�K�縙C5qgL;��:ű	[0N/7�K����	NT��.�L��V=t�\�WB#[���D��p�
j��W��v]�y@���|�3,�&�1(�csč��J����0(fymk[������|�ƒ72�.�'i6��%��\%[Wq�����<���{�@�k���y{o��� �m�����P �&Y�]�#�5MI�Z�Pr�}�!�tG3ܺ�um�"W�2���z�х�������v��*:S	�/���١�ľX��Ǝ8S2��$Q�EE��mS>���v�b�Dũh�*� ',<�7?��<cs�ӣ�b�U�(�ck��lM6듵C.<��,'�O�VC)��./�.�c��! ��� �#V@a��iɸwW���}���mj,��=��2���?����.�D� ��܉�:Q���~��i���	SIn(��#��3��Z ]�t�^W.̦��[G�lQ5&QS���Y�����皧}o��;q�_�P�g�睞�f�����b�<�1�"�����Y�q�'��q��EAAe=��9�ƞ3.᫇��N@�)�沜|y�A���hZl�_8�8���[�eX��:� ��#CSN<ϼuw�!�bH��m�ר��0�8͠��k���@UC��O�g-hŷWi`�ӓ������QG��}�}�>���8g[e{"��Z���4��Rw��ȼ�8n�u��w�JH���8�[��\ ��_��� �Ez�-� 4ٍg��#J�	�4�����2���FE����!�t��ebE�p!ٶD]���k#�����U�\��[���x�?E�2C��n�	�9�K�)OT`-뎿3��]f��K+�r��1d -9^�^��:��U��7b8�䈵t�
�O�'���s8�J��o7��XsC�80�����vc��E9{>r+s�W��h��J<�����B��.Y��e�.F��b��L_� 5�R���KJ3�>X� Xh�{��O6��C��p̸�A��C������U��=m�w�bx���N�7�'p<zZc&��H��l�p��`��X�f��m�(�t��u�ɧ��TR������4��7%x �v7�r���RR���+�&g��}[��Op�XIգ�Bp�9�)���b�\�?�6��÷�o�Mt%[��y]I!mF�y�ն8�k Xa�(�m�ܶ�D��J��\�<�(���&r�P����O�Zwg�ʪ�AE�Zz�����>% ���+F�����7��G-�o��-�aNy<���T�fP��Y���#bG۶�3O|���~��H/>_�� N��n�l�c&<m��Q�Ұ%W�3�I�evPB4�4βtZ�+�jE��[�8Do��z�ta��/{(�r��		����t�c��9��us�8�h��}�ĉ9�K� ��G���Fd��	�s�;�/�C� �<�
v���!c�'X{OEXx�8�Û»�x�S�})��3�B��7:J��N�J��p��ŷ�4F�:�s	9]KR��U�u�]���l�K�+k�=ߝ���C7��{(�|C�o^;�&�dc��̿&�e�G���ʀ|�*A��5�2߉z^jX�a��'�7��y8\�mwE�pT�A�A���p`[y#x��4SB�f5ɕ����L���/�c�B�=��O�f�
l���r�N�v9�k0a=6&�H���3�O�+���zn5Ǝ~�M�;CA#����X������x�F?:P@�'���L���-����!V�5i��)�(s�o��1��>����$�&���u~��*�Dr����rR���h8R�_�љ��J3m���:ֲ' yC���j U �!�(6�Z8���2�0��L�8�jw<�n���QQNZdIգn����c�P��]�K��x���_��{�h(]�LØek������+��,����� �]Y������H�E�RX��5�A��&�X����X���w!� G:;�8�+�������'�h|3J|�K�:${_�WQ�^3����,���t���E�y��y)1�c��\�%��"���ڊ�e��h�!ק�h��q�u�u�T:x*$��*k����c��9&	�lE�����K�<�*�&3�oJ*���3]�6i��
0�P(�(��3�dQ!�;X�קbz�~��FD2+k�����U���k>%��� ������:����q��bZ��@b|�b-��f�%��5���䖕9��Ԁ��Qr�v���~�5龋-����Kj�Ƚ���u�t��h����K%��[Hy�f�h�7�O9;>H%���!A�_�WPN7����NrC�X����q��h��������7lK�"��)zx��su%c{(~-7���A�/�z��W˥��B�Іy�3��?ާ��r� M*��!+R0q�ئ@ɋ�l,I���Ի[8���<j!�@��W�Ң�:��u�Xڤ�w��e�i�H��GO�j~F�m��/�{]�3�<R��Ȧ��v�]�ZW����e�~�92��XTs�-�<�����R���&�}Q�`���!��
��Mr����:(	�ʉF�E����i�F:�W�q5G�;�S�,���h1y��E�j���R~�@��9\�}#���GSr���~R���?�_^s*��9��\���k>< ��	??����~@r������g��9��rн���xO��g�}�Ŏ9�X��m9ij�t0r���d�W��_������LEbT����2A�.碸��g���N9���|��()X����	�F��Z4X��oJg��'���ɂ�C>sj]
����n$[)9į;���f�)���%c��]di l$qs�,U�G���Я2R+��Z�J5���W}#����&߈OQ�dD�P���1WE�Q/�c�]�͖��:b�qwO���H�C��ȅ�q��g�����PѰ��V�)�;dP'M����˔������7N���3�j&3�q������=�Q�;����`�{�i�,�D�:L�b�~���~��:�P57����� u�nI2��"�k�m��e�h��q煢�p��C�0#����{���v�:*7�,)?����"�Sh�%���t�ْ�?M�5�.X��U�q���(1Jh�Q�W6CO6�-ˑ`���z�L]?��1c����/u ��K��p�Ģ�FF�'�J�X�Uҽ�_7H/��_u�J;xo� ���h�/�6��ܤ�z�:٬Y|�5����*,�oAcG^ ��33��)�߾�o������!���y2��&q�~.�.9��t�0$�%-�������-y<��S~�Eҳ~��}�{&j>(hK�3�N=��N��f!�<0��&vؘS���$��L
xf;�_zPK�~)�z��wXRw�W��R�wE4�Y!̍�K����}��)k(�K�����\K�~�e�= ��%�4)�#l`�ۏ��"�ϱ~pE%�W�$��F	~o_���ʔb��|<���P��ؓ���Cyu�ǥ�]h7-���r��) ����g�l������.����B�C�;$>��p�]3���>��X,�������T}��,��0I<���v����Ե�SE�=9��Zr�!�rL�#�>z`�wh&^�9g�M1E5�g0)��Y>`�-�kNe��O��z�L�	Љ�U~�VVZ@A
y�iE���t���5���rfa9N�دB��G�V��$U�p���M�CO8���Ԗ_��M�4�V
s�zh�6?T4Hq(�o� gbS�>v�f47B��gg�tp����a�������rd/k�#S����[���EX�m�n0�^���ΐ��� R��7^e�m�h�sM](��([=�
��S���͍�����BM��Á���K���pCz�D��7m_db,=݋�g��!d����9��ύ��[��i\ʃR�C�ޑ��;����^,��/ui��#����d&={�.�w/s]:����x6&�~p��]�Z
����F�Ap<O��xF@J��K���;�u�(8 �ֳ�,	l��ė���h[*��>ú��Mw���9�n��"���1�i��@�&��r�Gn�����L�n|r��}�_�7�Vh�:��?D��Lc�̇�6"0�{���΃$�F`��{,GL��n�L�X�T1����N�4�\V��v_�
/��I�,�A �k=�����\GRS���+Vo�D���(R!��Jc � ��a�O�#���)�P@��J!�X�`��
q��'�|4~G�s�/��EA��2>��� ����I�.'ηh�&��;O���-"x���^p�!�\��TSmV��5Vf��[�#uһT' hv�~`D+�w������s;�~k�?@��r)Is�����1�h	���?=�C���J��wR�N�:P1k�/��~�NO!�&BX$&9�Q��نE2� ����UE��$��HH�_ps�7LƇ��o�Qj�.�y��F��`�:�2�lZ��%���
�T�ȕX]�� H��yV=���8�N6J�� ��t �#-~y���h��7�~���k�{u���	~�!�y�}�;phSZ�t��;l~΍ڕ�}���@@!gV�y���m_mO�~���8^�������I����J��6v$���_ݒ�����ho@/�K/�����<]�y��`�~��ޫK�$jQ\g����A�j����e-G�]KD�hg��(BO;2�;���
hS�[�&,�N>5ѯ�\K�<
�ȑ��r��ژM��֖�Z��έ���L7��NH�}��K��}�J���	ƊP$�u���Ҙ �28/B�� �O��%���]$K�L�B$lc
��ֺ��h�1f��Q�qX��;���,��yN�}f�@m�>E=�"���f�=f�t�@�UcڳN�+�ef1�yw흞s�;�>��}�����w�o})��t~\������J������s�$�'�~ɴM;�Q�v� �W�QrY�Ѩ��I��������6�
'�$�<">;xb-�l<��O&4̌����<DM����
�l�J������|�A��L�s1s���n�>5�ӣ����a`>�r&&λ����_Dl�4Ѥs�.D����Z�J���J�Uk|�ҨJ�<1,��P�z�/[d,�E�3��}�d$�1d�տ�h�b��_
 A�`R�n<��Ha-�w̘�+�;��%wG�C����n�`ws�au�\uIC�6�[Cݷ���?���l�=Ǝ��x0�	��[���7_k�s�-��s٘g�}v��|VXAْ+:�����k�b;�$�׋;{���>����U�wtӐ���;׊�w���Z�FAW��K� Kyc�{6+����c�P3-�t�p�88��<yy���+6l�PY�2L����[s���+�I�8����˚)~��ǚ���wD�M�I�<�  ����׵����"
�Z|\`�S�%�~��q��=�_Z��8 S.�bzfKV)�(�&�t���Ol1F�v� 5pPYr�a����v��	��R�u,��F9d�	j�e�� ���T�1�J��4����=o���~�e��V�P����E|q2C�9���rc7 }�=��5��]V'��De������i����b��(��٨�6��ς ?��W����@L��j@���c���d�.��GZ�ᢢ�h�L�>�rw3Ђ=W;=gpX۸?DMpt��b�����/'K�)*� ��lB(ius�k�\�����ZƷ��G�)��G�{���8���+"8č	�D$Կb@��Š�k�$5���s[�0k�hа�	!Q|5D���4���>R������9|���W�P�/�!	����3���4�UL$��YpB32Z�Mt�v�y��GLO*����z�]2��C�=���M({����X�Kt$ƥ���!�c�-l�(��.JU�g��v/Z
��`*���.����;3�S��	�Șﳤ���1@�DO����^�hv�[���R;�ߞ��u�}�1@�#b�Y�I�9�ѵ{@����/�Id���(of;�R�N��sXE�tY�5eZp���+ȭ�I���+�%���}�[�y�7�~��v􂴿��过b�#X˕���!��d�N� ��A�V9DSx"z�L)��z�FЈ=�ܒ
p������x���GA]��YTi�˘�&��;Uty~M=B��#�m��	oޫf���m�7��Z'ڌ5p{#�X��i�?_�đ�@*m��L
�"MSbB%�b��U�BM���n��/WT�*�S4����2��������cO���=d����2�5.�S��(t� �^��BW�2M�� ˟fKU{s��n��J����=�!,7_`K㋮����R�\:R���ږS�^�˗`��!3��^�jq�h�j��p��f�I��G�W�gH�lj�(Y��W4���/z���9�>��U�{�\�ɾ*����)�H����&mo�$\iC�Vcb����2	V����RY�.�s���6.H7N�2~,�KɳTl@Dɰ�.�4���޲W��簐� �qBz�z���VkR¿�,�-1�2P���& ���CБ�o��5�7�mȺ'RI�>�O��*�j�A=�S�(m���M����/�Co�q�<3�x���W�C+Fr��L
��kȄ���:K2�jF\ts H�Q�u���BJ�35�؁����1l�2��J4�����������[�����1wD��(iң⿗dc����"J�'�a��zD�L[�nZG��DWd�E�@�'g�rT��}^8��A��ǂ�y՛�L��v+>� ō�B~r��)��]���R��҃a�JG���#p��$�V���l*��]���u��U�^���=͍���d�H���1,�'�Z����?����qv�@���%V|���2B�����u���I�t�MN�c���������8C���)��_��1I��EV@�
�B�h*���2�����!�A���V�6OٴO���p�w�r8\�a�p7T�X\#|^�"F����9��a!T0���l�&.�Ð^��"su�!	��M��%2(�5x��5qdX��M�t��6��C�v	��͐���ʒ����=B8Z�,tƺ�� �%(}���6��~��xc��,Du����z�z�{A�Gڢ��+� �+u�s"C^���SS��SD��ZAէ���D"����l�Y�_��Ug�#	u�+ �k�(����%F
-��<���t��}f��`�E�.��h!<�U�F�A��+���n�6;���F;{���\��R�({.zr�|&O�������c����G��E�gr�O"3�V�sS���PsWE�����N|�lj2�Ќ�]m�p��� ��w,�a��F�����25����w�B}ke���U\lk�a�f�m���VD�N>e�<V���e�H�(�
8xV�P�k}���/�ɴqK�_�����L�$/q��J�	�s���_��xКk5�+��ќ	�b�P�h��݋�p,/ը�ˑ�
��.uw=�ɤ�[�.Y�[�ub[`�W{Ы5 %Cғ�I�-����Q�aliHP8�R�:&C ���8��eD��L������{�Ř`1�	��)wz�ר��B'�#�5�(�?�&��oz'��T�E�a�u�6��y�	(��9�r ���#�R�����9�K���¿�G���Y6���v��n!:���M�
p�9���e	��OP��n5���;�Tf�5�
�,ҪaC��������!I ƛy�%]yr�;t3t�����d���B6��c��>�]���(��v�{S�#a`��2�ˍ{$�mj�r�PH�c�fʪ������^��h�7DW.H�,�(�B���F`yg���47�vтG�IoV�o1Ѐ��b����Ʃc���̀9�t,�;XZۮ7+P�S��6}J����@3;����B�025��r�4���E�DB
�����($]3D�[�oR�N�o�oS�R�ǿ!��_و��h����_�W�uؤ��;��|��"$y<��Z����z�4���0��v
��9��r��
5,��O�#�S�qp"����kp��Y��zh�^����3���{˪�&�����Q��Q�
ſG���{��C�?��F�IC̖�T.aAפ���s�-���(#�,=-Hf�%��X���)_p2����8hĕ�&9?��5*���R���w�ʐ���E��M�(Ld�B�!�9�QڂI�լܕ�Et	NQ��M|�ْ`�5��*UE��U�ȋ묥��rY�]\믎h
���>L�S�6]C��/�.a�{�Z�����s�MFM�2������\<��C���4A>v|��Q�U5.@�8�G�8��T��ۺ9��2�.��֙�o���{	�1��fW�?;T��n�˙�F�l��[^DU��`��}�i3�XO��J�y<�%�x����g s�S�S����K�q�dNߢ��~��
&��-ٱPâXAv�%�����J�u{R�]�3���ƌ�?�8b��;ҫ`㉛�g4F}�bz�{E���[�.gG�x��A�i��i����4�P�Cl�z�O[4Z�	);z�Kl���xk��ԙ��2Rۻ�c呃|�Kǉ �
�n���Ƣ�B�L�.��9�*��ڀq4 i�hޣ�i��CA�q���t�Yd\����� �	ý�х���*��+�٨O��@j�0$`�ۗ��j�n�7ig�Q�5�ǮF�'��x��;�v!�lq�m�oݿ�n�؟}|�e3��#�H���i�J��i����A��K��xz�Ɋ����#&�!��ug�۵3]5������4	�W�'���h!pݽ���4}�T��4�&��n^,MBj��Jz���6��62g\�b�I{��7w�n��]��=����0N.�� 8w�NE���+d]�{O4x!��c�1�3
�nH�.��ͼ�m=��2�i����Z>�T�m�6ٓ�͖���`���:�S�@�-�XZz�ό�+/���	�H
W]����_������@�f��!��9G��;���&�����ȡ�4�؊�'!�=��0��;�pp�7]�7�X��(.�$!9�R�`�TB甃w��޼�/��nJ�ֺ̼@E+���|��v��ҵ�����|o����+Ӭ�E-�u��V�M�{k��y~f"�?f��76�z&�^�ģAs�&Kp�*�]���%l~���4*)3�b?��F���R$���������-���V�����:�kZ_s��O�E���(�����N�N] ���}�w�����K̈́llv�S6�k��]eJ���	O���n�<ە��.����� cU��SV+l�̤����4	�&!~�A
L���*�=jnu� �H_̭}O1ӎN̃�&�5y|��YE�R.YY̢�XІ��;��>��=���Pȸ1���i_�\�D4�����R�c�2�J�z��f�Y\����`#^%q���0��M~�
%|�l��9���P��`f�����w��y�N���p�A�c.y�
c������Ǌ�)ѯ�8Jz6��0����_��b�c�Zm�Q!��Ic3�ߟN1 �E���I��i�����~�&u̕K�	���V��*k�w��G����5�4@jB������5[�L���`��{�L�}�B
$��G))�moA2fe������ׁ��o��^|~�}�Q��A�~[Ո�*c�/j�+�C�n�f�+��J��l(e�.��WkG��7�Ӟ��h���	]Ç�^�������|�&2^�=��frQ���JR��+ɟOJ�������p�*��a�R�7D�;+��d���Q��2������M"#{!cX��p�H���R�3�[G�x�x��Zs"���ѷ�5]B+�Ő.�1�ȧ���Z1�Њ:~��4q��pẺ}o^�F�s�Ƴ�+,��Q��)�(s����(nP��<p�.���ӍE���2��R���M��7������e���\�$s"��n�����cjc���r˭|ʘ[�hͳHvh���0R��x̮:�� ��/�]�S	K�/���C����u�;X�{�B:}7>�t� �QQ�Y��m�Ʋ#����5�zzLAH�/C.����a�}�ӱ�B��z�p���E�5�c9�OM�	)N�G)(����(�m��{��ۂ�'�zI��f©g �&��E�8���L�ɗ���<�kܪ�^9�K���T��L�� ��g�΃;���C�\³L6����lt}a���i�NU��ej �լ�;`x�M�KX��䉄���GP˃��H�ˑt�����'i�q��
lI�r{K��]t�.�|���`��_A����K��>?Z#M��yip��X�,����Bq	xǼ�O��u���n=fq�f5�w���"~\H��pO�����$dW���o!A�B�!#�P�x�ͼi�oא�b��u�R�a5{��]��%q��
t�Z7MЇ�|�/�"��ʩ͋G������t�0�� ��v�դŚ�*_s����R3�Kq���
O��	�&`i�y��}�QG!i�A1�0&5�L�7�w�����;���[:߁��L�&J�V*�K� u��D�!؎���_df ����o��LQ_����5����i	Gg
�v��$kί�q:�&�Ɗ�֋i����H��X��YHh^��bUM�ΓM��E:�M�0��_u��f��Q9�9
�8��
u$cn].ERpjRL��Q�<�T��BO�S=f�/�u�0���^�H��D:	�Y��>**]��ǁ.],ik���GJ��sd�<E��@mގ��9����������p.2	�8,k�^�:v�� :�^��&;�R���;*pA��#f�Ds�}����&��]zKe�'*��� ���x�{�P.�'�D�t�)qk�xH-F��i&�>��&|���[g�$��W#ř�\_qO`�����h�27;�>D5���\�J#�N��B��!�,7" ��GO�ϓ@;�1��L`��]��f�W"��Z�e����L��5��E'qJ~��	RӨ����Xn�sX��wQH:����+�UV-�O�bq�z�GE:�K.}��1�ߘ3��^x��H��2b�@��pYcCa��dG�V�����S�#Am01}�+bt��գ7z��
w�I�,���6�tցo����8u�eI����e�����2�6�|h�x&f��>�I�۳#�����h#*kw^��O��U+Jf�h��Q�K�w��\�v��[���ϗ���b�S���ó��$TsH�=!�n=�rdL��Jn�Y�f��ܡz����f3t�6j�H�7c�؀���ʎ����ʝ�a�y��*hV�/�E����e�9�>�6�v�h�h/�
�W$�u,R��0ڟ3m>��f��d�۸�?�r��<�lO�$�K���2n�ޓL����H|,R�d��
r�78���t��]� �H,���C�h��:`m�������� (>�[-Q{�$��(�������I�T+�d�#��9S� ��"�sn���K#�ƌ]l��,s�����Mٻ����ƃ�1?����]r�+�@jJVz`R2[O�r�=�,cd͐�=��*y�p�u�Ϛ�H<�!���f}i���F���q

V8�J,'u����H;HX��5^~
�[5�؞gb��Y�������-�p�E�f-�\�<�����*���݀�pM�k�/ª���z���M)�v`�Ã�xY(ר��M��<zR#�a4�
q̾����L!�qUR����p��W�N+mh����fA�����	ܳ�3q��tǦj�+�P��?���)��о�%Ʒ3���y$	�j��b+��sK�d�X�F
��e=	/��%��1hc�����,$���al�&��SE���TFj���9 }g!<0�D���@2�XЅ�"�����}����O��2�Àw�f4#%�q�ӢӜ�g����[���y'�f��l\�<�J���o��)I���ʋ����օA��'�t�?F������o�p;*����;6S�z,S�]!=.0���d���[��a���_a�r0 �^`��oe��A�&��iͺ< �����&����}�&��hE&`.azG�W�Ĳ����#v��rn[#M~ .��J�oY�@t���?[�d݁��ׂh�zHf.b��>�!��܁��S�|��'�sn��W
w��G���a]�4M�Db�a�E���3V�����be�H�(@�%)�Hr�_����~_����^ؤ�r�iy�Xྜ��G*�S�}p��$��Z=�1:w*�Ө�9����P�$�>�kp��jK?��#o�⊸� Z�=p���o�o��J��P����C���$��6IOˌO�$���d������#9�����η^�~��y[�Qғ��vg<'#@T\v��x���˔�@ ��G����ڞ�M���ԗ�X�����O�B�ץ�?O��?�\X5�)PIUl�=��ƒ��4Kܢ@C;Hy����
��iF5�-q��TTn�w�9n~�]U��%��2�@�Pr���8
��3
��+�ʷd����M6��` ��Z',�����n�V�7��=n�!l{-\�Ϙ�(��Rz�����
��4�DL$Su��,(�#HǊȳ�S^���h�
��yT^�e�'����R^%dW�W��\Gc�(�yfF��6�v��u�C@eb�H�`m>�w�b)d�T\�pj��h]H�� Q��\�#?8Ǧ��gZ�r<s����`�ީ`z���v?�1�����V��GIg˵e�3d�<�3M�Z0SNx�YDsbG�p�؏��AOsYK�
^/U�Q�-��q~��=s������#_ 蕁C�O[�� .�f-.���YP���-�ފO��53�׉��>?�m�Y��}L�q�7ɭ�+�I61��͕V:����B`���O� ������zS(�wm����̶�᰸/����L�k�	͂�;6G\�!8� V��*r�$^�n�rm;����>P;f�_B��1	s�Á�	_����S�����������y]~�s9� ]�e�^��N����|g&lo*ڈ1�0���ws<�"��D����9}+�j�����OxoIѹ����e�cU��'�Q���b�0��җ�B�J�!&÷�it��kǺ6�:���'� v��e�Ԇ���U/*���}pV���ۇ����ř�໑)�i�L�1�%w$���>�#7mh/�A�'�
g�L:��[A^mk�,�d�M��uJ�l��#�j��	m/wة�0��C�Մ�Ɏ�i���Ň��>0` �fB�=;I�kAY�-?�C���R�S�Ic�~ނI�ͅ�pRh�B5�Be;����hzƧ���� ��R�#�����1Y��G�0QR�|�����U�H��#0�h�:�;?�&q�q2Uo�*,sϬ��qX�W��+��p�K��)l�l���}n[1�/��W��R�?��du���p�,���>�vo3ҫ:Vf�>Y��m�|�l�׭[X��ʀj�^#:�b�H��[��9y�F;8i󏩳�E��&�1a-�G�X��1�4Y]	�Yѕ\�ʬ�pPã!WU&"	�g��pk䢌�M5>ҎF�Ό|���wxFQ�s_|�x�$O�<���^a3��'l�8P�9%�oۧ���������K*�R�s��7�N��`�HvM����������1�9n�sѝ�0='�N��j��V3{���%���W��<�F���tG���o7/k<C�y�ez��sE�9|J:�p(��ȥl�����Dq)��[?��Z,Y�2����~���@��ø��9��ĶP�Ʋs4{��t�-+��i]0|�Jl�Kq%Yݎ�îl��e#xL��\r[o��Dr�r�^ w:���z�g.���
�ZEE��B���!!�o��s��ٗ�	�M��z2��i'�3�
�Us�yMO������W��o#H�|Qa[9��;io�|8��҅�8�|����F���O����'Gb��dTQHf�7��*��mx�TI�1mUJ�y���>#q3ZW�'�� 7�@�����7ĵ�9J��fs���b6!VN�$�0KݖE|��M��	e�lC�)��;��3����� љ���H���g��[Н�f�!����ʞ�^�h�)�;��BЛ�#��]5������ xbk�*�9ɑM���U�j��B�z��;��׀e��`���0
��9�J�@�h�ݦkp���GP��F����,"wi��4���mY�%���C���檖�AǮA�	�8X�#�y��n&T��Jk���#�+xs*�ӛ�m�,5�7"����Z��Sp�Ŏޔ��<w/�tiY��QC��1+��->�C��DpB�lHB����`�L����W
6��C@�[.����LB�dz�>�Sp�FOz!f�$�/��V��~��	�B�hqRC�P{C=�����ʒ�Hze�3�i�j�ϥ���.SS�u�?�Oa�U�P"��V;�. ��*�](���3ĚJ��ѣ���>\�]u��o7�;<͉�jՍ��7�{���<)������c��'C�*�t_l�*�<X� 9k-�2S�*��5ʱV��n�T���s��!��q��)�'�!P�`uVH��3Es�M�M�����խ�6��hhʪ�.e}��c�S�#�����Ӕx�k4�e�&(�<�?�
ذ��s+V�.��}`�c�"ᐡē�n~���Pǹ��n�S[�,آ��Z��᱘I�#�UV��[C�R�)�C̘m�
��'�j^C-����_��K���G�ėF�E����P�v�K��4���/G����!��z>1fW>	�2e�	b��N�����lf�?���(]�!/�b��^�T̓k*�䥲�P�r�j{�ZMt��/�O)����8�* W�j��PTK@>�g}�Y�8#̠�
Ҩ�(�_i\�̔�=���!�{w��>�dphi3����/#���o����'D�;�^�;G$�M��1Y����P��؆�b �%`��Ɔ@�&�x⧹���"L�_e�E�t@�r5����������I�Q�z	_tΚs!젥N-I���<�����5�2G�M�����S^ub3�$��Ul��\ȩ��J�/L�� �+ﱊ/{��q������c+�i���Z��K��K@�r���Z�.5"pԀv"W�MUb��d�s��6��qEɱ�xY���Л4�I���N1E+��j�5�>��t
e�)�� fCt5�L�Y{��1ig6tg�t`�nQ���j.������D������
JI)�m�h��c�,&dyC�/�,�)��Ej�܇QȏǪ�� RB�d7�b����ԃTX�㜖�J9�^��aKVN8l��j�r�a����>C!�9�s�~6���J[_���������>�Aq	]�q�nP>3��ʷ��*��q/��a���ix�_������7x�t.��H ����#�015�^�SI�:���M��z���Q�l4�hml��D\�W�L�Z����`V�2N��W��9��n�՝rtj?!���R\��]2kHx�% �8��Z���CD����Ug׷_Ѕˤ�&��Y�ŀ�ibd�����t8����� ��1%R�h��+?֦���k�"�㧾���.�mA�2`yI�h��W�W�p��V�Ia� �?�qaU,0=
��N�՟��h�������[<���m����]��F:��#�Y�����mD-V������%t�8�N�9����DG͝[vN4Y�'>���݊C��a�1w�ܛ� y��H!�G�;س� �ؙ7[�|��O�@57i�a����M`}D�K�>�O7��$�¨vl{=Ψ:�������P�o���*����Xg��,5��ql��FM�cG��%P6���枺P�Ɨ�������>R�aSH8!�1�a�b��S���U�%��A�ڲZ��B4o�*�#;�u6�D=C�'"��D��NQ�a_��_,�3�W�Z2B����QX�*޿S�8d�T9��n�E�,��rڈs�T�7���7�=����D��+�'��-j�a�ԍ�z8!���.s����i�К�aº!V�2�}�Iw3i��.�o�0���w��1�L
K�[�Z��P���$|)��	
�W!c˂��q)��R1gзy0u�`��і�w��`4��)�mZ���"�0����)���-�}���M��DA�s��{c�����Љ�[y���=jb��㯄��{#���c�=yɆ$Z��/5�,*~����8*�_?,NӁ��n�W�
��(��>S�J�z�/0��ud�a�L2�;Z��Mѷ:\5b���0`�� ���G��#��Z~體��/9f罪.�p��y~
�9fM4�,���'�7PJb��
�g��ns��Ӓײz����?�c����!qp�"�J�������+U��	��fS����">t��t#i1�f�r�r�Q݂��,��ČSF|�q��t�b�� �d;H��i^N�����yO�����3�o�^�v�(���:�q�4���~�Ɵ.��%�2�M���`W����#tF>��9��͠��6urz��B��yfX>z��-�D�H_m��R�"���(�D�=C������:g�Ȩ3({�.��nK�:�Z�@�L^�I����U� ,&�|���zy��zRdύ�����$�Ft���^
���î�b�b�iB:܅��SZwÕ"��㍒Ts�O�!����=�&'�`�Rz*m�q��
-)�$
u]�?:��{7�e�oa�VR����;юH���h6Wh�80V��f�Y+U�YF����`>G�y 䫒b�x��u�-N��5�1�ũ�ƈ2ꓞ�`*����ɛib��O�w�%��!�� M
�kב�[鋻>��$����֕�Z��ǎ�1�k�8�JBz3���b!�2Ci= "�,Y�s��Thq'������͘�nn�g��W��=Kn�; �7�I���==kh?̏\ �Q��!�����=���!��Uz0�A =#�u��t����J�B�o`���P� !y�����c���d�pO��rx���Sx���Q��>�����٫r���9\K�c�71v�f������Fd����汈^S<�OuG�}FRE!?�C�|l�g�'����9�y�9��%6-2B��*�F�zi�@���b"���]GI�<�_��18LҠ��t����N��l,D��R]e S��]�IE�5d
�`gT�r����0����! ޵�����:Raj���/Ȟ�y����S0�ҕ�B#���#'��}�>�K�5���AQ�	" ���8�6��u�ͻw��� �m^MUu��p��YB9S�J���TYo��s����Ԙ�v��T��8g}�Wy�ek!���'5&��PF8ǲ-'_�1�8v�Fl�i�~�Ӟ�����9ǈO�ѕe�����G�Q:���q��MD�BS׶�*A�[�/�I5�N���*�~KQ�FPѡe6u����A˘��DÂ=Mo��������Y���@E�h�!��J��1MKm�.l��J��Aˬ�4�8"M�h�c���܎o@�\DI�Y<eD+�ey_Ź�n��X�| <�ѡ�V��e�K�w�B\���g�ؑuQ�by�(\t�(GN�c��¿���1�����,9w�6�P��'K��;Y}t���C|��$-�n��	��3�����8���$m�E�F.��r�m]���J{$�=N�4�4q��7����I*���U���:`�B�� �������|�9L�- �֪4��;�nu�4���~���5��U�_s�]�-��
��t�P����V�D�%���Bd1l#���haJ7�� $^f"�;��n[J���}�	\^�0'����5UO^(���K��=�z"k����ܥ���9+)[Y�	�"�SadX����W�Q%������8wm��sF�6��!)�Ǥz�n��sb�z��	�J.��03��)�>�k-
S!���G��b��+f����0�Lx`��M�>3�x���Q�;Nj(��SIhQQ�]%����,É��Tb�!S!m���]#��V[����go����U��5�S����}G˦����n�H?qQ����_IQ�
[�]	��c8{y�~�ɷ���2�'�6
%�g��(�n9���)4'���9E�Ӳ?���c�:��u\﵌��&>�0x�����	�=$��}�#\��SAbA����-�R���ƶs@��e��-8�x鎜YT��xq�iܒ0�@N�ޔ-W>�����-`z&� y�Ƒ�_aM'w��z������ �֥W�Dj֙	�
#�)���b���(?�Z�\K��z�����Lk��ň?'S�zb�^80���j\�@B�y�Y{����U�1rFެ�^���e�6���[~رlAF��.���Dq��kVK����]��R�!��p~s6�oNz�Jhu���4c��,����K팜��k ��+����w+[e؎Z�S�w�*+<�[x���3T����d69�	�!���a�9w���J��h���5=5����L�'qqx���@ý��D��?΍3?��M��w;~��E0nh���-Aa�bུ���K<���z ��}-��?�1s�.�`2�k�O;�i)�o�C��ϡ�&����?�b��r�@��9��4� ��%0	M��Р#J^��		��q��KM�J�ဇ�<��>�`Cn��������#Ƙ>b�R�X(�D$y�w��f(Y�p޷�.�������_<l�W�~a�`�؅�/�Q���0]t@��4��p�BO��Є�C�h����O�F>	�|%iOѤ������i�<D�+���n��L|\�$ڑ���5v�!�e��6A�b��<�f�򍑄���_�Tg��A�
�}!xƶ�؈�'�aD��������А�(��P�L�g_(�xV����� H�oK)U��^k=WSv@ۂ��K��P�LǗ�Ί'�/9�.J\↯�����i�[�B�w!�iAkfv+�9������nn��H9�Q� ~N��ƛ���xc!��PD�q�	�m��:mF��������9���=5k�s!%���X��,�L:%%�7ŧ9��H�̼zf��گ��()"��EQF��iV�4!󒡈P�SA`R5@�(����v꽄BqDCkN�~�����ݛp��R��d�N8���c*1�^�,l�u:�Qs�Ct�����ط�2��q��n��\4p��d{�&�W�)�/U-�bb�+��Դ�+%���K��u�,A��˰��`���qg�OS��f���v&���M����Rg�#>�"��~�3��.��!�+������ΧaxOԨ��Al�7!���r�-�N�p�1�K$~��ĺ&�)l��f���s먯�ҷZ��|����ɧ���V")F�5��G[i�<�f1����+y�YI�b����N� Tၮ×�f7��8�E	ܯ�7��m;LF��{R�"2]��X�8�M���H���I����e����
��3��m��)>2�*^�L����2w-����>�Kc�־���X&�N���6k�{J�8�U�r�l2>}$w�Ż�i0�{|�t�E�"6$��
���H��Qb�O�n��$_柗��V�s��/r!F#�tǏ�+;�"�>�wǕ�a�:�A<1�nb:�B�9THX.�����w�6^�(C5�s�F�[z�	������C��	&�nN-4b(�� ,����񜉻)8��8�/+�9r���|����Pj�X��8u��ǿV�S/���:��4S�Tvo�:��o�yLki��L�b*�.�̓T���41H�@�A�f�o�u1��l-r���_�WL�`��n"H
�y�����5"W�������OLr��N T"��t�U���d�DP��eDi0��H�(_EH:��uX�&����HO��G��*��*Z��V#bk��~_�#��i-��c�!�=�r�!������[M[���+Qq��Ix$���`���?�Ky��Fo���X�$D@ĭy]<�O��N��'�1>btE}I+y@ُ\O�`�׈ ��m���A?"!PvޑؕG��!])��I2�Q9$����]TXG��7㱶� mD�c�x52�M�X����4����'���S�^�,L�ɫ�q43ˬ���v$en|m���NZ�o1���B���H�dZ��{����a�YXe�p�L�� ���� ��GWu��1�ss� � n+<�۲��Uw8���!�A���8�F�O�%�M�������ހ�[^�J�j��q.SqO����h?���6��Yg����T�����LI)�Dtm�h.
;*�g�-H��0Ca멀D�Gܚ�\R\�D��y9i�B��xSը+���w��U����"�wnR��)n�ˈ�;�4�b�ZB�"e����\O`����$4�4O����;����i�n��t?�R--/��i�����G��܅<@c��+��a�
���M7���A��N��U=s�ޏ.M�V��űG�9��%�_�.�u���y���)1SU(��se$vv��ى�r�9g��*�@N��7�M¡O��M��(/�}|�=Q	D��53s��+��;3ܦ�y��g �Uec�Ob����O�>�H�YF�?�������\�([���e����y�$�4�t�)g��U?��x.�sc��U�N����=�S)@�W��N���ߊf�]�Ush u���n�d����;w[`;BdzE�������
v͕JDyq���$4�>���U}y��=stVc��¬׼����R�]��8+g%���A��af5���}����2-��vx�A�C5t��:ӤH8��v.lT$G�� |+�p�����_�, ��<�)z��-�m�S/8ް�x�+{��~�3J~��RX��(��l&4�D$�D�U*�x5hc�mq�X!�x�h�!¡��w��N
���5�q{&5
g� Dvق���j�؅Kr��ch�vB^��|���t�	�EV���]M?�g�$���V��cC��l^s$T�5$��\��A3���Kg
�M�ɶ�P��\Ҝ(y�+9�z7C߄(����Ө���/��?�6E��k�������
���~})gA���sw��o�E&�dIe��r���(�`��:�㡹CB�	�Rʱ�&є9�{�̊� �����l)�gt q˄�íC'�_C`.B�d��g�r�_Rl���CcI_�_Jy��Վ=���V�#��}\�s�V��x�3�;���N��w�ye����{vnu�BY~��خ�^����tRƑI w�J��FhH�~߈�}ı%�u�Ɖ���[��F���8;��%��4��o�E]�َ/Fl� �b>�?!,2`�x����d'����T�����H�0*ӆe����1�?�j����ת���K��)�aY
j��a.�ht��X��R[�s<>��L��M��~�Y�88������9��t:�p!��Vơ!��t}�yS01f]9�5���;��f����C��޹B��x��,��lN/?�`�X��+㗩�+v(l���w�#�ྲ=0o�>������dq�%#
�xTNc����S歱���t���1/���A�1%���t�v��m�];:>�z��I|�N|4J|4"�"k�����:�Z6#_��g9k�R�b˾���ϰ��`�*��H֤������.�E���*�&�[@�N����G�>������̊�el��O��HJz�E?�uO�V�.�Qf�pi���Z�L!�wr�O �]�l.��	ڽ!f���� �eJ/x�|����۠"d�;�JU+C�������D]e��@M�`	��^�P�N���HIe��ߡ��\J�_Qr����\h�8&(���l�4UL�v~��,V)�I�F�mm�RU��T�&<�@�I��Rj�H#�]�̃v�S�D����R����{3���w#����)'|����Bl����(�@Fz���2 &�~.����J0�ű�jt�9ݎ1a���AV;�j���[�ī����V$��2ؠ��={B�������K��m���F�A��^�j���!�˄�8�-`VDO�Q��upd�h�g�T���v��W��$����i��E�t6w��������{�Z��_��= =��(J� �G�ߝu3��~G�d��b5{s#$/���/� r����`��{]j:�����.�.��n��a����5��@%]�4�@B�2��f���xҿq�n�fq��&kv9��n�%�^�p�
���G���!}^c+�m{��
�>�c��?&�Y��ր+X��TS!�῞xe+��>�u'��o��7r�ں0�Y0jn��Q����Z����*>+�����P�	�8daj	�N*�+�^m�1|M�q��ʫ#��䔔"e����xq_�UO�}�*��&��� ���� 6��H�+�L��fW��jS ����d�w2�����������z]��q�C\�RUC}r�#�Y�� \L�br:"!B�jae�r��Z_��}% ~4����A�	Vb	�m>lq�S�����4&�q����q��(�+c�{��V�[�y�z����9�L����o��?C��糸߼\z}��!�{O�Śd�ʦ(��KQJ�k�:�Ј(K�Җ����`ݏ��DM��qU|pK�|O�	~C��ւI�a���,��q7J�j���HJ�� ӈa�0%��j��E��t87�g7Zb�"��k�7��ᱨ��f�	Ct�XZU1Ĕ!m��������#����ɘ���� ��U��U�jF7�o�|��d0뵲a���%m�w��C#L飴��BR��Y�$�0�.ɀ���v���Ly $���R�_7��YP��e\�ʚh}sr���&��G�В�/v�����AS(�L���"]6�0G��K,4�v�����?n_�6 �"�����u����2΄�����@�/�/���H�=*4˴����NR`���&R}�s��3�2���2���8ps�#{���>k��(��9�#T��-ܖN��ſ�ds}�<��bM�K%�oܷ��TR�,���IJ���MfIk�A��6�l4�����Sܥ���smP+j[1���Bn(݃�0\����f���S@O�>�3JR�t:m����:�2���e*b���������E��6�ZU,7���z�i�Ʋ��}!��'a���,IU<��)�x1aҼ��'��������"�	a�>=�}����I�ln��a'Z�SƠ��6N1_j���&^� �<�S�|���+l�)o��D|ñ�Aq��(;���\5�H��e��ӻ|?�c;�g��g�B��/S̞ZL�%EX�~�_Pt,��a�&<N�dP��{fH4(l7�@��e���F�a@č��˺O{��<1���%��?�j�M"C����5�"�-P�ÈT�%Y��8��`�q�_�0�x���	��[s`��H�ՆB�M�s������;�-X�w��K�Ɏ�Y~\lY�gֿK}����SH�ZG~�9�o5���	���O��QB�Y��<3O#��L������U�)������siy5r�.:�v��m�̓��x�
?q�@�9��h����A:$�X��(8�h���s�̰���lN�b4�G�ޛ��Iۼ��҈�=Q���Q�O����{��2��*\w��s�J���pϠR+,\uH��RBu6���!���Z�h,�͋T  �U]����)L�b H �
�A�C6Q��k�	rtQr&8]F��-��Iz��wK��;�&?.l-Ś�C
�83$fJP����;P'k�����(<03�oJ���Ï�
~g����[���uwU�{GyS8�Lo�'����.��Ĕ�T����Z,��%�WVU��)b@7�{+C���P��~a�ZGXj��O�f=I5C�&�{}���"��fCU�+i|T���8����*��FZ��'�����!2�6�*_.��ʙ���V,AZ�1m޸��)t����0�JJ�V6�%�j
�{� z
68
�Q��04K U���L}b�D�������?��[,��:>�0�Iȳ0��|>Ս%)�8�gpZ���fS��v�3�� GKX�Mj�=#!�?�{Zx��R�3�!�O����K�ǒ��.��+߸��&�_]����ӻ?\��rY�	ŨjQ3��z��.YJ��U0��L:���KU��e�*rǁ��<K��Z�C����@\rR�xZ,ښ��1X�f�������3�@�/�{�<]/G��2q�v�b���oyk���.rm���?S��Ei�[���wjP.|�Ăչ"v/t��IL�o��DxanF��h�>� ;`з$%>A��u�Ϫ /��S	��P#ص��a���fo�Z�`]�E�8�0��~-F�wH��pl1�j�˗��ݽaC���f�Q�ם�������e��Y|I);�܇�¶o�H>P�9;OZ����@b��RÌb�Q3H��Gc>�5·}h$� ��;�C��;�¥z,���||���{�2|b�r��@3«e�b
���Q귚HN1O�{d�������*;�01��X�a|s����@E=�-xH_j�Q��7���◪�&�G�厞<���_�~ 7M{��kcɣ$���n�����|��Q(z\#����)�p������z]!�$�qsᴉ�����05��n�o�����N�Q��ob�:��M�}�+9ҵ�^��?Kͧ&�}G�:�6��T�ZW7�j?w�Z�kI\�W����ED!�M[�s��C�|��{n�Y!�J�О�Z2&���hJHB��L�,�ũ�	��x`�����;��Q��Oh�O�^Om �T�
��i���D�(5��R����@-�I�>�� �w��:������Z h��-�UP@BNx~Rz?�V"� x3����ENG�;�bv�����Ay����U0�r �ٚ�Vn_{\`��:�ZIZ0]����P�-�E��A�c�ve�ʟ:*�l8��O���zH��%Ē�ʮ�n��y�3B�F�AJ5B�ڷ�vK}���w)4���������H�ݩ�)�3*���ƮNʿ�J;@�+����L�����*,2���)������9�90�i��a~���R��~*7x&_N�݆�9!�|�K��iZ�V�/��wZ�D�/S�Q�ŧ�kF��R/�p�n�$���\���~b-Rx����u�������J�Ȧ�<3�K,o@N𵟗�L����b�����+Ι�$�a�r��s)�^�k���(����?�a/�����w-�1-X\rb#��.����gh��6*5#�n����^��i Ρ�*T���b�����T���<
���s{o$N�wDi2ۖS,�������{V�`h@�%ƀ:��Pчz,s[.|��ʀ���d�/X���Ji���)����^#��M*��
ڵ͊m����b��ɕ9���t��4���"*ȯ$̌��+[Tˍ�,X��!7��1����+Y��װ��'��<����\�\ɟ%����ss�]��KT��k���W���v"/p�Qv-N�
����`�e�N��u�,B���^��IL\�=b�\<kZi%��l*1�v_��4�(�3�b�6��e�y��؄ڴ�/�,���I�;r��W��(c�.ߌ#ƚR�۟��g�=Ə<��=?�4�psR�}f�I �z���_wi	��,i��#ݠ��� ��i쾚j4_[���G1�#���'4����꽉Ey}F�(�~ ց��\�������t�3�`��	x~�zAkU�B����7�o
���L�V��c� qu|��M�p?O��Qfv>�7���q���U$��S>���-}�p�`AE���t�l���m�b�{�*.� W*�l{"�[� ��c�d�:Q\�Z)i�;ok� �o��NR[@�w(bT:��y�)��?j�`��S2��d���債�/CHq��7<x�ğq7w�L���_
�a�ovv�Ǔڄ�Yǋ.3 �ޣ�u�3�7G��sGWcZ�#Q���7�13��4�u� #���, ܁"���������D�:����*���_^-�e��Xzz��X�D�'��nGp�z��:�˸TcLT��͵,.��WQ����v�)/B������s��"h���&�yPop�zg����/$�2�`�����Ib&�Y�M��B�)����t�Y���C��o��H�s5����8��d��+��.���d�8�DLA�9J����F�D.Un���e�����MH��/��NcAU&��'��y���;(c�Wz5��O(]D���th�� c��tCG�,Eosxt COM��><�ΰ���T�lM�x�e�S;۬��a����@=�	e��s�G�x\�/�K���[B�|��pC�]�»�v�[Ǹ�o���u��א�I�e}g�ƪb}1`���&�P>_]�՘2/�y��tv�Ov�IK��]1[cb3%�ԁ;��In'n��3§��M�&��7��녠t�����)���,-L	�#r|~hY�G+*�~[�Gbg�8�����OK�YF�c̡�+v��� ��+Vc�'��k��2�j��>*�$�@-<�SfIO/҅��d���~m�I0��1/l�?�<� �潳Bc�@|fDܭ%~5��y�RF�kL�-��mR��YŲ�ݘ�T�'�p�l�.?n�Q�R����ǋ1�C���fF&};�O���X}�x,خQ�&�I�D����Ƭ|�{2�kr���	)@�RB�+�d��B?z\���*�S��<.Nk^���F^J�x;m�'K���MUTn�`4,�@׎pQ䎡L�h"���	�г�������Es�J�H��Y�3���c�mS?�l�G��Q�`����JsNN������ގ�2`Գc�;$k�����Xr�ri�g�V#��ۧ_Q[����Y�������z���h�qG�l��~�K���OދN@�F����(w�Ţ�5�@=}W�f��q�`�N����;S�C��n1�'��:1�?\�s�Q�O-�1�v V8��"
�_[���NU�)�
�su�.ju0JA"�J��G���XL���H�{/�j�;$�1d�ϋ{��D����F�t��6���E��d�l����p�i�-�{x}�#w��_|ΚW'q���rpP��=܎�"{L):IT�<ݴ��>���yt"9�lR&��S�\C�M?.j6p����+���:Aُ���|C���e��Q������b���e������&��N�'�g�(�UmCO�n���Ϊ�[q�_�.�=n8�!�!Ht^`0zo�p��r�B�>#���������w�h�'��hEQ^�r�[��	'�h4�Ԧ �O��[</S�v�Qr��{�����g<S��<�U���a��-��VH�+Gf@�ǣ��U�a�E�̆�8YY�?��%AЩ��[}Tr�?*��_�nf�hvE/Q4��/��Go�V�
_���e#���e�'��d4��7���m���`�� ����$@s�e���Ʊ�VqÐ���~�C��f�-�ضW@�Z���oi�������)����;>ʸ%{�.�!�L��FY��Q�[�N����I�`�����ܭŉ�����Vl���x���>�HO��!�4$��ڻG\�y�����+��MAdF��!��z%��ysSb�V�jG^ǿ��)�1���nU�G��>jNZ���r���n3��=��J�)2��z@��lC�F�w�^�������Ls����_)�|�l��,`ct��3�����S��4j*��T�x���,���lg8�bmq��߻��^nf�90�TTX�Y�Z���s������ԬH1��9��+���>,F��Er1���IK~|�����(ry�Y����p��
��n�B����C����,����WC�Y��U���$��"gW�T&����qV�B<�i�$�y8��6S�d�+����t{�/4�M����/A�ҝL ��.S���F��d��b�>�fx��\wj�(r�԰�[ �åvݢ�B97q���TCB<pGi��b�t�Wj*R66��<�1P���}�[�=\��/��2�3m�_�"�6[�#��	 ���'�\����f�M�6̇�`o��T�s�]���΀�`�.K�ͬ���:�m�NKB�\�M>
"r���XЂ�5T�N=����6]�>(�	+�p�0ɳ=��/AЛ��*&R ����m
���hM��^�;HD�zZv�������ϴ��o�V�c�6�N95��I��D��x|�/> -&�Y٭K����6V��e̯�~<�����xT�m�_H����9�֘��E vI[h�kJ^�t���$��͉0#F�����;����ժk8��o��D�b��t9�~��W��X(��T����eI����bH4����lI�����@���tK�>����պ?K7�1�Kb]�٫x<����LU��(�A�>�(�4��� �f侗I�X� ����&Fo�����{mVJ�8�M����kM�3����ֵ��͢u�*>7Z�z4�]V�S���/U�FrQ�g���.�u�^�J�UyL<�z`��U�'��M����f����"��=j<G�V�J5h@�u�C��6-G��&��t{��{�^�|�ݬ�Q�c�O�s�;��q�!��Hf����&/_��౥��8���S���,+����(_m���i���"��F�^d�]�3��T��c��/�N'��KF�<�  �;��f�tl�^C��,ٷ"0�m�Q1A���A0�2�Z�<�F6_";�C�C��L9qR��,��e�[�_H��s�Ԥ�����+�$�p�s��}I�%B� /9{�������p>@��ɹ��P~��s�g���ۅB�#3#S�z�9i0�|y��#�ƶ�W]:N�|������P�*�4<��]!�Pd�-���RҺ�Lo����8b����XY��#r���gSx��(F����6��"Vew��Tde(uV�$�\\�߽<p�(�|��e'_���=��#7�R�h�7A�>��V8�n��0�Χ[�m��D�œ��;���׎�@�)��a[J����-fU�;����H	fn�Rx���&�k�̕�w�͏��GIl$|oƍJ�.Ta�pm�]���z~6z�QiU�&��8hO}�w6I����:i��M>zHU��/v���s|0R�}\�}��s����;���g��`�z������"8���ak&HX^�'lE�Wp*9����&�ˊ�%��X qzd�|��vno7�g�N/@M��Ӊ�
��Z�N�n*��&�j�\�������"gA߃O`�a�.Gp�
���0���w��A�����jo7��'wq���w~ho����&C��T�*"�QLf�j�9!4Ϡvl���̳P�}�XZ�Ubm{�����~KI�JԀ�^�'��\��IȄ���DJ�U�X]�k��4��J��lU��^bg�ͫ�ܙ�O� �c3�-��ޙ�e��aߣ��ǹ�P�+��w������	L� 3YU��5s�'۽��cR��^���k�-^ùm�-D����*h%n3�{�_X�n��j���*t�bf�Q�l����Dg.cvP��O�c+^	�E+�����*�\*�PT�����j���o_g�f@���?F�$­x�|(��.�ߡ#]�����0��
�m��8Ի�t�!�y��l���g��'��T�Y��B�b� d2�&��I���s�I����,�}�6�E^~��	/TL?#�W�!]d^�Ɨ���b������C̗����rv��M���0߻�2��\
A�,9���+PՍ�=؛,h�0�x��U�qj�v��45���vf��\ :�(���Q�TLd���K2dk����;�Y�6�߯$��U�4&w���r$�S4f���fH���" r��/M�����@�Fk��c������@��!�?�M�ib]?�G�Η
�ͺ0��C�����r��)o��|�N	qZO*�4�I})�\���+�?�mW�zC�Y<��f�����.�~���B���%�ɦ�az�5����_�Z�&�L;O�k�C��H�°�P�Vy�����扲��Y���߸�!�a�	�z�v�T�s���(C�f�L�fa<| �؃R�+a����u׆S���~�v�f-�ϓ�գ%+T���O�t� �қ2
���ѷ�������kB��d �.�O%x/��1�����%Z@e:�6i���*�� ��E�j^<O	a�{����J�:��F����q��vS�4;D�N�|N�F��h�B/��9���Є����h�� E,�JN�t3,���\�^a�o8���O���r1���S�WW|}��FLe<� A]�j=�������L5�]sg�E��ݲWlG>���}�X�{�B��#�䶉yxBOe���V��SF��b)����?�'=|f��@Q(�]d0���b���^��?���Ǧ��z�QzI����#��]��Y��I�(/���L��9�|v���"?{�8C��dB�5��N�m_���|�M�s�Dr�o��!1L\F�E�)�k��~�T"������绺����i>�}�#ƴ�8�f�g*��� �ՊE��/H:�L�Q���Vh�c�E�A�J0��CM��w���aH�����ِ��n��������<��w/P�=��+U !?�������6��K��]1@<UYF��g�+�|�h���@_Ups�Zh�-�g�O����������4�zV1.�2��������_͚�����ϯr�Yt��J��2gz0B����o,m09"2��K��ݬ��'�!Lo���\�fm�}S:zwd�f��]�#����P��y)��.����v�Y���[h��D��	�x�,�ȅ�����_eW�>*�F�D�=�j�^�W��Լ�u7.[�R�넻z���qx-����^���'�A���S[h��u�	�)\
���L�l�jc��Є�h��QW�?��n���J`��l� �=�,
�5\���#ţ��a_о�W6}��yaO�mڨ�;W�Zk�Go'br&-�ZY��?��C6d!+�8��j�D9|��8ZQ��(���?3�g�H�å���'�r�d�)��Mv�qd�,�J��ؙ!�Ó2�A���4�!�(�0��c��I�f�����Fh�����(�ƦkcP+]�@��*��r�x��������!ߡ.C04d &�{�����g-�'.4{vcsg��N�|%I$�J�s����Ԇ{.��mH+���o�>������Z@�2�Gk�h�[��s��1Kh҆��ť���*�Zl�n"KO1df��1A��{08�����Ak�u��Z� D))�Ԗ�mz�'���*�A�l�}��.���V��ii�r!�z:˾�.Ү�ȷ}S/�)M�j��@0����Y�E�y���]���4��˟w@˚�6�C��֯�o&�[�o�/���i�[ek���W�k2
@��H��=Q��b���|'��V�����o�<u��O(�e��*��&5Ʉ�,�2(1\3�C���:��A
�НrC�j��gã��:�w2����ٱ�V��r�l'�FT�fW�Q��@��w�#]Ul}�0�y�`����f;��]@�a<-w�^��;����5\v"���`��[�5	%�����3���)�J	.��~�h���[0�x�|J֋�l���_��Q�>�r�t��i��f��Q��ST��\�� b
�l��L[lI�}�é����P�R��v��t�O����X��f��.I}O���'�x})���� s�Uk����z���z�qv6bD�T��.�WT}�Jᓽ�*�c'X�zx]�T�]G���@�;N�=��)?l�P3���kTq\��c�跖J��f����'��Kk��.=]OD��.c���q3�X�3녯/\�3���¼��+�޻��l�R�d�"TV�5ԧ@�=�U���r%!�j����_�!���b���)�tnzʳJn	�=��?�R��vd�ܥ�����5�~�����>�u�R��!������5K��^)ȬV�fڠ9���H;ͣ#S\���"o٥L�_0[o%Ne5,��������{."���$�%���$c�g1����:*� �n]I���"�v� ����w��z�^eZ�-Д�S�#x����& ���'�1Lvg�q�U �*���Ӳ�ZE���+X���ř~�b]B��Ǻ�,���d�����bn��v�i�j�8?��{&>�ZO���[���3~Ы���$�����L���j.��	���3��۳N/�h\@!�m��g�A�ke�W k!�ʜ��Mg;�WO\�����f��0������Ю�AZ���(5��j�}�zS1c�����=@�<��qٗ�O�m��=���y=��$p��#�jD�NH��܉r��I	b&, �E��O��ϫ��~�����$gp%��>J��HY6�V��1a/�<��z�i0�@;����q���|�N���bl7Q�-c!�s�/�A';	���ڣ� �fJ�Rua����1��&.�� {H���O�LS`�Xɯ$�T� L<�Ҕ�̊����TR*����2�#��I�[������UH��ʹ[�/n�a��M)O?�Ha���!�e�,ſ�2q�d����x� ���ٓ2���g�܅�=��q�)����Y=����s�9�q�{����1�f��Jӯ�#]���$���Ƴr�4@���I�)�,��5������@m;����[�{3���4�62��o:�qϖ	��wlLP=ˣu�%�T��g�iꙜ�?K)4�ý�NMȜ.+Zɱ�~��3�<�S���X�=K��m��ꢙݼ�����D.����ⓕ�X�l��yrp��TW
�����݈�+w�MeVwX��DL�γ��=R�}&���Yr# �k��!��G���P�b�;g2M�u��Ud -��c���	�c�-�����[>�9ֵ����Z�@=����y5t|��r�§4.-ԉ��ɍXd�Yc��- �����Tњᶱ8����L${�/1KLR�u�:�@�|P��XU�X(P�{T����0	�)Ay%�Ch�[��G:e
�dn#��F�Kcsp��w?���#	�3L6^��dB�"H�ݠ8�}o�l?����)K�j4�t��A�"��#�7{��5xJ�ZD��wb {eK�l�R��9#yo����)���D�����b�65N�U���Ot�#�c&p�G�#*�+ʉ_�vQ�Vs��-r�*$����0.b�(��������mA(4;�R�)�?��|�3��ЛXL)6�&�ȶ�CpM� �X��﯁=�!��ù���[p�?b���4ٽ0�q5�SX/p����&�F��x���Yz+�f�B"�V7�='�(�X���dAqG�»�F��jL*�~Ʋ�?aWA��4$	)��XP��e��tb~��IK�#��e��!����*L�竹׹e���s�����I��}�0a+��qϣ8�b���,ݑU�ҖD	����@ۈD���.LEL"u��Z7n�]C��x�憊]�D�>��ltKi����|`�k"��>p�A=>�s�F��@�*6�ڑZ-���o
���	�� �N1��ʭQ����h�T�p���'	�+Y��f�~i�쮹�=�b�3�$=V�ۄ�yΧ�����$r���Gm#F	t��&� *H��/¯Ǧ�d�X7'����:_\���ī d��#�[�Y?F�j�5	���˳�����֊8�Y3�`)���m-�r&�"u5���QĈU�m���-��P�흃��#v휬�m�������� "���|�0� ���� rP�����s��9qz�Uk��������@b@��-}����d�"�g]�@�U�P
�g�U�LVU��i���h��2�b���� ����^r�}w�������cK�.����,�OE~L�@�n�q��IW�%ԍ�$���\v'�� ��B�D9gt*3wݚ�mqב�ʩ$-B��+�~�y5�9�=��!�2"`�)��u��*R	 ��;~
8U�ـ�����Rܬ�n���PE�U¸P)-/����D��߅�c �ٶ8�݁?��{�ĳg���濈H�5�2U�mn�tq �PV$f����y��=����ƽ���m3����ޭ�D�(_ʏ�����I{�T��K����;�G2P?����Xp=0$��ר����4� �{�m�#��4�V���X& ���:By�fU����xrЉų�hO�<K� X�:Ea>'s�w�b�P�z�5�{ͤ��(���o��>�MS`ɮp}�n���w4/�zr���\��-��a�2��3'��_��-�3��f��a-��f�X��{��>ѷ����$�0��u���55�hW�����hb����� ���e`�2������p#���x{�>s
�[�ӫ5%��4���1��s�p�v�U½h
�j��~��\���tM!�9*,+R��3�`��B�t:�z�%+�7̕㷰<��!b΍dJX/��TU�#��Vx�����Zw< <6�s�*���"��oi�𚱂�Ռ�.Ѷ
�uÿ�{�}�#(�R�w�#Q��IX�u�K߾��F���5��@,O��V0Q��A��o��~t��<5,խTrE�Wu��\��8�~�ݔ �sC8�į=�&���a/0��J���Vj������e�v��,���|�Y� \s�	�x"����?��lEФUﲥc5����T�oHC�����4UK�ɻ��1�jv��6�Eȫ�M	o�B�~�݆������q٘C.,i��^�  5�u�L� ���2��?⣂腸����2�JŽ�g!O�lӦ�hʸ��H�7��>�Wh^R#���>()��Cr�s.��.K(�Ϯ�
�?���������_��ڊP:��ONg����`���mɻ}i�gk��:�z�.�]w�v���i�N�wT�5T�
,��̅5�޷杻�lz�	>ע�A4U��p���_��G\���z`K�D�A�1�r��0&�Ԑ��̗O+(�-�?h�5�倯	�G�k:�%�M&Ҁ�s]2��GR�B'��4){<-n��Zt�ID�T%�`�7������sn��,}:�D=���3�IV<a����C�2���rBjԽkr�[1���Q��H�������U�A���j��^K(@������D
�@4⎢�B��lB�W�x�|����0%r��!�tj8�s��6[ܚ#*�ǵ�B1o��!fK��VO�gw|^��,S����ڪH�Qav�ݬ�9c\�Zz-<%f�yc��cH� e���<a� �!-�gNg��Oڔ����V��Y�~���i̓0���nگF�vy�e1���J����������z8=�;��{��*Z~W_�sz��'���g)��X��d2�'�Ne��� �����̃�ؐt��q/���!	��51�5� �z��*��1���os=>�c��ӌy9�Q��h��Um��t��E�۵�$�SD�=d��ֈ@��	CQ>�n�:��%����s�����1,F�t�rj-y�Lt� ���$p	�����a�c��Y�*�?l���4@	D8���"ֈox��h���Ǵ/��9���9 �n�M�������7|�];����~p�� S���u,"݈�<~�g�}ڤ_���nbG�>�@@/|�X:9{a�#��3i��
�[gi  �@�߶��u(L����̠L���&�n���N �U�^�x��M�b���G��C��-#�X�[�z��'�ww�:o�$ �N="3D�\���B�j�~l3�P�`<�J���g�	���F&[��
z�h����pg�H�x��3�i¬a*XR��_[MFEX<E�U�-qA{SD�e��U}03�S��8$�_�4Ρ��'�(w��*������~nH6/X�3��U����jӾ4�.q�e�ux�1w������`�:`�������M�=UQ��c3�o)(0�1=����W��|�j&�����lY�>�4��x(td����Ag�|�՛�9d%٣���WIࣵںd��!�s��em��B-*��4�<\u��$�s�d�WO����k����� d�:n�������JG��g
�ꢎ�� �먃��wp�"�N��NS �w�Vi7F;ʹ����Gq??ު`H�q�4��_�j�0�]�F�hg��K�iOWt�p��%6�S���[�6�XM9�1%_~����_� ��Ӷ�����U��&\��S�E╲~a��n]UZ!uðF�1Ď�����.��B	��������X�g��0����&(�y+{T���'cu��Y�Xkv�x�/8I�r�[)-<1���'3V8V��4��b���S����<5K?�zS��A�GR�cl��w�y��A>g'��q���Y�?�;�iHuY�a^���ϔ��=�U�**d�R8Jf6�[l&.�N��@ب�� <q���>%�śN՟&T_����Ƃ��b)\]cc�bi`U����XP�{�9�̺��H&�z3�).�A��Dbݓ�5io|��酮<{�#�[X�S���Y��z�w&��=ډ�[6%0�0֫���������vV-�-���|UE�o�D�#��3wZ��`޾���z���<��"O '�q	-�[�w�bG���!�ʱ��`�洍�"A#i�c�����F�k��l=!�@�[ꉨ�=,S�j����8����.N�!T*��#A����l��wۍ濵��$�F5�pQZ�e;Dz�N0HhL��y����*�Tm�YM���Sg�9�m!P��H����cKm5TX�e�s�KZ���Dg��8�5���sT��ЕPՕVݯ��r��t�C��V�[NJ����)�g� ���Kn�ğ$\.����D��z��:1|�#I�Yw�g��������Lg+�ğz�«�ߠ���- O��sa���	�U�E��_�����s\k�����؂ܖm�5�%˶���L6��S��*��24;L#�3�����K�<3��p���������]���S32W>(��������=����1�>�b��yZZ)�:��ݿ&}��^�N�~d�9��|�T�qn>7ֆg��A�	�P��O�F�G�ukqs��_�5��]��~��'�n�����cSo���W���hf=�_5��i1������u��q�]�3�#�o��X˴�s�+���	g��jه�P,�;��Z:�#vJ�^���4���Y�vB
 ����J:-�Q
O60DhX����C,;��ֆ��+�DOP�o��Ғ$Q�<Q��4�������3�R�I-�x���&�n杂���6����R�ݍ�АZ)	��������wa��	$�펿W�~�E�jFBǿ�5�H!��,�⥆�z�WK�h~mo\�#Jc�x��� F (��Ӱ�S���TX_"r�5��(�#�J�d����4�S�����aGC[�46��dZ�ӓ5�fИ{䗍�$�^�U�>~$`H�	<� *&�PIc�*��
�$���E�	5�9�q=B����R  ��ۑ��+v��;������%2���o�B�.����큝��M�����kf� ���5%�"�NS�po�η<vݸ?;�1�\�L�He1aV=���|1��m�;��7	���eg�r���mG����Rmwq�&zR��W/����+F�Pˢ��W�ō�6�G��P#�G9lH!�UA�9�x�1�O}����N�7��F�]���'�(u/=���]*��|��;k�4�D%��i�[�*=�>2:- ��m_��tc'��b�a�Q��s���;f�>��/��lXn$woM���S���QCj�a���D�R�'����ܺ�K,���,���;Ӧ0���Ь,�E������5H�Đ��9�@0h���iٍ��?�?���.v�U�q���W����͋��^�����V�l�}|�W<��� �;�`Ke�s����@�CAQ�p�V\(|�E;e�*oN��F�-q��j��Fo7weq�����+�b�9y�ZwR����؆1�f����p���Z�_v�#��-�����(C!k��V��*8��>"��L��*e	@��ΓրD�+'��ӿ!��iZ���Ğ��[�*<���-e�E��X�����18}d�R�y=|Ň������9
m�2|��u��!�b�`��[�'��Q6�Ƀ���4	���H��@*������Mca���r]ߺ��^Y�a��H�Q�1e��/s�-�h|���d��,g���H,��He��2K�l9j��X�T~����Ѕ)������7���ӟa�!-������ix��Z�@]��Ѧ�u�ǿ��w,�	�Q*J�c���E�9�`�'P]������AB��a�!��_Y�S�����O��Z 3�=|Х���]!�\�E�j3���V��`�j�p����ZԌ7IM���c��WC�}l�V8xg����;b�	����
���m+��Z`M=�k0�"�|��%�gN�U�Q��O���r��n�|r=���|0:1�+��拍��}U���J��Y��fH�;Yv��LL!*���]9�h�q2��%��s̈_%��hv4��p�@�eD��0^��Kf��+@Fev@ќ[j�� �c4��7uO�u/;��(����:��8:�\�m��p-!O󫯛"��Bĺ�1D�Z�7ŘA��Fo�p���)�u�m��ήvTosOu9�&����i�+F�jzuD��DIɹ3���!�O��!��Y��Vr� >���gC��E�o�ji�$��L7;��r*�gA�A�晧q��a�0��\q���[i\¸9C��\��P�ɰ���L;�����#�1�I�<9f^W�6�)��-�r22�q�!�Y��%�'�تDR��}=�bq8V鬞9й���/������%kt�V�OaDX�mZ��=�^<�(�7�����ׄC˞�?���<XX��k�7j@/Ii�7��:�}j��u7�Oj5�䑮J�8&T��~9#�%VL�xD-�����d#��0��]�h���7�)���N��|+�2t^���7U�n�JLަ�u�k���Qt�?!�}R�c�<�ۗ�r�z��4�t�~yVJ-�)L���r~��>�6�!{�lCR�ٛ�o*.�q����m{�S�;�|1�H�}81��j����Ur�gΔp�d��AtH����Y7*@Z��(0t���&a�\��-��L?�]�D�H�m)e�>��[ʇp�a���9��hm]�|W�H������$e.�Fm�	u��0W[Z�/B�g���8` Mlmj��Uo��: 5�e�$&@�x�?ʷF$��q8���;��0^=6g��D��6�����:����v�ݼ㈵F��{�aҞA�hϣ����]�$�- ��E����8�bn�p6W:���o�T�*�jr(��_E*� ���!�h��x�F�q��9X��τߛ?��B���;l�2lU2�|�sDiy'�jFE��5��ɰ=�uOԸ����ڐ�X�;2��S��`Ud�M>f�PR�$^b�;��������s���j�q$�"���xp,����Eɇ��`[�I&�):D�=b�M[S�ƘB`&Kbi��ΊI�󍚈��/x����NI��}c^㰌in�����+N���+�Ē]Չ�'����c�kI��~�n7OҔ t@,������鲥����b�������A_��J��(3��Ɇ��Y�U�1ٳ�5	%��7�3����p�ݬ?�vhoF91�҆ƒ����k�Ȭ�U����jۘ`��Ş�TeгU'���A�vo]���CcS�&��6�u���R�����%y�xKs�&�a#������5��
���@Ov�钞{��Ϟɑ`Ӊ��C{3նXp46i���|�Vdl����-�A�c�YQ{��-����-HiJa�t�$�%f[fhxBX���b�f0�����M�0������˗�����n��A�\ʿ��o��ƙ/uK��Kf��\:�n�
�ws�j�`��Z�$����ɺ���2�<ѕ��-7POu�E�4dF�s�N;9�WGԨ����$�!��A�m�E�o{�w��ԕ�'P�Y�,���>��/0�p�~�W!;��P��YPu��*p��V�py?c��0C�t�L��u���y���#�E�){	���\̉�Ɗ~�2v�8��F�ׯy\�l���ĳ"��ƨ,� h��S-x�C�"a6�1�Pjz1�r���:�pվ���i`	l&|����܋�h$�[��4�ѵ�(34X�E���S(��6��G]?��PЖ@�瓛�SgH��9��x��kDY�Z�+�x����xYPv	�)��.�dڿ����4~2���+͋��s`�~�'�.j�ӞUR� ���;w�)0W�#���ǖ�� t�J�߬A!��#�zQZ��ר?<|#�x͘إLe/��]�N�J����ud[��ࢋ�9iMZy��]h��-�͚��Pt����#Ī0=x�5�W�҉���`��Q�̦�\�/�����+º?£�W��	�|����lǽ��U�s��:Z��y��
}nD摾���GR�Оn�~v��R���19����u�D���V:S��b��׊Y�~�����?B�.������xb���a���z�s�P	�ٟf5����ـ�Gs��E2�����8���މ��|������ Q��D��ܹ��}Sq���m�pG�+��B�����M厭r1�E��P�m���K��)���`_�Rg׼�ҡ��I@Ȍ���*����Ϲ���`n�ڐ���wY/�*Ts��9��u�o
-Ѷr�������&<��)Wm�U!ݱ�(����ݕ����^M0M�A�&��b'Fw���~H���"8��A�V�x>�J��O�*ј����x�a>�ٟ��/	�}���(�~&|�@��,Kq�a����?��ƈ )6���=���j{�.=�Lp��n[r?�I,gpCڄ�l���t@Na�mf���vKg���Z�(�m��?;i`�Y9��»H�
{���VG�~��.P��+�>=�"W*�V�Z�=:�z1���Z_iQ��/�-��=���1�j̘1�袼H~�i�v �%� P�h��P���QX�&�[tVNy�{���a@�%�h�m8�����m���h�w�y䉬��j�G���}O�6[0� �Bs¿b�lE]��fNK���"#X^'^��d7�l����؎��҂��ŷ����?X���C� p���Z�q�'_�
��D	46��7������B���8�4Lk^�?#�� g�zC�E����º%���rd��٫;w�&l��r�V�9ǧ� +A;����%�R���:�a�-���	��	f����Sa�^�1�\�q�[`���<\�ڬC�Tlb��5��a��*q�Y���%OM�sDg/�	�V�ioO�c���5PK<�����L�n �'?��6{",�!?�̥�/K��K�g#��bG�vg?�n��\�� vf���c�V2d�q]��zcIX�����b}�o�"��p$j�N�HI��Ͳ4�uH����݋��4u��͇fnL�D���P�J3�[]A�|�@�,�41��pI�G��Y���}�}"2�h��ɮ����~����#=l
�s���`�|9�v�	/�U�:ģ�-�������{���´z�� '�q��0?3"�=6f�EV[���p�`�u���k�����m,;rm ��qgq�4(lT2����n Bp��j�$��j\��Iv����R�@wH��5����H�1�r�������ǏX�яo�x9r��Z���
߼6ؚ��:����at/@p��=�h
�5s��Ry�[��+v$��L+�\ni����9�=��M���	h�[4&�
���|&�=�iNwH��H�$db�ٸ�>�i��i��2�Af��W�v|�{@�����R�A�H���)]$�U�O��Z���8�����I�8�^��?�#��H�m��fоm[������n2��(�qKt��`>ș��(!�NO�/��5��C6���5��q2Sˮ��=����KYZ.�<&e#��Ef��77S��&��-���,��v�����
`XR� 4
��JPߏ����ҁE+w��_b�w�϶�X.�'�!,��7�;"�����]�.'VA������)(�o��(?/ab"����,�IzZ1bfg� �w�� �T�r2H�޻_�|�>-���Y������U��#�Ǳ�����_���	�� �@g�2,S֤֦��?��G>o��1x!�}��Bz˪
�\��@;#,AJSg�W��z/M�ޓt=���P��3؞�Y�����\>Id�q�Xo��F4�E��>�e�b���"�л���E������cr&v�x	i�Il��RP�$��!�Z���^����~}F��8�0����K4�� H�K<s0��*�s`��-�q���W[2ˈ.�����7�Ş5X������2Rkr����P����K8m.9�I�>"j:�ɬX�9*+|dH%�0��&ad�;"�B� ����D� �!v���x���0l��̚7މ^���+@ȯ��[­�l.��;9f��Qj��r�e�S��^ �9_Om��P��0m�*}
��9A}��s;H��z�d<��Ӓ?J���U�I3Z�r��K���B p�}o������ۙtΣ��'(<6s'���n�#{���M3�ؓ8fּ�伥��� !������4��E��(�R��z�h|���J�)�h�[J�h�짼�V��H�/�<��#��i���+o�K�]v9�#�з?o(w�n�`$uy��!6UW�;Ĕs�f���o�&�ܮ�a�u3
o4�����|(m�%%�tfaB��m�LW$���;>�A�*k�SVso�:A�0���	T�����I���
���15檗CR����@ ��2�P����YzÞ2{��║��53l�i�|B��ܯÅK� ���g�����5<I�o�nK�/�,�h
M(�e�47uw�^�@�)|�����A��C��|�v��+\��M��9���`�;8�5ڢ�_���9��%�Ȼ� ��A���<Ռ�r؋�������C@0K{�n�,0;�ւB��nm�G0fH���e��j{f��1UЧ|�={�v���&L�V�ѯ$%�kJđ ��"�\:Bn�[�b5�(x�[-6�ࢀ�sζv7&�o6��@׌�I�P��p̉g�#�-���w >�j�@��6�La�'N�q���ͫ�abO!T
�Y?�KHU�>��HN�-~L�P5����{g!t�y��'�:n/N�`�Xy��`��l(d��e�[�^� �"�'86Wnk�_.Ƒ��1x� ��]�`F�uȡ��77�R��&�H ���
M׈��	B��D�\&��+��"-Z��N��	�^�
��D��x�ew��y^���i^�%,X/`'y�����@0��]v%W�d�]�<�Ip��e��A��*L�1�ۺ;E��	~j-�ދ8�$& JU5s[i^a�4`*�N�#]Q2��oQ}�d�g�����E��ɐ�Äywds7OY�s��v��b��b6��\�`��z����;�RεM5?p+�{}c?�������^����959�odb�g�˩��ӘG���i"�����+�[��E��@�ρ���N��9�Ʀ�R�d��kwK F*i3\h#T?]��jJ�S��?��VH�j��+YHU����2H�_���� ��[�1
�;���?z���w=Q�H�A~��t��:C��i�L��f@��M�/�ob�p�Sr��r,��V�g�z�b3	]��W��,�窷<TK;t�/�����WL[��[��{T�9k�<� �KM����<a�H�,����x������|��DD�l��BXqS�Ƹ)�g�[;QZ��1(M�i��9E�eǣ��զlvUI 8d�
+d��.�2���p���:T	^!O |!�j)N���e��[��6r[���;x�>h��UM%�YM���)<�n���'����X�B�j'�/�+�?�M��U�N���/:ˤ�9�xH�}��h+8^~����<6����^��%���W��nVW�%�6{>�Fa�<R6��N�M�T��nr����GV2��.U3ON?����'w-�#�R�Nl��A�����ԩ�.��|O����
w��'!�~���|���4�.�#�1����R+��9��i�ݮb�2HZ&N�l�0A��re����C-�F;���D��)���>�)/?�pBYƪ�Q�5�"��s��L7��ȣG�\�U9�kp_$�t'ZH���a>���$�>�T�6`�ԯ'X��<�'8ե��e8B�3e�4�m_�d7��5 N�m��d6��'�ǔ"]m��kDI�?��Bt�(��4��ﺷ�x_`��u<�ä�]׬��>���N$�n��g�j���M�V�|_ex�RWW ܅g��'���s~C���jÉn˯VL8R���D[�3�U)'�B2S3�$�����S/T� ��|0q�A��ǰ�ľF���Yr�@����)��!~#׹�\��蠌?󰢫�^���s&R�mm�B�H��SŻs'��>x��̆��,TH�rM�����@�L[h4B�x:��6P�"�[Fh�� �C�˭�ra��������u>��I���W�B`����,���R��]���o�H�[D)vo��(�':]�Fi��抄hR~�s�2W��Z�	PY,�@��Na22f��ⴔ�Kox5�A�	���ȮZ�xc�{$��xY��Z�Jn��Gb����-GFEpEm�n�ǔ��y���qA&�T�Q5̈��Ơe��1��t���~��{�L���5�6.�;�Dhug�/���N+�m1�ǘ�^@�<%;�����ē��i���8�ڱ%��x?��c�O������N��IH9�	0ݟ���R�?�uX�n���Zc����Rw�|��s��<��
tiƛ�:�L�|���{�'�w&"NG�	�Em��(�?�M%�$��l@�]� f"���Ϩ�v.W 0$b������ާ?nr����^ C�|�$T5��YVޗ4���w�#��
��WH�=�j
��j&��t��� `�N�O�^��w�5��Ý>�vRh��� Rrw�^,�#ᷯNI�a�
A�&!I��r�H ����p�.���p,�^�[[�i��!OR�[��c�G�g@}�!�]��;���P]��7�!�)��}0|�7���o�X����߁��W*�DU!xX��vv'(�w�~L�JQ�+�E��f=эe}<��z�֮����e�3�!��n��N��-��P����t#����rfY��)�!�
^���U$|ARot�������AA�"�f����$��(µG.���$H �����И�L��hj�nXi0ԷV��]��V��ɍ��5+8��xW�tX���yޅ撡��	��e����Ut�6L�h����?����d����8���t^I"j��Ү|��ŮZ��N3C�?[��5u���>;���߅i�I��ن6��C0��G�IH�^�-�j��M�?�V������a0cT��W�&K�Fv%�e��9w���l�]��,�%��3����X8�
���r�+b$� f5�@j��_]1tZ��8�4,x��F�0zZ��a���DMl)�8Y��M6E��RF����d�M��MG���_'����;���'�Mn���ƌڍj����������wzL�d4�Ô�^.���=K�W�wRJ�u齚��X��������׼ݣ'q�A�e��Օ�4��
�	��ܵ��*��zސ��'��r��>��#SZ�V(��c�HS悼��Ǖ}�s� ?�u��GZvj��cY�X�O	� l+���0[��X��z��Oq�'t��v
9�I{���2�}�|��vT����F�)�����<@NO��z��A'J`k$�=&x�4 �d)rJ�����}.P����L� �r���2���A%���0� �����bju�%gF�P �m�z�i&�G2��C�_�7��yt�� �q*���8C]X��`A�9�����]�	ړt��T�Hh��2ko����R2)M}�5,����X�J�-�c>���{}�mױ^R{��xK�Ǭ��cu`	�\N��aɣ�.CT� �K��3xԧ��K�-��Ԕ�4�[~��>�
6��u����F�esO� 
���E	�S}-�w\�+. ovis��y�U%zs�Ȉ�*�jhTn�;�
��L�u���T��ݡo�H��9��GE8��?>���<$s֫����Z�q`���pv��V���t3�@9�A3pTg�ŉ�S�SH�s�
B.��7HI=�M��~�|�~_@z�kݿ��b��Qg�=zߞN��ml��C�떰��q0�����5'ͫ�*ť���ZU��R����+vksJ�G�7�߈�xO4��k�%�&�e�r;6{�ųg�w�I�������T�Pol�ƹ��/�-&�@}0�ӹި �;��If�v3G�Lխ�R<?�FN�(٬	b��+K�=d;��>��Ri�v�jU�@.s!�s�ʸ%Y�{
a�F��8Q�����`fR�6��9gŪ�Q��;�9����E�ٴ{;p�"�;z��~đ�l��Q!pO\~���c��%�8�
��QWEP',r��x�_��Pcʮ[gVN�=H�^xd߰��b_�0�&8���ll�� ��3�SsP�RE�a�7��d�m/5�㴞l1_wsS�� ���%����q"�|T�UG>J3��P!���8w9�P~ �R��nO�ca���8��wQP���t�˭ɫ��!�/����B�YW}�2mS��U#�|�C;�xH (�5)%�c[�4�<��-E�(�Ж���5�^H��}����0��~�q�fW��I*�!��v��tíT�Qt"�<��*bʰvw8��8 ��P�@AzPiEq�/ӛ݂W9�����B��aK�U���ǂ��������;�ڼ|�-��؏` o���)���>l�߲���~�^�6�ޫi�u��k�ҽ��z9BA  w��k7��-P����Rxe���Ƅ�E��t|;w�y���yuxc��N��4UC ����;\_褓����|�m�Z�ߖ�Gs	[0�2���
�� &$�
��eN��#�����l�j^~�	E�t��ɔRw�fi#�b+֑ɇ�Ś��zQ���Lꓮ� pԟ���+&X�&͉��i`���U^o�~44�ӛZNq#{$���;X��Oh>uKt��X��W>��+��$p�m�u�Kŏ�4��2Lʛj�W��fgϋ�X�&��k�j_��^���\�Y�h
F�0�XMR���H��ћ
"��ё�?캯��^9���?5��;R������'���gi���_#a1ˠ&8
�LL��g��D{�و����|�:{;+�n�G�(�=�obx����O�M=G�!%1Ԅ��c�I]���@Z�As�
������*���]i2J]�2�T�#|s��t���c0��o�O��}߹���f�~�"���r�Do� �}`Z�%���'>��e�v�
��F;))p;ȝ-v��u��#Q�8�f�����L�@�J��+�n7�Mm�b�s,� �[Tȃ�����<\��R��Y7?���h�4�
-��J �^�[%�?��
��R�p�ث4ZW�Ǣ��8X��\QO���?��_�̢�j��L�f�#Gϯ�(��dK[�#��51���f��R�\�ÿ`��
�C������2"s�Tz~����¬+���;���
��y��K�H�F�/
�dA��������Ҽ�+`{f��J��c�@	����!��i{W�xt��ԅ�U�;�^	y?�O�6�d�A{���m�%��׆���Ɵ����a��o�^��쫆fr��k��Rr�|~u�����h��H@dS.� ?����ꁪU��j4�T~}���q���K�1j�iI�ڢ�<�E�r	q*�� ��3o�CF���lt.�$� p�����!���z �H��)#�����A�J:>.�5��V�@u�n�߫ͳ^�n���hEg���ʝ�N�P{��ʭV�IR=���N�g��$����W/�=�Ĵ,�x;�僮C�XF,g�k��vH�1�9�e�xy4-�Ͼ�������s6�9T�[���4�cC��<]h�U|����{s��D�[O�/.�tWTJ:l1����ٝ�3�ټ=�z��^��:_vܫp���h@4..u;M��]���<z�X�L�����ʐ�(�\t(6�z^k��F~��-� �P�僖�d/k�t/�w�O���1�8��~��z��|y�Te��?��5�7��~��}�0�x�u,t!(s���>:7��\�I����6������"�~7e�%�����&(�e}�3�A�6�<�����	���+��v��(݉��/%��Ux��M	I��.ĩsʸ�wn.�I*O�C�߻�Oyª������h��r���9�s��aHy9��I5@P������w���Fփ���Y���$�A��R_�a%�q\u�����7s���P�cӍz�:���4m��~�ċr�{�af@|`\j�1�fq��d�/���P�"]M�AG~g�j�a`1���/>I��s��M�����h*'=���O����V*̅��QVA�	�-�Μ�����4~{��)��G�����x�O��2�J��1&���R2�gƆ)n��I$a�!n�Q�6�o��@^a��èA��lS)�Q]��'�Zwbh@��}�B�@�]Y:'��e����ܠ���H`�`�mD<����RXw(�-�!�}*&�����H�t@�W�	�����	���S��B&v�e(Έ^絩6'@b<I`��i�Q�"LP��V��/�՚ǒ{�|�U`�fd�Wů�*bCS�;�o2;^��ig�m�];�N�A�2(4�1�z�W�R4�ͩ~�����tH��������8+�X�<_�)x�ݙ�;�y?�K�Y�wA�Ӵ�P������X�u2\�@��I)b���\3�53�Õ�L�UÞ�V�!/�߰��`xS1����Z���m����c!�4��������9����n��F�NtLrY]v�L�
X��	���0c�U#��m�	(�`fL����_��f+A2��J>�sw�C|7^^���~:�k7y�AV��o��]�b�Q��F�n&\��2Qh�{��YVt�� �lH��������Vdz�1�&!if�S��51�L�-�+�(�@���ܘbf����7[�˥$Ɯ��GA���b"�a��4;�0y�Ag���Ij��9����,	ȗ�����-�kѵ��tŤϨ��?Qvc�Qđ�Tz������&����{X���
�� ����l�ݲb�M[�3
�{��l�f��Yx���sj
a�x�K�'2��s��ȔFf:eWL��'Z!�����`���(Q7��T|b��)�Z�N�VL�A��RHPE@��`:G
�I�s���VP�J�d��g�=
�O�����~<"]3��Z�E�/�f��o��|֞ds�I�ݕo2)�:4�sN2B2��\O������3�O���"�)�Ԯ	��'�7�X�f��b^��7��RSÿ�`#E�䁓m�xѥ�7F�/P��?�()O(�gv�Z���a�S�czv��>��E��}��.�Ep�`E4������t�;�����K��5U�^o$�6ɆޗϟS��ݏ�DI��|+HjѬ?L���{�fA��������v��eY�ª*���@(�fH��@E��W9?j{8
E��j>�6���*oњF����qJ������{��_�J'�]'%���wF켕̱1+���}%���]#RFCb�����wL0;��Lƴ�1H���em�k��_}+!K������Yi�Z��!�H~6���ȥ��s��J�pmxr���|-cD$:�
��Z�q�"�_%�iUG8P �*��)] �G�㏴P1�V'E�k&�`c�a�on����}E�ύ�p��
�kf(k� =E�h�JS|YB'����G�5�P��=�:8$�ZK�$��5��ڧ���^$)�S�����K�"gϣ�S��$���v>��ܲR�
�ֲ(Iބxu�X�
8�w]��
�N��<�ڒ�/܇Q�6�G����>T�@���WZB�e��2y��H�{��d̔�m�x���ΐ��nl�N�:`dܝ�P��gN�c��Tď��!/qq�>����@A���@S9�qi�Npj�nn�H�k�*�v�Ǯ-��FSB�fm���+�
g��1�W崉ɷ��%�y��1���͠E�ϣ5z!G�D�־:��?ќ��}�O�[eڈn���5Oif��;ӗrF����%�.�2�y��/T�c���O�d!|k|8��v�[\��YN��n?wqDd��̶wfsx0�(��1�q�
������0Qcv���d�����,2ޏ�F�Τ�c��Cj(о8O�Fi�1:�6>�
�:���w���R�=b3��#�Q�b�}��ʚ��p
E��X����&�)%��g���VϠ/�2��d�I�̣{T�V�,�7����@*ǋԒ��9�E���('���W�g����1Ճ�+
K��I�x<��kT�I������;^��|�c��pda�qN\�!V���1�
5�4�/���`�ɽ������������rg7�q�/�ma�#�[52%��5+�N�i=�4��..nT[� h���g�t�p4ޔ�Q����R/�+���U`{�R���M�T(���¿��R��
�E���
ԣ��,=�r�"&rXh�	0�$fD�&\su|4�w@Ǘ���K��`��1�zL���jB5(���88S�,���Ғ�q/"@�d�&�ч�R/'����MQP����,2��&^���#P���/05z��X���5��Rğ[OAa�0P������\�+$-ܧ݌�����yA� "�
�Ѯ�_�����R�n�;<��#5�6BSX{�ĬU���	dXs���j�zGdC��������Eҍ��,VpCT�\�d�����ePC@N؁i�I��yO|��5����;� �s�o%>�Z0�o���z���&�7��������d��HP��{�2Ӡ�/H㗒,S�*)3������ݽ� k�<�ah7G���0c@�?�{�0�d�r�g�_5X�G����;R�'&�Q�_�L8`�aU9.�k��cN�@�O�@�g� �̍��㔀+��D�������S�,~
d�,��♠�*tfO���f^H�
�ŏ �vZ���v}��w�W�������4�bD�9�:I�ǐ�B�C	����s�&BjK���zK��jU:\�5a_>&�8t-իl���/V$�$�`js��۲��Wx�a3��WJS��`0u� ���+����
Z�*���E�Rz+����9��G��-t%n��!��3��,��J���]��7�&����P]5;Ns-B,%s:IMF(��HU�ҸWAK��|�����b<�0)'=gg��,�԰�0�)d`���o�4^f$�h�<��\����ٕ;$K�J˧�*/sVu��o�4�LÎ�n�&��W���.����ͥCǴ�X��9;{�_����S���w�ظ��X}�}y�5<ԁ�!�x9�xM�csh�&�YoX��:�w.#`���ǃL�	�����j;���oB셥�����3=[�ѭ�,��R�є�U�乣��-+4n��UL��@�n�J����Z����楷:����{h����3�/f���T���c+�<k�:U�P��1��
u�K�h]��F+�ͪ�騒W'�G�3�U��]�G�+q��<H��'�i���u�c2�4����)������tT�`�iU��mf�N��(���_�{ND4Ŀ~5�kH|��^�0�4$��ă.��4�����R[�W��$߹]J��6�U��uk��Ok�����-U�f��ΕR��E㘭.c��22gqܩ"��$Nq�٫��A�.-�#,��o�5hA~:e�N �݅�%��F������U0���z�2�!,Q��I��b�Q&ST��X]��vA\����F�� �<z&ȫ=*-�8���&ڌO>��m���o���9j޼p��Ď�ICl�ǭ�9�/F��D;@��t����鸧�����������d���>���=��6����ii���Ǿ`� ��w�[{���h�b���(�oP��.݆��~|�_+I����:����RÚ"D<K!v��x�c��WL�BX;>��/R�������HHFBզC�yy��qH^��B�NQC*��W(�~ꅚ�vsak$� �R��rӏ�M�H��{�.R�(]�M8�ܢ>ő������m�J�]cC�VK
��^�H	�* ���1���:�zL���O8�ڣ�[H�6��cj�Ȼ��q�!�K�G���N�*2ן��܅
d�Ɵ�u��
�x�q�;D�MD;�Q�n#�w�j���\��В5B|�E�Y�㝝�i K ��H�b�Y�|i4lP+-9�R�	��ᴿ��V�w�u�������=|/ι�a�zkby�_�ήl�ucL���!�mƯ0�jK����b��m	.S�\?U�>Q掗E��]*����p�!��0��1=��_���x���7"#��8/�g�����Pv���\�Ex��.�P���v��>�k��y��W2�u�sP{�A�z[�^TIt9��&ؑѺ,X�ÃN�;M4ct��uL��q-'iN�o��R�"5U���3�"�l�"��r~�H� +JYJ}�~.ܹ��_��a�`�MV��,�����W6�.��8�o�yH~nb�<o����U�U���m��iF��|`<�������f��Uȸ��8c��{\j
rй]v�+��^��]O�����p^�a�h�Ӿ�좉�A牎�`�5a���)��n60��D��K��X�����A]x���ɭ����E��D�R���!l���)*V��r�Ґ�Q�q����6��Ũ���O���JJo@�����.������2���B L��t�j^�g����H��JZzh��U.'��]�JdJ��.vFj	����wҩ>��<I/҆H�.`ڸ� _�����la�e���<�'��H�Wƀ���ׇ�cs�>3<�]U8g�kl;A��~0����>���W
�b���$�(�u I�'V�qo' �=��:��:	u��-!�<��z.���9Ȳ��kV��l��>��ڨ81L;u����^��)�]o(lW�m8�_�BC��:e����q3���;+F%;Vb���&WUـ@�N���#�N�َ�Vgӂ�)��4"J���`���ް�o�x�@k[���VZ[;�B3��͋�T�����`#�Wg��|uGGV����5}ѧ�hJ�g�J.z��`��
{%;)vY���^���"����N'_��D���X��Hc�Oy�I&E|�G��17���T�w\�,.[�q$Lgx���G� vQGxce�&Xl�_��4��a'l����h�4�M���Zo�
�Os��c:���\����8�Vz˭���&��
l�ND�Cd,��<;V��6B6Q���,t��4�v�8[�ً`Kdp�^���9[��_�u�`��n�qs	B�.U�Aqi�$�
c������y�a��8�_���Q������1ߖ!S����k"q/�������1�W��8�O�k�կ��lrC�����p���I���߅[�\9���k3�|������3%~��
��|��~%'�ͻ���F[���`K��- ��e�͜�g@��2�p���<C_��D$|c�K�L(A�lk����5�<�`�.Wև�\Ch�Y�e�֔�x�z&�p�����+j3ږ��l`0��[r��pG�f�����n(� 8N�o�r�aHqQ]3�佨��6P�a,JB�f\��%@Wh܍��>�he:���c;�g��0cxU�l1�3s�������F1�G�C�\����C�8����S�%#�z{��x0�W������X��zcz7�j_y��Ϯ�n�pT��Ƚ��\�ɍGn��.@�WvH��fI�M|��ʔ�S)�[�H�!�{>����'UKy71��n����xs���ҫb��T����h�F�3�����h�^�L�|R��� LX����ޖ�t���I��0=�IOs�X��5T�ո+���t� �\��6��у~R/��d���%Y���
C�U m�t�A�k���#����.�f��_�'� e�4��D��i���!���&щ�֫`�R��d��=�Qv��[/��.�rˣ�%*� l����bI�9���L=���m���U�VsP}�q����X�P�p��F:e����e�in�|\����3}�_��*��1wl(�磖weO��d��=��tKlع���F��
SٱY���?�!J��{�2(e�N�,/����mR�95�^�z|/vg��eڶ+3�E�o�9yZ�M5ON~�و��s�t&�]����Ķ�ص#�� ���T���<�.3*�D������ޞ<P���&(����Z?��ݹ]A�&6�tE�r"�`.�q��5 xE� ��Q�����m� �3$J1�]�CuVgt=��^�7���g%(	�P�*	���=:G%�,�n�q�6��ѱ-j�7��_��P�N����Z����QҐ�Q=�Y%ʂ�8rx�%^g�V����OB��`}S�]i�i�?#� '��|����_�7MsG��ϓ�b�xD۷e
5���j��xɐ��Rn��1Hb�ñ�E�BU�Ax����0���h��k��Z�G`��N�}��7E}���sH]�MRXi��OFl�$��$T��Z
���sq��jr{)T�"�QJ��i9F�i7���5 ��sL!v���S���f{�$��$�`mJii��ً���!���r�V�����>�:���ʛ
g;v+��}@=/����L׌��Ji��Df�|^�=>���y�nz��v�-�9����/�H]U�D���U�
���������O)V��y��W��T�D���Ԍ�0£�$��)�V��@tj}j��q.P�Բ_���l��A�	4���H#l˿
��ֵ
�"�<f��*�{b���Q+��g��
2"b�T;�*֞�#%@�+���,�(�6��I������ �ίm�k
y@o���|���u����7ZA�`j��G�^��n�	4���\���WY\O�5�*f����'f�9�c���е\�D�iesC�b}>��e�yGD��M-uf=`�)�~P�`WB��͸���[6$��E���EV*�[؈F7�	r�mf�֣CI��Q̎W��V�9��H�ETO�ݤ��Q#''�D����;}����i��ڬ�T`�`�xÆ*���}��aD���n�C�_j`�lo��۵SVhh[܂(�t���h8/HJ(ICCb5�� �w{l���sev��mm�?��tA�؟
+:~J�!�P?�y�O�ʻ�8�B�� ��.�>c�v�`��?�|���h���>T����������?�aW���ȸ�n�#àO��~�_�scWs��H����s�;�G�Ʀf��E�#D�AET;��JcY���'B�ӆ"$0h���mx#n�g���"�`���:�zC����	���Z�c���%fn	���4�!U��aO'�Ԥ�ԤG�ewo��*��L��ER���w�̪h��JC��"|Y�"����F)��P`���rf��X�1XT�	�t�Ÿ��;z���6p:��1��	*�l
2t�Aw��:R+� ��2�/7%O3;_��(Q�� E�'ˬHE7��e-e,f���+�������ƫ�틤�����,j�yiK'I�RO}>˰V	v����&�Z3L���0�m�j�n	��(����>gvD��T��4��*۳ދ�ѩ�}�\�n{�e:4<YC��QV�5�>�����N�)~ȡ�J7g:��/ص'���Ņ�dYd5_����(���w:�&K�,�A�$�ʩ0(Fj���L��fܳHN�'3k	���#� *w�+
_�H؟7"�X��DN��#�
u��
^!�gG�H���r*	�Im����9m�\d����/DD��kT�]�������cc�2&E�cD9D�9q�� %�J����J8���m1'J�@��m��d�-A�妙�t���yQk;@M�e����$�v�)�͸P���4���y7
Ki��b6���l��e����|?��#�Z�>��-a��&oX��0��w1-���Fl�i��6`ݡ�����[��&��	������n��/�n���s��=g�S� ^ݮz����5rtXy�:��	ܪ�v�E�"��[0Q���^�2]����2,�Tl��RB��GO�_�I���I�rfS�VM0��Wq�A�Z!�OX���t4�����������7A\���*��m��I������QϠ�x����"Y]�VV$�rƨgZ�*�o�!��n��ນuEV���	]?��msM�U�o2�]a��	��e��m�}����1}?��v�VԐ�Xd`	���Dg+��x�/�`�e�V�>�r�b���O|}���d�]��]U�?B2��w��z�B�arl�����z$vy��|G�6���� v�ؚ��͛�.f9��ŉ�X�& &&��I����q�]@S*7L��~8�#aJC�cJ�A:f�w{�3_�^Ȓw����-y�B���F)������ö�+�r��{'��VF�������'�s�	�\�	�
�t)wNڕ	�7v'�;�ͫ��3��X��ݑd}D2�!�x�
8#�f��#��A�r�ǚ�l�Ds +}�J�n7�*�ؘ�*�4-Q�G��R�8����co�A�o�{%�[c�B��Ȁ��T����
�ڱl�l��@ ��\!o�';��|�v�x�� l �-����ݸ��Jދ��OQX(j{�qmɷ�b���ۮH��7/�3M$�<@�1n�R����o�$��B
��s�%��6�¦.#a�@�I�W���㩲�Qs��$��~��*	-�\N+c��s%l�V)�P?�@�>/�xk��1���!��v���R���&�r��v�Ș䟬�?k�4���Z���l����t���ʵC8�n��9�a�ͩύD��HT�=�'Q*���'+���p4�`�nn�J�J�>�8�+K.n����Q-g_ߨX6��J>���	�=2���
1��lV���nƊ�u���T�v7I^��S�9��7���4�ٻ���LܖJR���:���_�w9$^-o��y.L��@�9�HZ���ŧƙ���"}�������6WY�$]5���0N�/	^o�A5]������~�����V���#dꑷ`FUr�c��V��Tm��C��!�?����/�Uֱ��Ix�KkjJ���N ��e�m=��ĕT�7�;S�r��V�=����/D��������D܋�����8�)�a#��6q���,P[�#퉢r��Z9w��7�|A��{�	� �66%u���ڴ�DŊ,.z�u�Z�}э0�<��TOހ���!d��Оpu���{3$��ͱ)�4}�d녁L0��$�4ئ\�հ���K���8�SL���TL��4�('"�1�S��q��FZ9Yq�͡�-�����a/*$03��#u���^#V���W�O���<պT�����P4�+<%��Ta�H~��N�~��H�c��B���Xt0�h�jjCY �a5VI��8^�:q.��Ϡ1E;��;v�k0��&�B�v�bNF:�$f�������9��ֽ	Ě:{���N���$X ��� 5JknmZ��H�2"Ʌw�8������`��/z2JWL~��=��� ���T~O�ǀo+ۅ�f��/}�L�=���V�,�*��3�,�ܳE���8�E�*!��Δ���Y��)�@J��<�u�'_��A��N�shpχ�3��F9���j�-6(����R���L" �)��#��j� 9]	8q��j��3���tج�8�Z���a��Ť&#n4t׎�}�y�~���
��`�{̹��ә�[�;�$��z���|:+�]��%�p�ޟ��D=�(8_�H%�E�	H��2h��#��F3����Z~e���	D�G��*����1���^�P��F�;4����QP~`]_���s�!��`�1wB+�SP���q�&>"�Z!�����"�k�l��G�&,��^Bg��sQ�Ť���$
0��u	i��w�� ��h��!�*�z����|C��Z�~�>\^T�y[��:C)��۫ԻP����B�7F+�r�B]�]��!��H�}�	�u�u�l?6����2L*��U�淳�>�b6��4@��w[m�3a�VQ�������(���!iKB�l8�%'kǞqg��G���Ǥ�f�u1�s�?P�[�ok3�(1��� L kz���P>�|��$����v	�FH�v��AyM	Q�-�Ot4�#�Tj��}��LN��X�y��;E���4�~x�?wJ8�$��	��C�7D\L����ME��D�v�٤����MD�-oBI����:D�Pb~T{<:*=�ު�*�j��0�>���UW^�T�S7lPvF4���Q�L��%Ѩ0JAu�̎�#PN���VPA*=Nxv�����|��Ƨ�{[�%��+Gd�5�~�Y�k�n�D���#������0�)�w�	Œ+$�cn�\z����.���%�U�=�Q,�%#���<q����_�g�ќH]n���%ȩ���U?`��LMr���k����Z��̾����t��O.��,�oY���I���� SJ�- �J�t�0!lO��?�d�J���q�yp�ew�@=qӌ��rj`CAw^��@�g����{��5�x	���js���0�;�<�$p�cT�8��5&�P{=JǊ���ދf�..F��I�wN5�l2|�Gc�Z!��?HQ�$?��AּՇ|���k�0�����߽���'��������Z�u���B��t�+�r�	�CY�*#�׽y@�<�U:F��Nk�#g���44;�j��K����S>�7+��L��u6BN�ߖ����\�찦`����z�d$�x��0y�E� ص�x��i�s��D��������o�����`��l�T,1Y�$}K���� �3����
Ng���k0�m��֍�~�J���0�Ikw��)�Z�_�:+���_�� 5�o��::�mcH�e���͹o��w��ʗ���NLm=��}����o��-d��BJ����ck�į���D�'EUGP�D������͍�wkc�l���D�p#
�!߮m�(U7NBM,/�E��rj��.����Ѳ��X_(��*��z�ts��9��"1l9W�ydhZc��2A&�2�[�܅�w��G����S��������lt"�~Uv" �-Xi=9�� 6U7Okޑ\�G�Esɬ���L-�kӌ�;�_�ʷ�9ne�|�l=�Yf_7��@���Z)���X��W��о �C�Hd�}�4I�7c&@H`L(?^��1B�BBևd��3���ql�����b9N��<̶yf�U!�TB��K�x+3Q�����}��r~�EE��`oO8$�SL]H���H�����~T�j��$�vI#�gn�n|����-��{�sI$r�#+N��F���:���)���#)�ιJ��XQ²�-Im\|)s1v8���� �VS��Q��l���#ɳ��
k��ѰW��\��w׭�1B��[Y~!���۪�uФaz_��gQ�]�(�Ƽ�y����6�X0f/D��_��R" ��I�聝X�!�s����#�ሑKRgu��ޜ|ׄ�@�4�g�HE������<|���86�>r�;2~W��V�-�B���hӦ�n��wU����R��y�-�p�3Z:���!��]s����m�@��g�i�U�d�u͈�Z��i9�󵛘�7���$�'������6G�%���I����\�����T�z�����5�]��Ab�sdu�d��I��sa.iQӐ1M��������{�9[��מ,��W�*��^�)o�ғ�O�� ��-G�H�����a �I�=�I��������I�=�Ξmz��x����i!�E���3����By�'�(�ݸ7O��B,ֻB�]ҢN@�{>��˔��2�����<�/�%BǸ�ۯ���ʎ��e&��1���Xў �k㚐@R���;����m"{`fn��^�z��F�e;;>��k����Z���hR��LA�sM_���=�T����|�9���N� N�4&�����_�vb^�����J���X��	��n���t#^�yfh�k�	�B�Y�J�g^�����7h�CŴ�_:+�)$��]��F=.�L^h��""G,�6�Ip7�����n�ӱ	V�X������t�o	�v(�1���
m�t�]C�P|4��V��I�D8�[�Ѝq`k<G����(9^]"���!���^H�>���Mvu|+��m�J�B�	!�|���@���+�U-.<��X�U���>��b+Ol�9\��yJ��S��Q8�T����_��q�(Tݘxb�;��Ӌ��:�x Q#]*n1�m9����Q/�����T� �(��KO��S����݇C�SҔg���>=���PV�M�/Dȯ�k^@>p��R���͠*��.�4 ǩ�x������[s��xS����-��(�;h������[�s�a�?l�� ������*��ChKy�	�I`쵧�~P�үQPo��޾��k�Q�����G~δS(U�=��ARI_�<�Ê�I�}"%G00�΍����Z�ܻY�LKO%��V2Y%�e8L#3:>����^#���ӥ�݇wu�i�þ���|c�|��B3�:_Ue�D��!�x�i�(��8YG7o��v�,	E��r@��}z?��߯fE��mn"�A�p#��+N��l��ǭٍ߯ǒ�ĚAT,��]��4�d˶'d�$�x��o㉸�t�|�?�tCZl+^̑����%�N]Mu�6�4���"Pޖ ��I�8�7�yY�jzIm�l�ͪ5�Qej%A�]��w� �/�Ŵ��͛�G �+�?�j�����G�ES��+Ԓ��'3���F��}M���7`�5��H�:�>�g�ur(#|{�X�5	d��]F���H�
�� HE�����O���g���"�-Q�E�Ğ��L�{;|W�tc:t�Y�@�Y��@��E8?e$ ]Uݨ�hex`��Y3���A�����\�<�R�E�	a��e�
��C<���6��v�d�/�;<�J���qi�:Dx�u��p%�����7ս�K2Hs�|Kh$F5�L���A��ďVkYܳ����J�9[��Vv)wf`J���|�I�� �ٝ��qCM��Ip�H�p�(=���D�gQ$C�2�sc��j%�M�̰��!w0n'�x@[��z��B&�����
��e@����u��m�%�Bǉ�D��<fݣ���Q��>��v�&�B�Ej_�-�P�_W2�;�B�%0�8q�u&����6��$y�bpݵ1�h<4�����wQ�[�>ˬ[�2�WU���A�-�������B���+�hO�#TqU�2O�!�y=�\�4���I���K��
��]1lN
��~����+��&ӭ�~�:���*z�E'�4�u��>Eό���Ē�S^rwB��%n	珠�|s������.p���V���1<��w�Ҏ�	iW���!l�<�Q��9M�4���A
�"��d'���N�P`�ս�TD�*�N��.	>�NE��@E9O�\���u ���ƞt���6~�C4�me7T�)=Sy��΢e�jj�M��(I��W�}�+Hސ�$Ot��n#7�~kWJ.E��H���B��o
���]�V{=}-�w_>Aru/:|G�	^�V��� П��!R�%�l%������H��E^t�GM<D���^_d��_g�_or1g�K������XgyE�������3��-�g�AE���Z�Ӿ��İF��Wp��.4�C:ϻ���;��������?Nje.��~�c��-���'ySC�r�h�/�q����jc6��n��[�-q?/�4
�m���@�a�y"����;�A3�2��zg�Y����L�k#L|��u��c�{h��>n2f���=� ����F������Yn�X�;p�����"��m�;�;�:m��������������o!���D����[�&��f��=[C�#�m��r
v5Cr�ӂ��d�rFfpK�ǜ�N������`�>%(K7�����6S�����{ _=^sTY���Yo5C��h�)��Ӟ��s���T	�$���;*%O\�$9������������g��|�S�		�׌[&�f�� cc}f��.���νel�nD��"��s�N��.Ĵ�v�Ex���JFk�(�K�%B18��1bB��4�#��zCU.��+��cQ��T���g�>)ϱI�������[دI+ �M]��j"�z�E��}K��i'=ڑyAcR�'<��(�Ԏ�]�}�x�$��V�p�_�A@�Xxa��:h�)��e��{!G�S�4Ql(���>�w��#����H�^��S?d�ف���T8k���9sẐY��� �ZY��.(�I���"�]�%�,���k}�'�0���ɴ2z]��L����q����
�1*�3kXY�<��@�@Wȗ-�����I�E��|I,��a��"E�̀z��;����R ��}҈`�a�p|u�*�y���
Dfb���[E��mu���l�q1D����v��dNF�T1Z���$b��Ei'Bd4˲�Қ���q�x��9皛S�Ys���9��}�`�{�S���3S@�� ��}���6M�?�c�NqSObjEP����(�
*��Pm�J�� aC;T8�i��C�Rqg͒�<�qv�0��,pY��4�y�^Ox�����ܪD	 2��J"��O=�����:�-��95�_�zi2��KB�k�_���e[�a���\��3k�o�݌ E�P�<EUm�.y��.�����h�M���~�2`%n]������I��`�p7db�������	fNp�J3���3�#5->W�Z�]�����}���jÚ�\[�A�lu�i���-��v���U����T�*R��^�V�0.��P(l�p�pg'!{��uF�Ժ��Q�,rMM������?�d��k[H�n:�����VZ<!�jc�Bg2*b7#�枓�zI�Uv��_'5&����+eĖ�!m��hM���{dL4�5�$�\��-#��JhN%`�Lp:8�|��ݡ��h�H'�����/���y$a�|��ss���5Ft�&���
�^aw�Tt&u��+u�������d��/�ڎ"K��Qf���#!t�
�4�i_{�_�%�9�P4{Ń�=?u@M�(��z�;'��K���&zvHR��M*&�N�A�{ϡ2��T�ULю��������L��Q�q`+��^oٚ��2���D5�Hc*��F��tzW�{]�L�̥�?�ڳ�j�������2�Sd�lh��"L��]������-w�Ċ>$i�/���>y�����R���H�qt<.�/ɨ�5ӗ��h����ewԕ8rI�s`�X�ᓌ�"Ї�	�ZLBO>:�(���w���'"pi����ɉ�S�$�W�3�����	 /��+}P����� �6J�~I�/�#��ò�@�"o�A�4��m�����"m#zn;*�E�hw�Gb�]��
�1���N���)���Q.8����%��}j�@��L�o`i�}aݼ=�p�U�w��8�#�+��gmE�.�T��� G��D�����ƣ�.�>I{����@���cgRor�ҷ�GKx\}O5�?�pL�w"�Sߏd��>}�T��<��酲R���\���M��z�Z�=�dKOX��W�q���H&��c��㙴��p�@�	;�'�1���ے[H�u�Tw�-k��S�%H)D`���!���Cmp&@w+� �&�Mj�t���Y�L�z���0���64e�Ri���ƞ��Y�汧�PA�rwx�={�R��V�n"p��k�-^W"w���ڧ�@��5Hҏ�`XYs
��JH��Z"�L���o���=�=^�+�P��^eTM}�̰jK�����9�V�a��n�9�&�v��?��z���?�o�����8@��^�=fe��P�|c���Y�m�a���wRU��W� ��<�}Ð��鲳>���٭�9	����|i9>9Ы
FLe6��c"�T=��c|c {8^3�0!�P���
�F9�9t-z��m��:-H��Y��s���%]$��?a(&��@�<;m�	�D0�AQ�2�͗��/��Ȫ�q���`��ok5��j^��z��ǡ�� ��'�+$�N^}�4�C�ȶ��o8��/~w	������󮂜���m�$;H���h#0TՃ��7i7Kh��T^�����������0�L4?�H�|�芑y)���H"X��#���j���A�pro0+H�x�h�BM�K9!�V�7W�)$�s��D��u�$���>Nt%��1��'OWVb�3'�w�G^� �Y��"�����|`��3�Q�nQΦ�$o�GU��^1���TO?F�+�QFF+��ޒ�'�Qlv�-%8�cd�pf�����X�]){��7�~��k'w�*B��K�v8;�|�/�����[ɂ��d���y�fZ/�Ɍ�߮iQ�0v�fJñZ����愭jǅ��Ȉ��#��:�9[�V!U;=��N��
>��jn��W���~��TP�~!iU ��B-Ļ�FQ�����z�Wȗ��	V_"�e{�O�҉
��v(^�H�|��b0$��<ň6lC��o��`ۧw�D�L���u�U$�3�*>_`�4���@�
��U�>D���vv\��:���F���1���-�W����VŎg��g0���Ӈ:��D+
4(3�}�̃b�%i���O�q0�Q0`��<[ly�	-=\-���0q9��M��m,T�u��t~�r��)#���8�'�3� B�h����]�ߨ���,���0_F��}[1���<�א� ����p���\�����?�b}�K��On���A3��s�N$�n�׃�s����Ox wʻMl��g7�?SM͝���6�+�{�3��dR��5l 0Bcj���]YQ]^W�,}4���1lQ K)z8U.�0{÷��ة�����lehD��w�B
�7��j�{�?8*h HW�Sv����|��%�p���DHg��J`4����\ҿ�
�������}ͿS�fp�N8{��;�v�(��>t��:U|a)f�0�E��!���Wz1���2u#���qf}5�")n�qR�Z�g�nC�у����ujLk*
�T|����C���[���)ჅQ�GY\f+m�9���!�rd����z���)���#'V���f���(��$��׍�Al��=L��>��Go�II0���s����*�j�A�+���%��iw/%��Af
^�xi��~���0C��k��&���$A��Pʻ^���)��%�e���|!��^����"9l�w� ��9�]W3�!�u��1��a���	�����]=��ߕ����	�;�(�2V����,7�����tT(�lB:�[�3�$V�ֽ�/�5�7�f0��i�˛0��81�q�5��A�Ҹ���3���?6�ظCRsT���,�{�6/�u|�t�}�����o,LIbF5Ҕ�7�7���x�)�j/^!|9'@�9���e�Y���$,���7�PfpF~)��66q��䅆gv�e-�G'��i�ޚ6Tw���=�����9a��^
�4L�Ы?^91����
Wz7�O�L�)��^	+�d�H�|�7�Ҁ�D����]r��0�Q�������"+@��?�JWV���*c�#颊�y>t'�x�X}13�h��%�3?#��ɉ��b$KV|Kb��Mz�oT�`x�N�������yL[Z��o�����nA٤(��4l���%z?��oO��p�!b[gΛ?#IH����JXӍ��6����0+�������;+��%4(��jŦ�᎑� �3��|���5��yy�!Ԋ��w2��<CGK{�*�������z��Q�0y���4;���q�����\��p��Ǜ㺟b������/)�V1�7թ�? /K�����
I_�w�;��9.g~�[B�(Qk����z=���,����?|����=Ăqm�(�c]K\]�1-E�c֍�r��1��Љ�:M��XH���r :��[?�v��t�l�
�w��B�����י���f�$�\-a%�d%��3��>�y Ǽ�/����C��v'�X�	����BR�c��ʨ�L���A=�v�0�<v��f����ǔ;�ů嘯�j�=n��i ��6ō�Nz^]PaLe����@�:�B�<��ǖI�+*���y-r�"ߦ���F��r6�=A� ~�f�h��4M�QL���w�X�p�p\T@"�RF��k�k'����梾HO���)�Gv�7b�S
�y ��Np����G�
;f]��E�w�*k��RR<���k���{vY�E≣#u"�q�I��(�E�ە�}��*;S����B�)��)$�>����&�$.i�9�f�}~�e廵l����,�*h�/2�<�B��ށ��!�DV7i��SV�G�X�d���2�@{@����Z���|�[��F���zG��M@��p� �v��i��j��U%������;f�����?��s�ו�NN_���8h���~�x^�=�j7�_h'�H��(�%�	�ɑ#�k�һ/fS�,&��sBW�B~V��U#o��K����G��4��9m�,��������L?�(�S٘+'�{v5�)��k8+1w:K�:4Eṇ�o�,�lƹ��a���A���%�����/$�i�6�o��P>�J)�^��D��4�к怒��¦���<��|ښ�"3�(3J�J����1 ɾ�����@�tWQZ�����T�~�E�G�\���_���jHX�����^n�{�p���6�֡W�l 2��)kn �s�C�j�Y>�E�N�qo�5f����O����=�pE��
�.^�!����59���V�T_F�B�G��-��w������?r�h�׬�4���룴����&�R(�{\,r�#r�8E�iQ��T���[\T�Z�oY��D�` ŗ/�̻yU$�����2O�_ï���n�@�a��:(R7��/m��x��G������~G�C}��%��T�P��G������'���@`̼���HD>�K3�vt�_��!o���L4����F�c9^��J�Y�ߋ?��>O���wa�l�~�q縴�$#�=��":$��D����.�p��Py�J��Sq�"��.�a#au�1q���y6�ʢ�[�-ؙ�A�@��O,�a��	�=&����eШ'>MM���{��2�D�>��P�8����W����W�w���W ����S��T���.��;�|�d��Q��Ͽ>y1�]�d(8�+=����k�+]}��Ўd-`�.h"D�8��ҷ��J�K��p��d<�aK����>����\j.������X�n~'���y���`ÑU~}���y��Of���i�+��g��_}ԥ$kO�6 [�mHUv+�q,0��3ѵ���@�Wf���k�m-��V4�^���}�j��� IIH��\~͢�aL,�?(�T��=g���Jq�� ��n�e{�9���4x������fGr^]��O+�Q�ȞJ�[c�ࣕg�m[��0$sB#���\��&����	���n9� �zOH# E�\Yc�c��$�����:S���	%H��u�Y��ߤŞ���a ��G
	)�XO� ���[��jR������͵Q�r�h����:3����7�>>F8����o˭����\/��F��x�ecƢ7�>��v�_D	?�I���J9<��u�"E�t�l���~/�T���,�^��r�Lp���t��䂚ǎ����(~pJ�d�q+�̎��xiI�L"���_�T1e�럇��QJy�x����Q�HS��kҾуv;��;��t��W8���bL3�g�"�� �C�V�{sg�1�l�k.]�9�����U��x�(����6�%;���Of���H-B��frq��}�������� ���X�"�wt�~���*y�~ e����!��]��@~i�L�
p8���2���#[P(���ڠ���W΋�'06	t�FÒ���s��he|V9JrS�QH�ߎ��ȹb�qu��ۢhO��s�_�$��>�1��D�\a=$c争�#����H��r`�n&���C�+K�;����7m�IP�*����|�x�����(t��s��ǜ���C����6��s�Vs�xTN�d9H�pw�_Ƞ!�&H��ۊa�9��qW�)�rT�Տ�B�w��HF�p�-Ւĉ%�4z���� Y$p�T3�kV�{���c��܃���Sg��	���'�_v������ܓ�%�2wpmt*�5O������ȍ<7�؄���A�%/�ǹ�'�j�
�F�� Ym6u[f���t}����P��^D�S�ne�Kz���R�?8����;woH�>��16����-�@f��7a��Yד�綞VѦ��V���D�:W�aXc����,�����g�� �%�<μ�O�]9��=�<7+��*p��� �e�K�&y<�4-�݆�/�\L��J@$=F���!�h����^��"����>�|��$�1�1ki�����z�_�\�'e2N�Yj����F�l�UX���I���n�)3���J������:�x4�57���*VZ8��?��w�X��t:r��M�Y֥��	{��j���UW����k���o�W�D�D�H��T1��:¢rl�9l�>� Oj��.��8� �) �T�8J�cؕGZX�Ox���;a#����CP�ji=��>���R��׻��.��f��1��5%�������$�2���XV��������~+����]+�N�/���6]1���jc9(t�QS�5ݍ��v%�����L{�nw{�x��-R(A������]�&���[E-p���D`�q��cfM^c�ҷ$GV'R1��	lkȡ�4�+��Z�j�.�q��V`��]H�I|0ɔE��i�ڇU��Uk�^��}]��G5��0�ڧ�(�b��IDCh��=���D�A�c�+�	��$F�n��u���E����g<ǉ��� �rN���Ŏ
�B|��EׂǄk�+_�Ļ�ٷ
��y���pp��.Ӵ�_�r��}b�)�j�%?��7Y�����T+,�y/�_�R���e+�>��w���aO��N��;N������� Oл'U��>�g����$,��s�ZYx3�!��Z�<�ք�\�Z��u#�*CƑ�-��ɒ�������9�?;�D{󦁒,z�q�2����ɴ�%0��U��� ,t��\,࣫ͱ��!���M7瘂�	w��L�a�����W.sN���a#�$��J������������i]������'��D� ¯�q�``�Ar�Qi�;CO�൮�����M7�6b�7 �'���v��C����PA�n�������p���at���(t�`gr�x+�D�#�n�Ul�S?5�H!�>��k&2�s�����=x��O�o���CC�v��D���/^|�l� ���=ǫ�D$􁔸U����j=W����]�C,5s�Co,~?p�J��:?�|�٘!��Nw���ώXۑ�/��|�҃�U��MНB��jt���,�Ǜ�#�a�M=�{ϰ��,9��a�)�Q����3a����"������}�e;�t�Ԣ?9!)f2��)�mek�YyGU�����lf�2a؜�e��!�T��%;����ķq�9�rr�M�kV<s���N]���A�?��YHc��Y�xw�k�-��ꠔ�������ѳ��*��}^�����t,�kڎ$���z1aN�I��]��`KI�O����{��V\�c2��}�ʐ��5��7��G�]�J����K&#��B'�T���#)�:�m0IKt�Zw=�j�niי맫CZ>��x۬��5.���-4�H.s����K�l־�iߵ-	�9���8Aѝ7�w�'p.r4�����vM�m��]��{�gۊ�e��d��F,p�U�ҥ?P����ك|���AN���! �q�>`���`�HO�R�*uC)�4�瀂oӯ����U�v����]m��$�_`�2=m���r�Ŝ!iI�Ao}h�(A��!��� ��18�Z1�6(�oa`ꀛ3�k	z��XFLx�dEC�q0ڠ!�3P���Id��k�u���m`���cJ3m�u�'�hl��q#��S�h�˕�����2vB��'���b�������y�ښ��IO�BA6 �;�IU�N�F��7�Ņ(ޕ�D��SQ/?�?+�=��a���Ζ�駸Z���e��mA��/Fq�<�Cbu�tb-��F��%���;<�@]jgIdHٖ-��3�����s|h�p��Z{�y�?���뎖X7�):�4�_4�}:q�֥:����`����f�$;)�{�g��D��+��`o��Vt9��!����^	�l�8���tބގ[t�>%�ɪQ��K�-s���i�N-���d֛���ъ���Ŕ�p&�+!+j�4�k}���<�F]�V�*r��EL�Ʒ
D�V��l���M����w��1&��P='cZ ��r{�D���*)�[��g ��-�G�Tp�׮��S�@��Qc��%3��%��C���e:d��ϚmL�#��W�}�ʫ�˳F�,��u�G����T1�����@���,4����
Q��FE��/��h%��(×�BB!�
B���u��Գ�NO�#� q}�.��A_ďI����wP8�t��"4@Mˬ�gi�9�r�����݋-Ls��~cA -k�k�tV��Nt��
|����cl�����!���Þ!���އ�hx��8�zC\u�T��l�G�K(�հ���K}�,�]aB�p5����ڿ��¡�	�'���A��z=O�
���gE�4�q�x���;٭�gUc�X7�m������m*�ñ]�kn��R��5�+/�h����4G�������p���,lW���������@�{y��:�"N��5T��at�Q~��������F��kL����y	�7g�����YUǽt%۳���$��s�J	��>��@+Qow�L��8��y{�K��
�;�x�#sU�?*Kl��$�9ъB�pQ�W&
�p�_2kz嫝y��Pn}5�J@ZUƛ���!A`Q�><!�����E!�S=?U��΅��m���$QW)�c!2K��2�.+���`��H�+��R�(��� ����,�?��2L&��!�&մ�/���g�$Q��%��PcW/f�8X��u�d���C%��-���-84��ݜSl��+=Q�����D��;-@�+�{�a,9���� �ރh�/������&���������T[Κ9���\h�Ì��/���7����2k�V�r�l��&�hJ� .^��rʐ[/(�&�Nݓ�k������b+	�gB��,��{Lӫ���n+��ͭ�r"�ʬ&՛S�%e����+hҰ�t̀�∭z���}��9D�o�U�~i�8�}���&�7Ti��V쯼�Z�{r�M�9n��O����y߄^ݝ�JH���Zؕ�KE RT����d�Ҭ��a�9MU?��[��+$)Bƣ0��MQ�I��-u�]���+=�7f=3����I.p�Q�A�A9=L�6i��S�=R�"��$:� ���Ԑ�X	��b"`.�"Ze$��k1 )b�}�5WtZ��t;���<pVoR�|�U����V��m�E�\9#�}�m�K�K�}����%�
U��,�R*aL��Of0)L ��&�䡙��C
���S��[N>��'�1b���k�X�		=��ew��NF8�� ���%�c�1��;����M��O#�6��j�s�u�nKp*��j���SJ�4[�����Vo6cc�x��}Sy-É��i@���Mm��"�ȸ/e8#��'Ț�t$Y��ޝ՟j]=����ȴ|���7�|JH���C�][yt ��/���(5b*�̱�q��
?�����[�|����#��(��X���d���c��S}����D0'�L�e����������ci�Z���;��X�̏��B��]z��[�ȁ��������)��ˣ�2���5}E_V���X�2o�l����,� ��eeTqQ;�ї����t�85##^��}�~O��-˻vF�Vs `9~L��yh��1�Q��[.n�~�~Ք�W|X���
��XA:�ʓgCP��K�p�)�s�ű��JK���#�Tj�)�� (�Z�5t�	g�Y5Dz����r"� ���r4v��wdg7Xr�r���8Y�ܫ�+��ݥm��c�;�x�P�d�`' �U���� ����w�C��Vƛ�)�;H�
�R�ئ�(r����g\�ז u_O�� ��1���Ƶh�����v� /z�fo�0�-V���C𼙨.�`~���è��X�P����V�g#U��hd��@ ^��Q޺���J�r��lg[K2�#@w�o���.·�S߆W�' H��$l��_/��
�4=�V���N����
�:	�^8��I��:@i_��N��Uu��efd�X�+�񀽛��$bN���P%�{#C��O��YѴd3{v�Qpt�|�����*��1�ڢ�,.�2�':>K�ƹ}�E�m���|j&	�wErތ��3��-�7wM}֍E�cSH��J��:��w�Z��9�?��
����%"i��s��AkG�P�d<n�����Xw=L�����@A�å��j2���4��vR�jTj�g�^xȊp{vGKPv�V�b^��>̼YxkcZ�~@N~_�qT��*hP�W
�lC�{C;�
��?Ν�m3�K��.sz*?&\M�s����'�q}���݃ѝ�%D
!W�,������a;�'!��|�e���_�i,J�,ϐ�笂6�,G�@�4:k���[�l��"�J�ɱK�9������	�R)�,�#Yų�<��<�u.+�	��h�L���H���}	�+��Irϒ�z��Y񵑪�����e @�o�LH����Gy���N�Want�c&���������hv�.�࿞-�
��N�a�g�%	�޷@x�X�N�&��� �"��&iu��OZ�3����6�V^`2B�zy^c�IV�pN�,屶����7��~��Q���qO��&�@���E�Җ��z����kg����	�:�C��3�'6l�4������̭�� &F�7IrG�vJ�3*�]�\�NF\�_�Oyek�"Iq3��ɘ�Rc�Ӵ�_����
�:�j7J��V�9�����7{'���K.��=��[����Z��e���F(FI��Q��%�x�F���mH��$�@R�Z1�� Lw���u���
�e�F�;��������]�j*u���{�C���<޽Gn���2�3P�7���H�-f��������ĩj1~͐_�pȂ
C�M�ú*���Hb�Fg�a����/���A�佯Je���{%`L�臠3k�"3""����32q_�2t��p���a+2;b��ws$�H����Ƨ%��>N����`Y������ѫL���
L�I��\��X����L#E�'�5�R f$mQ�B�8�8(�@������)�iuD5�#Hj���Z1B���>�-�y���7�¢^KV�e��N���D� !��:Բ���G�kGVEF+c}{����iM�y���{p�K�d�%09�|�w���|�"OO�	�}c��V�;���\	���ֶ/1)-ć|�z&���]y>_N�BF�.�Pjo˞�Z���)n�`P8Ū�8�͖Ҡ!�R��i^h�܀��w\��R*荏��0	�"u��"�U�ϡ�l��{�e2QFkѨ��,����FF,)��[q�R"���zx�����'���U�����W���ԃsWԃ��9 H,��n�i��M�H�~N�fa��YȽ�~�w{�+2��~a����D��F������eJpY���	U˛��hb{	C06�;���w=~�l,�G���8� � u5�,D�L̲��1�k���)��lF�N�����/&(��"g3}	hū���z2��F��p��,0��H�JwF�#)R��N��̻�g`�����(@�7Y{�z�Ӎ�&������� ř5گA���<��A�\�x�Gr6���O�t��Y�z�)[3B�׻�z��i;�}hK��u�5�V
��N�����3{a�m$}����L?ʶ��j45��	4xz��{�iu�-�=�`��pIO��� �~m�q"����dB��v�?��E4H�w��~`����q����������iEAQ��2� ��E��ܜ�N�(���D������X[� ��{�^qmT��G���k��A��"T9��;���b��r1oɵ�Xm�����y��}�߁�P�P�k��d�}�j�b�U�4�,S�?<�ڃu�Y�m�3Ȅ�X���_�Zxw;j�e�(��yIM5yϾƫ�b]b�q�5丢�ڝK]F]�\\��}�,���;gH�r���]h� ���\*t�o�Cb�g~c#^�F}��^S�T���a,�vm�xtX����@���a]�}��Uu«��N�t�j�h�_al~H՞h�L��/������0�W���E$rw���z`�X,)"����=��M ��L8�N���)g��rZ.p�"͹�l�dB���ο�ӈ$n�-bv#���s�ujBX@K�<z�q��
vg��q�����:2ܖ�N��}%�y��m,5�%�����U�G7���P��H�w$�8!$W���~��N-7W��xcە��2Б���+�W'I-4��� |��ڹ��σ�����wAʩ�!�F��Tt�;���4��J	9�c�F<���S�h�//;X��4�bB�O���4g�[	�t���I����!}	��nE#VhLd�����+X/B�q獷�*>�Y����3�&��1�ɳ�O���%W�
��7d��d�h�D*��Lؽ�EN���0�v�F�Mz��A�	�0���Z�����F�TJ'0��}X/F�Ņ �R|M��q5uAI��'�U�eg�'��R�n��1|��tnl�\�����ֱ��T�`tt�ȁ"W���L�ӄ��94n�Hv�I��p�G���zEj���6�wˁ�[��~��c�-�a�I���M� ��]{�N�c���i��X���̺F�*�1@�;�-�)X������Ժ���w�>\�ؒ�Q��蘟���������q���)����3o���y�sb�2q��`���8Zy����p{Q%�qR^ַ�fo�j�U�a�܍����Z�w�	�6�N��8�e������d���g�P�"���?_����x.�~�4����3��*����%tw�k|Zr@�E�H���k)�G�|Kx��^�����m�^Za����~��^�\���"�*�vT �	B�D���=�ݭ�ϙ1�?�C��ª��f#䝁��L��m����Ĥ��t�h��o�CaQ��6�߮[��0Ȟ�FѢ���M=���],߹ �Ψ��A !����;����d�kfк"<�
�:s�Ĕ 4�^n���Q�{g�7p�
m/��P}�{�W�[Mq�c�C��A���&Kof �
�*�&�V��<�iZփ��0Ǉ�����x׵������5�c-E��:�?�6R��W���>憐"�M8�E9�Fu�
b�*�:���{�$�b�b�/�)�+�.�o7��%��b���q�� �|:ƈ}_��k~y1�b�҇-
�8~ HMQ�ŗL��l���������: �;��O`�����v���.��N�f���Уo�̍Zy��]�5�
 ����.��I�l@�=hܛn���i��w;#��=z4i�S��O �{�� THD͓��H25�ibދv,�tؗ�����6ڔغِl̮�S��IH�K��#_�rO��f�w������5��7�%��tVC0.�O�|7U�$fd4��;V����J!ˠ���˭�w�Zϼ	2�EF����~T�v)	I���2������}C۸Z�:��R�-��������B Ӝ��!7xg.�iϊz,��)��%m*G�+L���p�����@����%��z�X��̡Q
�ַ�ȏ��FѼh�B������*�p�S,�/�����2G{���}�X읢��m�SV�����|��S�Fn�š�� `�/��/q�/ϓUCX��p�m��r��
������L}��bm�j��&:�����W˫C�2F��	�Ll�
 %�hz~���0�
_��;q1	j@�r��8��~h@=Wʡ]�(BDKܰ� "���n_t�?��N�F'm� ����a"=Z�%��*�&���JXw�f¨(`�i�4��(i�Fye����R��Mf7s����0-1�~kz���I���8k��N9F�$y$�%���Es���8��§[W��ϴX�������9����>$�7�$%Gƭ2�2��Tp�)�Q��� 7{Լ��{�8����<{ѳ�pv���(�>!l� ��w"�<�+�f���*L�/�osV_Q�-�_���O(J&�.Vm0\��O��W���u9�r)�O	V�`�7��SZ6_���#nRE]��1([���F�5�K��_�:I�M��]@�E�����jd+�:X�Fl�>�r�f��[���dR�'�AI�/w85�5�	��V'��ߵ쒢£{��$:�t,�8����$�'������G����2��I��b�t�e/�}��ҳ��l˝9q�)�;*.����v�#�ݔ�1���-o������w���YF��rĄM�����cm� #��� �`^�#�`,�K�c�yeZ!���*	��J*5����eZ��8�o�`�4K�['�T>�0�1�K�/��T��c�1��ba�HA�ZL�A\.�Ⱓ����܌6tѠ~��H7L�ϋ��A8kŘ>�բ���0�J˗�D�u�'V���8��6 ��CX�M����y����/�HC���<�#I��[\��P������ë?
_!�h����?6N�Iˑ%�:|��~�#��2�[v��	���̚�4�����W���نu�����T:����3!s�ˆ1�X�dQ�8ES�lH��%��Ő�L�~��,LĀ۝�M�� �͌��*"��H6m�Z �)�;4|�����&J�����p�zZ���nL�5HsOjI����~N7�r�����u�f՚.$�_�9�2\�n"�گ��*R5���e����Ö�O�Y�Po���\i�q'�.ÕN��٥�I��nM�OL�N���:hxm�c2t	��|8Ḏ�����h?g: ��{�ь����:",�X�A�j%O���ՙ�=�Uְ���=��\3 pD%�Z"�Kd����q���`}��%����|'[
\�ǌ.&��x������5Wk��?_����G�<Y��B�$C��[>���C$9ǋ׶0U�lֶ����;�h���'�3���zoˮ������B������/��mGv��sSqdHns��33S"ԛ�Y7%'�ZT�NR�M�4��Q �P�<��@������-��\�D~D�l��1�Pzf��Vf��5���I/��L	ǫz�����P��3�z�1�l�Q��L�UY2 Tdz9�?h�ϻB3������M������HRQ���v�%I����؉���GC����r������U���^Q&g��ϠvXξu��-��i��L�XZ�Jͣob��D]��}�q����_���Tc���s&#���H_s�\��r������6��!���8�����3���[��t�%Kmd_��|w|�^�/�~����Ky���@+���ޞl/�{�kIq&�8�\��5q����1�1^A\u����X�ۭ-"��ȡ�U:�)���P����Ecp?�r��~X�lq��+�����	�r�(F)��r��-v./��ܯ«�c�N0���4���ʊa��:�e��ZXW��0^$�DV����(��tӮ;�0��)�6���m��z@�MJ�g)=�����?�O��MU�&��]�;V���X�����{�#�F��J��j�����,�,�D���x�
b�4��3�oJo�?��B�'dj�ȜՔ���7?�Ņn�������SI�:��|D��eB�`��P&�[ZRRw]u+�'���Q� y�-��	$	�b��ܷ�>Ӯ�Z	���-
ȫK���9&0T�9J�WkJ�?<M��F�P��	�ٰ^���浻\��$���Ip�,Y%$�|ߝ���@m�ءQ)�3�Q@�hwd��>䜱1�hR�oYc�kx$[���CW,M;]A3��M������f4�Ց�Xf<�����+w~�]�ԘB�m
��Yɸŋ1��&lm~�6-3v4gs�f����xk!�׭cg�����!4;���1	|����D2�0c��4�[�=�Mx|@`g�!-㩁���H&�`��.��Ç��ϛ>�.����_�7�6�9��\��p��}�`,/��+�ē6�f�&K�G҆��"~^Z����>孪~R�>|�vD�:@�Ӂ�5�wo(jɎa~`�."�^�np�$�g��1��~���_����t��:-�\ma8�q�3'P��:�Ix��0t��FީȉW��q���Y}��Mоً�G���SF�RA8)=�I��@�Y�4M��.���Q�.2&���	��zz�su���6��ޭ�N��8�-��d�`���:>Y��2��y<�Ԭ�,K:�H�K>%C�pp��'{m��?\�3�J��n����R�9�~�BB���X]�S�+��*�Z�y����h;��@���2㍋�{7ʼӂܫVC�l�:�>��'B(4 ��Z��o�|��F�9ܧ�{n/�9�ɣ1Ϣ��g����N[6jF_rn������Da���B�$5�l���zef�-�K��\<��C��@ܣ��~n�����z�vO�r��*4��~{�P�JQ`�a�S�����r�R��&iJ�B8�/>�v�27:k��_�D��5���"u�����.F�K�eL[(6�c�H-21?��g���/�ܻV%��Y� ʬ��]b���FO�y�/��2��JA�������a�R��,�B���F��b���l��^g�{ѓ-8�N�Լb��$
3w����S�m� ũ	�bS&�+��s���7�����>^�L�$��#z��܊؋���s,�EH*������ՖaV0�S~�jb��^
'�nq��6
y%x��&�f�؅���,����h�J��AC��,\���DT,�QRا钱�y��J+��-=[�ҷӢ�h��q��o���u�Ǫ��p�B����ߴ-��P����� �s%�i���.ș#q�g��[M!k�1Q�g����HJ��2��|y������X �(k��zGI���b{$7���"%[�����i`�X-'���b���ϡ���3,^�`��p7܄��9���s�1Y�arP��0��	���raF�M��>?�����Vib�zi���t����*h&j�[�m)����6A���*�r� �,�Q� �� +��Bn�k��������F��כֿ����G����v�,U&1w� a���п�g���?:C�C��r
�S�����DyC@��3��!3��N�.�G�R2Dr��_l�~il�ٺ�$�@�3B(�B%�^�6Pwm�l!jŶ�	��� �pti��%{��R�'��[��Ӏ���!թ����Z���&��19�Q=�2O�i���m��$܃� �&Z!GQ3����S��x��	@��m�)Q:�e\�*���O!XX�6MR_�*�w �$�8�[;������Y�QƉ��1c����v=ʺ���C�lh�R�����6w�s�}ŕT��r�O���>ZMf���1�Lf-oG��Y"��P��ʂ��Lw� �d��yӻ	�|��c1��A\��� xgm�ի3�2`� �_���y�IF���]'s�%;^N��Ó�%����[B��!�P�Mׅo�����N������qĈfX��z�J�b�5=�"i�F�e�7Ӽ�&�i��)��/�����=ҙ>j�-VC뭁TFDؐ���*ߵ's�+��M�?f��h!�g:У4�*�ش���������Ģҁ�l��)�.;7�./9z��#i�.�|�Qd���bG&c�l��e��*/}霴<�v?J����c\��ȌAn��yN��S�e}M�6U_���nxc' �Q�;�����pb?^�@9Q�qRZF�:<�"ɷ��0q#�Hv��i��6fG���0�;��S��#�0@x
���b�\7����� p��2B�@�r�[�����l`ZFkEo��2N��%f4�,���(������0?0��K�<�3��@CU���ݠ�.u���4Ys��B��J�]�����eZ��lm��2�X����AfZ�Dg�u^�S|c�
��?
�n>�g�r��D*�n���E
d�#n�*�V��q���Q˞%|��4q��ڵ���d��\�\��oU�֖19_�q��V�7�9������Aй�ظq��F7�S���"w��d��5ߢE����l�>S�)`Bʟ����)���EY���Hһ�P34�?#|�!����nG�rM�����X3�G癈0�鐁i���o2��e����M/�@���z���Aԕ�Ó�x����V�Zjt_D����2���M��2�z^��L��nF����O�i0�dj�T���ĄZ7)�QJ�c�L9�*X٠Dc^��m����gJI1�!˴-A��Q%�[#���p5R���u�����9�V�?�Z|ŭ���9&�K���,_*'t�����F�A�-���hX�$�e�\+gv��Uy�����+^�6~P�r��ů	��E�ި�h=:�w�|Xk������l�^ۙ�|�%��zf��-}���� ��Sϗ�KVsU�W����C���P�<KI3���٭
����|�r��{D�A���*��0e�bH)����Z���Ko�J�Q�	<�����$�x| ��'c�8�"r�$�s��@Ѻ �6g�m�\|h��)'I[���B��J|1��}���a!���{D�Y�@��`(�+o� Jo����w6��.�ݸx8�^W���T��:��,�h�9������5I�ę@7G2�V�%6�Ț�$K̭�œ��!�q����{Om�B����:DˆZbs���JSa�������t�� SW���zG��ߪ�ʭ�w�1e�d7�{�X��G�7,*�97˒��! �eH�+sA�P�Ё/����]�W�� V���<P�sԸ��k�����1120��]�M--[���p/�bĭꙇ�b�$���	E��H�vX�{ө��"`w��#����d��{h�i�O�KR:�i\KL	9Z٬��lp����yg�;� ��48P.�$��PEoo��(p�2�����f�M(~��o�v�Z�D��@��؋ݵ8�������{�0/�-��`��1K�`{��*��[�{{x�VU��]�=�$9�������Kj�d�g)l�/�́���o�G_/,��ͥC��+ڂ��A�5]����KB�{�0��QJ)n}�9���rr�Nw� ��/���b�t�Ɵ�?k��{<
��ࠥR�C�+��gݖ����?y�<Cy�7�;EmJ,��A�5�t�[��3�:R���ß�P, 9����%��~��w�;�j�P�)�R����G��kWcXNt�bYp׏�\������q��$����_l4��|�c�<����7Wㆪ�,h�ڷu���W"n�E虭U7�I
�<�cg�����"���|���N6�M��UT?W�s��_�BAi6z_�!MC��o�����P�U���(���8�~k�S:�,�@��;O���"�`��g���oʪtf�~� �R`.".
Z��e�'���L".����P�mn7\<(˞��)���k>H��6�l6!D�����i6ݏ���]?��=��?`���2V�0����RN�g��= A~��6�E�)lR�EP.�Ř�B�~z������$�h-}.m���horK�0}��:��{6�Br�2���A��a]g�����Lʻ�z�f-�V�S��$�+�a�d�� yp�p�iuĝ/{��nUT���ۧ-FJާ�y���GJ�l>��Q�lJ��-ӑ�Le���S2�yI�?F����%��ŻRC��?E�;��Y�� ݧJ5�����M�|T���Xs�y[E+�?��eh���SAH�;���z��և�?����~��H@ekN���B�31)��:����^G�'ٿ���V��\�=�a5מ�j���o�=2}���=�w!��;�
^A{��d ��Sc���?�Q��3Y6����;7
��0� ���E��I�3<���'1�S�%�A��[c�HS�Z	l��
ׯ|~����.���%t��i�_.'6�A��nǙ��{Ê5�$�����d{�����ž��ƥ.K�n��R�[��G�^ݎ�՘�Wˉe�N�C�Kw!�MvS�J�$�D��	-���a,��!�o	�<��>�@��pք���K��Z��	�@z5��؁��kΒo[��Z{D�8�0.��Cо���+F}{q��.�E�T��umav�C<��ֈOO֖;��'� }�6�$�c\4^�^M����,���պ�STH���ߟ��f�W!��=���&^LaEtș#����M�ɚ�F<���ta��g��42�,�������W2��#����F�ؐnE �y��{�N�_��7v��Yk;�e�d���~�n�����	qR�����}�҂I}6�v?�M�Xij[�@���%�;��'�`��b��_���b�JML�K!Q�"�4	C�_8'Ž�M$Nî��gl�E�@��I�#�gmXc�J5�Q�H,��4���Bl6����TT��5y0: (jԜsc�5���$�I�وUr���zћ��ɭ�ɎD�ۊo4�TwjU"]��á#��~�0�����.�a~D��0yc��Έ2O�Q�z�Q%_³r��)���G'>�76�w�R�TR�ߪ6lP׶u�"�u�{��LZ{.�{�6�E n�%q�鍵��5:\��)<��0'9x.�q��K1{�3�� �Υi���+b��4����7�<V��J�ľ	�J�ku�*04K85HQ?�=�f���ڎ�EsAv�Dg&�H�Z�	�Ĉ�%[(2�oT ѷ�u[)l���G0��)�s���p�=����z�Uٳ�@��s��>.�T����ۂ�l�/����ū��Y��������=wT�R.��nB����Ϋ�k���2������F�XT���V�R�ff�|N��ܫ\���� �^�h{,�i�]�5��o	�ɬj�&gD�}�2(6�
�wT�ې"���qP�-�!�xH*�OaB���2��hv ��䆤i<���<�BH-��7F��*�]Nt�{�Z���`��������vy�Ms7	O�&�Dd»n��?��Ti-�.���;mX4���R�Mq����UwB��|V�u>�q�t��'��X�"
n�;]r��gM>�G܄��8��!������W>f_L���/�ϫ��ٝ��k��	�,x��8�:���`�
��OL�����,��R�'�-*�x�$��wŔ|>kM?��F��r\� �TM�Ɨ��8
�N�Yj��S �#�T�B勗�W���d�4���m�l�Vv�m���6�0��y0���^����v$�����-U�U|&d�_�W��_�J���0hr��F��u_"�$~"A� M�Q��A�������H��Ff�Gk"l)���y�څ��=���b��BP|}����A�Ɲ�wݡ���:�22��\mnA����ha�K*� [�R,f�a���ݢ<��G^�����!�Z�-oU�D�j�/W��e���U�w����\��.aI�׸�
�090�5��d��¶J5��~�m�ȱ9
f|�u͚-ǂWP양���f�N����Dyx�I�h��
ԝ���)�q����C|�\��Jפ \��tG3P��{l�d�y�Z��T﮾�eYf��eAF>D�Y^1��p�6�2 ��ht��"����ю���m�V!��;B�
�up4�HIn�t
ɲ��MT�������i�#<���x
�/�|��{jמ�»�+G*���*\��^��|$'��}(7H������ j�(̢&;s��VD���t�I=@$���u\�=�&dc�*�j��T���J�6)[YΣ��h[�1b��pgN�����9~T�M�Id���-�/���jM�9h�����,�*�.5��d����{~�%��xf�x5Ф�m+� � 
�f�hJPq�0(�^��4S�h1zY������B㘈F*�s%聅&0��Ć���: "U>���o�-����P��i���@ʟʴSl~�
̠4��&U.H��t�&�pZ5�ڿj�(�qcq�Yց���[.��M_Z� ���WD-���fOjDtR���ϵt�o6��2�&��e4E�YB��5E�h����O�Xa��}c�LCX�A�e�!�ݺ7�ZXd�7OS�.6�3�g�Z����`V,0��$�-c$�#=id'�rV�楝G�I��z�{�2�8X���7���$�T��AŬ�
�򗝧�X<v��*Lj_����%����]h��e>z#y?V��x�S,AdH������K��:�^@H���rc�3�_�����T��l�/��6+�p�Ӌ����Nk$;�垖[%�0#��[Q��y��7�;P_�A}��nb&_����lk�h���Kx��uv���K�	1TnC$���W�΄�SI��[�7�cgR_��0�k�J���4�)�f����h���1S�N��y�A։����6��Y'%6A-&�~�K(TϏzkV��n�u���-[�s��m�t�0x��s6�o�«�	7P�1l�t�i��F���:t��Q��i&_�J��(��>+1�gmb��u��q蜁bS�3e���1�ar���  ���d�&)�۴��qKw��w?�}K(_��auZ|3��S��`H��|r���P�hi��ޟ���.m�:g�ˡ����d*B�	���DrO��	)^q�G�|.6+1�HI�Ǹ��A7 ?�N�H�M�3�2%B��M�?�y3�"T����&k�EO`ϸδs�o�Ry:og+�/ShH)_9�LQk���E/Pa��#Y����]{&)�~�Fj��F���<��
���z��_��K2�ta�S�y�_�_l.Ґ��x	{B��91_J5�%�C��o������$X�s(�Ց�� �7_�"e}�T �1��`�3b�`���MP�c�_��)��ʤy������S��h��/>�#F�
tsvc[��^e%=�[s�l̈���q�\J��r)�%�;��=��>�w{#��ZE�n�7]��He~��A��ǂ�}�E�?�"�Rg�Њ�Ш%�L�RQ+������"�6���|���V�쟝�"{��:0��:v-ݤ��ė"'��]Չ�ȏ�a,M�
f���tx�8�R��>.����c|2%u���X��d�uj%K��A�.=_��C(n�c�7��Xr�f;�[� �J:����19�h���-ۀ^�
�].��P\�ʠO��U�����M�ि0�&x���t2�O�ZS�Dw�n��v�����9:o����P-������`�M��(��ϰ����a?�g��O~N�h�;=��=��I]�W��?]�σ��ÐC��j��$R�d���{�"���|B�O�]���j���
/u�B���' a�SS�d�J$�u�F²ES�#GAΑ���Q�hM�DٵN�#�T��G��!��6G9̇���)QRl��<7���f�]9c�͝��sx���+��y3*�V�sn���홁z���Y�����^XM���Az���|,>7�tQ�i��\(+uX7
�S�F]��
rZ��c%-`��TB����e�Z0Dt��:�F`B;�)�{15v��dC���1k��ga��:��i!�o�-'kF/��D���l\��c_`C��O"�!���e��.IgZ�H���O⦽�TE�&������tƝ6��� �CFk$�e�ۯ�(k
����11M���&p��=�@�!��>�e��p�V�*�zQ��A�#{Z� ���:��֚����A2;A�.�	w{~���R@(~��p��e��NF��t|�R���pP�O��ax&��D���GR�W�ѐ(	+e�\��"^�-��b��U��-$�i��ׯ�'�V�6o%�w�������=M��Lי^P7�̒�q��~UϾ�⛦��3�dgT�BNon�"��|x�t���~,2�`�Bi���G������
q��]0�������P0iұz/��{
�3�f�g-��y����0S$_�O@�R/|�6�-��\����Ѯ~�yi�P����8�R�+�a؎�5-f�1<s�>$G�Cj��Z�O�34(�������^*��bb񲾀�Uc�{.�,N0�s䃁&>��9	%};m|�w���P�9o[hM��.aۢj��[;��K�X���9����,.%�Dn����4����L��P
��/^���D�z�*�I��4Z���+O�%�[#ĈXwa��,Z7��l�]�޴�Lu���c-�r�J���z����$��u+�!Q�e�rM2n:�,���"U���*�����#ہ�� **|�u�7C.GnX������8��(ͷ�9Y�1,���5�0|�5��KD�<Ʉ(,�kR� dj�u�]���"�X�= �f�
�^ۙ:�bʟY�/��)��ׇ^a�Y�I���L>i�"���.B��6�n$��3?��5�u�ﹸ���1���*)�>U5�]�W���y��H|xwwL������vꦩ��B]���ME���8D,��;�l�6��4J���s����9_����؊����xm�qh�e퉙�X�+6O�.�-9�^ΐ��q=a�Qw'�	+ߵ�@93HXzR��(�8�-�<��㑻���#���$aң�{,}���$��|�zC������iE.���(pN��:��<���	`Cq�-D\k�v4���Fn��M���#��@��s�*�k�*]����Y6����^� .+�����_j�x��~���?l��ܰ|��:�k�Xo=N�;�cE�ĕ^sL�=;�	ϗ��,�fҙ�֍�!rV�m+A�H��TlGNy����幨q��3��F��,UI@�u��x"^���<1�X	���y_Ŋ�<Mc\C��)�ѷK�M. o]>��<*�04�,��y�M�����a�nI�ﯜ(F��_�����S��6U4��,��m� V��jR5X��/�y���^��"{m9R��$�t��U��ԫ�#���
�>)`X�������m���~Zt�0	�<0��-�d�e4~�h���4�d�� �y;����v��O����{8z�5,�N��l�eX�F�/�@5x���+bF��w�i�� D���Mofڅ�dy�wհ���v!������$:p�}���0ؼJPO?���Ek��H��*\0��N�m�}�ļK�����w�h���
�7�W�rKdj��	��VRI�����s��fc��Y���M��u�=z3þ�2Dg�~���!������d녂���N�������Ks���A��ln�Gm�(֗iJ��j��D�egb�fc�_�x��7t��L#�!QnY�0٨��F�i�;���x�/���&��:o�lK��-QR�>Ut#�ɐ���<�7��?!�lO��WL�e讔ʯL���5�$"=L%�x=+2�x�mE,��v��U���v��V5�BL/��ATˌ4��?�1t0$��3��d��~�A�C]�[+�����Ӗ��5���>o�g ވ��nP�����ɚ;��ݢ/Z$Z�S�蔧ߝ�8J�B��#k7X�_6wJ��W�t�.5�%�hN�te�q�K=,��
Dd�`���3h���$�S���x!�\j}�ﵨ�i&t!U�) f�f
���~���(�^1pT�6e���N����WB"�Y1{����F��|�K�Dn?~��H�s�6c
"�P��/P�����H")���~�C�f8���9r�s���b��H���3[��������Ǭ=_o�*I���9�s��* �����5Ԁ��������2����a��A�9�����u���k{QSx��io���P�PP	���A�11��$|(�d�1�嘍���+y�S�����ő!�>�=��V󲣱����?�˗9k�.*=0�S�o�7�֍J���n^;����K {\����2�E $�t��rt\��SS�,��Y	��צo�lA������6"�ii��H=a����#=)+/`k
7Y�[��3��������|@�Z��(�E~7ה-�0W6	���\VTν�X	t���I�W=�0����B8.ڍ���	��3���1�z˽珆�*�8��v'�V��IG!��O��TDO��eM�`��ɥP���/��2?��L����J� �]��C�(0�،�J4&Wߞ^<O�lW�Oj�������Q��Q�𿞈hh
��~;����T�#*w��n��p�d�܃�W���a@��ޠ��l~7i���"�0�=di�Ȑ~0�)o���b���a^Y���F���?R�B��m�q�7���e�j�k���a���ȴ���,o��&
7�%�Z�K�u�k�ﷆ�V_9���u�����5{�5��hy�hHu�N��f�u)�6o�8�땭-��{1�rc�H�����vmG@9��0�o�o�k#'x!��xKE��� 0�h>��
�]������\�92��)8�	&1c���%|K��
���4&r�0j�7P'�Ip&�:�%�b49��d�f��X����e��qlA�U�W3��+=,�!;@y>�X�`��	N�ݸ��"�}�vXjj`��G���xj�;B�D"v��٘��n���g�Ƚ<Q�U��E�]r�vl&�}�n�+�$B��l�6�8#jC"��j���7��əo;2�U.��{	��^ef{D��@��l��f͜smwC������9�L�ǒ7�7���^�sJH�1��}p]�p�^9qzI}+
����BR"Hes�?B\��|_���n�i��G���h͋r���R��=
y���Sx-C��4���-��>ʧS���gyb\T">��^�2b±#�p��
�Թ�"F�c=Y?	'������l�^x�BQnF.``�#�LN�Y^�'_����q'���R�ie!�$fx��vg�&�L�����ۿX�Wa\�|#�a�����S�v<��F�5{��sU��>j#��8ߙ�U	Q�?e�]�9��7~:�B� Qs�� '�2��h'�i�x=k!�-!�����rE� ����m���˼����c�l<�8$T�/|P�p	�a!���o11���v-�%� ��O�ߍ�sX�}�1Orڦ����L��R���xe��J9���Ѣr������ͥ�����A 
���@���1����L��M�ͺ�
)�:<%z�����29��fe�{��;���nz��v߸Fw�>O��q�F5~��%�y�t~%�D�ۣb5��v���X�&{x���G\yj��.�M��ؐun��}���S;gAF�t��5���[nÛR�ЇE�'G,�J5|BFh7����r�J�?y*n�F����Z{Q���Y`M����i�4���L�-��G���af�q�n�{%.��H\qP�<����[��g(m�Y��ҍ����o�;X���D��,�h����o�H+\��5����B v���`GW��EE`E�j��1��,�;��qk��s�b�SH�ܚ.qǉ�4�n��k=�o'U!��hvDv��@L�oT0_�$�on���gU��bYŷ�Pz��%[tn�#ɳ����Kik��X{EHb�7�h�L�p*�s{��0/� ��o2�ǈb����Ֆx������**r�7pM4eԝY6̭z��__L��te�;���[G�8Z>���S?��֩wck���	r5&��A��.؝�.����zaWg�6~h���SN��!L����W��:���w3�����\o�����ή(q7(�:`� �����|���ɍ�#Ʃ�4V4$��+�ΒҮ�cX~5:[	�h �-��e����Ԑ�m: ��SgV�O����4{�3�Ja���з2!��]���6E5�7r�4�� �e;�R�$�kuЩ��qK�MӦ�Z3�;�������� V\�cm�!�Fв. q9�J����\������M^Gu��O��WiM5�ن��0w�����:�W���yY�𡳹h7g)���\c��f�[2����a�%��v>q�3^ٱ�*&.R㗴~�9��0Y��Z�\�����sk!9��(b�ˎ�d��l���d�ʣ��3.8x;}vV�M�-\!��u�x}.r�b*L��e�p������抄N�@4� 2�"F�T�M�:uae�]Y,�KU~;��&��-�o�$!��� �
u6�bЁ�Af�
7ܱ��^�݉3
P!1�#�D�r���~�wMyP�U���0G�:�{Wt:��|�_ǒ�m͢��~���v��N�x�A >�}G齑���iЇ�{�r5�#��I��(nW�+!sbK��o�<YZ���\v.w��E�r���׼T�2K���!5��qJ`Ա�;����K��~������D��)��>dϼM�	����M�ζNz��o��f�B�]���ʦ��k<������u��)��b!Ƽ̔�d��q[BR<#1�K0�x^�����C�z�V��f�������-L׶���;[��n(}g�Fٛ�[�*	r�m���EĐt��C������|q�"[�i�V4�m�q9�����`kḅ�c���AN��of��z�	�@�Z�W�N\,��¿��gpV�	 �ج��������K`��v
�t����H	�'1��j��n1BO�-o�?|+�C����r���$#�>�hkH��wL�ݝ�g�l>���#{(H-�A�,,p>�$ɲ�L� �mT�G$ltI�w����%Su��B �,�{��hB3�M����uy�! q�z�Ω����;3o����$K��G"�	�gU���BR�?-�R���4��ܕ&�ȶ��p��c:K������n�xv��F����)�J��w�`�z}L����.�a5����YZ�~1h����$�Q�Q� �N��F�K�>_E��l�]����'�FuI�nH����o8E�G;^���: k�,��`��6�> ��-���E&�<�\2���Bh��ַ�y-�a�Z�H��3�\���<�:v��m=�E�e6?�.}y�ybLS���~������Ɋh	[K�@dK5�|�)�
,\�4���̗r�t���ޔe�`�J��|�!ڼ����vP�k1�0,��
����èx��w9��p?8�t#x����[0��^�G��g��@�g
�&�'�rk�R7�0#��7}�y�)X<sZu�z4W������<���x��A$��@�\�l�_��Y��L�R�΀-�U���m��ѓh���� �!�M[�@�]�L�v�k�V����]y� ���"1�O�茥?ԁ�����8u�s� �+~����n{ꝋW ߌ%�3�H��׹*��[Ž��۽�0��|*��IW��0�3�������Fe�_����-��o�&������c��HD3x�o&�̝%D� ��鏳������;�Ph�	֯}#}�D�>8x��a#�݂i	*īo��e����+�,�%O�E=������I<�j�~�?lo*m�9��÷�:pz7ld��B�ƅ��˴�!M*z������8���4�\1�]H���>D����]l�#�&m�F�+o~��%P���M���M���?H��4�ߓv�1�$� ��۸_��s�����{D��-���܇K����Ĕ��u�pR�Q���_+��9 B�^,=�DG�9��MZ��䀴�f>�FH�LKX_���*F�y4 ɋ%�U�%&�I^z�1K+�}3r�F�<L��݆@o+(*W�h/��ՙ�?p���8W�U���=�F��=�,>�t���'�Z�O�o�����{bj��E]lԒw�}q�P�!��Қq�>[JZT�N�ӟ��&ԃ�b)�~���ye����bh��`g�iy���X���t�م�UP��hd�z��m��HA���32�sv��AIWa����;��N�N���j&�
S��ZC܀!>�Z޻l�m��_��8(���n�>%���0�޺-_�{���S���;.:��j���ْ�$����9��)c�WBg��얘���apt�S��ޘ*��U%EpG�j���R�������O5ש�� *��/+�S���3�5ک>���}��*u���IY7'I?��B��|Ё�!����� ��!��BȒV6��$8a���C�	`R��ן�ltv��4s��e�]��Ia.�q�(���g�.R~�%H|��<k�\�Y��i�=���f_O�t�t��q����˭��v�C�:�qÓ��lP"�������`o�`6 ���T��]���������Ѫk��D�j�q����D�{�0�O
�|V�]s�s
k�h�����sI�V��v��=��G
f�Fo���lԱ(񪁳LEkKȜ��+�����<�x0x"E����\;"]��Hݘ�{�
?m�)gEmн�;�±����y�h�Ĉe��nO�޼�{�J~���a��hT����\_J���Ԃ�M� ��A &����;��*��6�L��?�J�xfv�|u;�c:�I3f��b�]���{�圮�	���"����%]��+��*>�D�!,�Q�)�q�w���Jƾ�=wjT]�����a��;W&	�yj.^7�*�9�����a�w���\̲�ԧgKj�w����q��Y%��@���G��i���֝�����d�?J���%)�L���ba��wyJ�b��3�_T�brcؠcD4o(�xf�5_��ց�D��v�?�*��'��QCq) ����aW���MH�3��zR�ݶ=�g��$\�?�s\.���m�5��	�(Jf*��A(y��2S�L��*z��G����z�z���ӈ\6�F���,}�j���j�QHq�x�6]�`��^M\�:�����$%q���A-^�5�@�ծ�~�h2�A�i���&r�it���
!�[E��� ���!ݏ��?'�hOI��y��1�^['��L;Ֆ2��@g�v��9���5&��G!Mo���=�w�������#��e'��T�uGby��'��ߐA��؊�����~��(�x�5��Ҿsǅ�/�b�NX���#C��B_N�����x a��)N�O&�XT"Ρ�3ݩ1�yQ�=w��=�qX��M؉���,�}��ѡ6���$lcAR�-Š���[+48��F��jy�3�6VJ��V3	ū�����\�z�)�B�ɧOD���5�oyf�jI怺�B6k*���B����(�ge���M��tc��
t.�Z[i���<���p�˙:�}��|���M+���#�fׂepi/]7e( ��q���}�Z�H�M���ǎo������8�<��z'm�7=%�*�ɤ�M��p�:Y]XM~_0���F��:,�o��,�+�Um�8�7�kH"��.,X�����:���:�ל�Hb',���Z8�˳�k����6�߽fx����Qb��|�86IEe(d:��`�,h���ش�� �N��s�?e�!0��Ą��3���Rq�S@C�d+|[{���2z��)E���*���4j�6�v��e������,YD��y�2����d��f���������V�ai1*�����Yk<��0�?��?����=]��{��L���4��ѽ�J��w�����B<�&�IOٓ˄O*X�x��sK��������@x� 6<�W����'�S���sZ>�$����M�h3ט	�;�e�ֹ�	��2��q���=`4	���IPqe�P�1G��2ɹ�Ռ)J�~;qu-��P��b	�\�R8�:pw�� �`�"��E�~v�r_QL��4�勫A3ۄ�"�֪��T�2�znD��!���bd	�'��}���yM"J�vi4��0�U�!��
�P^��И7;���|S�Çg�z���E0�Üog�o�1{�$�fq���Y�᧨G^���2�i��H�I�t^��5�E��+��ϖao�r߸�@yτ��������}l���Kc� Z���'�(1Q#�������$��~'6R�,���J�8�7'S>� �~7
LΩ�#��F�M�*ϡ�nH�����	�!�a�S�E�
t�E7@S/�1���s�Q;�F�^�;x��:�"�������F=,�w�H��(W���3��Ť����U��G���Fl �Tp����?�a3q��ީ�7S��S$����I9��:�u�Χ)��ĵ��
��X�41o�w�l�-�����	�6�:�>�ՖM��0�*�ƿ��-<�M����$��W=��A	���? SȑVC�t��R�!)v�A6ʝIc�B�:$(���}��,�{��S��V��5\�/yT������G�í�Y?�t�+�TJht8�5��<R3���Q��	4P�4��hGF���(��C�W!�'�|r������}���ήv��ʰ�mB�	�i�m���&I)��; ���f��{OH�Sҥ�3m�j|���N)���$EeW��V8�&úu�nF{>{fy�4���GR,�H��;���{���؅�'oG�y���R�	p�Cݤ�e�����q�s2�*aߧ.�������$���~{����f_���^^�RH�N׺)�0E ����eC�d���у�gn�6��e���
�-��n�����!Iz%Ssu�A��z���E�cUb'`�3Cb&�� ��+����q5]�����M��l	���������X'=�qQ�A�]<\4pޏ^0Y���{j�>��s'u�MLv���)u4��Q$�,��h���Bǵא2�D�:O�����b�m9[�R�%�i����/�g��wy�;s"�Jz%��l��~�ԃ�ī+?c��z� ��Yu�r��2ѐ@ȗ��f0���u-�`���`�����F����r<U�VD8���H��ĎĬ��ʀ��&���t�Nd�bh�,��)s��'M|��T�����n�s�)�,`��jmٓ���Z('����m��K���R'H�jt�)��������/ɋԯV��d2'ָ/����
n���+z*���j�ȗ'�nT�5X�_|l�ȍ�7q��ы�g}�W_|�'���c���+�&�!]���l%aޯ>�ޠ����H�>Hmr��5��!�v`e5o�;��ѭ�/ׅ���mmZI4���=vB�L� �s�N�݇���q8��)�W�V���;QX7��`�+��f��~=�!1� d3���`�Ӽ�u���j4��4�oFG������fܝ�Vo�|��/�FLt�(��h��Yq����=�@��c@AO�)�S3���4$�6�)o�B��(PW��`�X�O;�S�̚�yT��Dmcβ �A�ˈ��#"�ɐ?&(�H36}&0L�KX7�T��5�B^h$�猨;XGz1ˊV��̩�/N���~6!���ckn�*�Y��ο���{��d��D٧}E��TXu]
A=����u@D�Ƿ��Ϗ��U��ǜ�fR��Rg�ࢋ��9w�,��Y���rJ�i$�"K��Wp��B�q:��{ι#�9`��m�?g�gu
T��&�|�W;����@b0�HYC8��<��zjA��$�?�heA�A*�w��/5�r���$�^�26��.��9�q�J9��i��_U�	�X�/���5q4�L�0�,���ұ��]B�h��8��R��Y���7�9�*~�VT����X�J1����[���좙!�����\Q���ʸ��?�!3ܥ|�^�5��uZg���l�"|v��dȧ����o%��Z�'a&+�K�&%aLˌ�X�T�R_�XwԾ�au�om/Q���u�Y[S�"�I� ��d��)d�m,���F�*�TshJ#����O�Mʐmlwv�ݳ�ko+��K�oE%���	��4m�<	��
�kx�-�ҍ2<���qA2)���<�ݾ�xS�>�,�ǚb�kX�A�D�nt�������jK/��7���ɯr(5�/�:��~����N-�47�dp@X�e��j�����}�ޞ�T8lK��zo�~g�QbZ�#k��3�SM����0�ݒ����Ѷ�Ht����u_F+])�v]J�ԥo6Ɓ�S��`�@`��-��#�D�>����d�z�7V�u_���Wm�G�����n�2���1P8Κ2��@z��ct�?9z��c��GK�����8�WE�� �u39�7������ d��L6z���]��!�}*w�nK	`<Γ�������	�\�ָl��-hY�.�Qv��ƅmt@r7��7�b��ϗ�ri3�K��q�:�
,��F�dxw���w%�Z#kK��t7);�)=�d�/A"z@pT�γY�L�f*_�6�ˇ`{z^���$HQD�B`:��eYe1�@[�7�M��l$�;�R���E6h��T�'� &�c&4TP)��RUC��� ���z�o���%^��IlB�pX������`����s� ��|Y,��&��oV����a{�֏c8I��+����S%�n�JIN��-��d*����k���R]׀G���܆��^�����f�͝+�JN�u7S�jH�l�+@��ɘu��ay�56΃߇(�c�4˅٬HgLݯ����s�Q΄�w��Sz���w�HO	�o����) J	�n)iw}�.�rc�.�h\�e���
\l�8ˌ�'��2��7�Ɵ�5u��~O! �4��g�E��t�>a��`+�{liѷ~�ѵ�����UXr����y;>��<��[��@T����}�`�r���+2:g��%&+���?;*��� 8����h������$�?+�R��1���)/׮�!K�rS�׆J�j��k��\�_���pK	�F)S�p�����/�]��vn�ƹ;����T�
�����m�5]X�������|Ϯ�E6�4u[��m�t&e~:�xʛ�����7����+�p�C{(���	y��Ȉ������&0�M�o=9�a]��h���Ff'��O�
D�@�"�1�}pv�LY24�H䍿��y �n�� �l����5S����hG�-��H�@[9��z��*�yz��+�K}�B"�H�Cx� ?�Ԇ'ھ�8|o?�T��@�*>�L^�!b$)��fN������a��Qu�=�0�_nC#�m�F������!'�A��_���B���4��F�979��1c�h#�nˈ��������OJI��!V����0��d�a�Og������ ��Gڊ��VX�+�Gb�8ܚ�я����8$(�Q�Y��=��qVo��Q\yZ+ r
6�v:�/l�fw�e�'<�ɬ�h�j���� ��q�V/�L^pXLp힨D ��G�/���s�[���9�R-��}��<�bܟ��o�����ǰ�Ϻ1���gg��&{R"�u�����zif�s*��� 49�{Eچ#����|��w:S!������3��;����*�pUM���b��y4KtV�s�a♫�c�Ʀ����se����e�t��%�!e�:C������/	H6�_3�Aޫ�pb�g��c '�]ZUL�y� ¹ǿ����!U�pE)� �:Ө���\D�x=>/���G�9�s2z��sߌ�9+�|����D Uߥ�6�r')�~�`q5����c���|��@�ɲDt�J�<�L���M?��إNan���M�����t���;&�H��j;}��ۺ�)P���@2l���y���Z�=����ٿ�#�Jھ��O�P�a�6/e��`Y e���y̥�����&��Ɉ?��y#%3(�L�6�:�s1�e���C��� 0���)�SZH@?��U��9��0zf����7	="Zע��Hk1���NN-r�EO���E��J��� �E���U����)�� 8u��s>�撈k�f��9��"��o�~#>�����ʠ<6tj�B6�����r����D�XAD9��z��1�brJ,gF��%�eT�Ė�z�c9�h%�F�K�e�_�s/���f�tA@��=�[��i��C�iMys���Vۉ��K/�_����
u9��9[H��?ݍ��w��s��D��r���zN��?��Zn�k3ѼE��BBH���[�Fo���֕�� 0<��W5��nr`�$��{�4�|��R�����֖�9�UZ����K��Q9�Hiֹ
O,�]k��#����{q���Y�~t��--���؏�H�N� �j�_��!Dn]!%u��W�4��QA;aA����_�����@����}B�D�:c�	3�R��Z2~o�m���Y3kj�nx�|J���1'�O��[NU��N�T@f1�{Y�8;��؉���M �u?3Af�n)�42���x��2���&!'�!@�Z��7pt��hx��'���3%MG��8�F��!��7��1�٪��eߟ�o�O�n���^���8XԂ���Ky����ӵk�NE�)d����p�$h���%9�(�7숞,��+���]|ס�+P{��L=n:�a����UY�h�k�2�<���ђI���P�,�_����ɻ���,�u�\�I�^U�8�gbʑ��anKG�JhϴlA�̀p��\�k�j��99���4���{�m�v�s�ϯ�ޯ�V4it��̠�,}(�7^K-��ԘzfV>�jØ�rq2��0���F�խ���8cJN]珞Q����Cgf���D���q����+�;��D�>�Q@�#8��W�s�V����-"Ϋ.C����$�$c�R`}0ɬ('TSU�u9d"#����=�s�&�9���ߙw�J#�e���6�C.�<�af�X�Eֱ&����������쮇���w����@<��~7���Q�,�b;�\��N��3�K�X޳�c}� 㚬��s�K��0�5@Xׄ�h�Vb��Ku (ٶl-+��)���{/P\����5��tߗc��-A��k7�+	>9�/�+�i�d*���s�O���ؘ��<�&��=m*W����0��ݧN��<z�(���j�܈���🎈W�d
ogrxS/��l��Њ��N�T���mC��<bG%����#=ט�Z���A�Q��� ��#(�k|��Z~d�� ⋡m�M-�߼l#A��;}6{,�m���,;8*���$��4q�Ѝ;�=�#��o��E�,�������,����r���
{�f����o045'A|>;c�?++����P��z��y�G�~s�>�h�w=��뮎���+���ڏ�D<�$���I�)�����o7���EV%�ݮ�KU1I�����2gM�u@�LJԋ�����*w�-��}�]�d�H���C�R�Β�� �$��;��7�l�	�;�2d�?�	���d�y+	��W/�e>�!C�P���ZU	��(9�$�����Du��D���V���G�?�k��'KF�]�2u���q\Ze�ee��gc��i� Aj6_Z>�Q�F���j+���V���r��5�g�Ӑ��}W$	������W	b{ª"|�i�t�o�c`7�˥��-_Ԯ���W�BL�GҠjr����KF�di�<��G��*~Iru%_M#�-U��	�c��=����A	�V�8p��<sձ��84=o�ʟ��Gfӽ
~�������=mO��}�����\ۢx �[����ZX)�A8�tmx�
0�2b�s�5��nP��yk��(��c�;Ot��h?9�ٗ�Wn��Gl�D���b$��{��JqQT��	҃�Cݠ���6�/J*�M�_)_��~''���E�)r�2�rrrԕ�9��������s�r�7�$l�-ۦMJz���eA��hm��p|_U�{D�������}����mR�@8]�+�KX�����
��$\
 �K�@q��P��2��n<���!j��g"�2وW6F0����9�tv�WE�g�"T�� ����ڶ컉��  ̋K�40
<�s� \�L>84�*�-�PQ�~��RG����t�d�L���)*�y���7}�l(��	�B��\"�?/���g����偯��hjS��<,4��)���s�7�u�r�k��Y�nI����-`_��5w�_CF4P�u�L��ܲw�*e�/�^v����f�D���Vs'#e�U%��\ܷ��cSS��T�,t���'Ù2c�G�D��ӹ��g�q�.<�2m�����z
�ڎ6����
�h�v�ljW��<���!RP!f�+pJZ����F#Vy"�s!r_!T��F ��`%�t~���N@�lFg�H�;���U���0��j�qf���8 L���f=B`Y�ExWDĝ��|�H�4  g�{a�"�32ںn7|yݑ�]BV���ms��u�9Ƃ�1�ag�Zְ.�R���o�I�mS��4�vy�j�u��<'�������@� �+M��%��[�y|K�b�Y����;���!7TLŏ��G^�)�ddT5a��>��4\QQit���8�g�NB�4p��1�ﷶ)&��hp�@*٪V$!��$ԙ���bp��kd,_�h�i�ܴ��d�dȨ�����?���-.��;#�'�����!v�Z_q3�� ��j#Z�0��qG4�%2����BӰy_W3s=}�Y�Bq]���z|i��y1��`��;��ml�5$�>	������Y��
oI�y�;I����;$�ED���Rd�|�@�/� �l�"y���B?Y�[�Q4���C҈	#a�O��6f�)g!�d�Q/qb��@��a�	ͬn�jzٱ&�'�e�q��g��r�=��1��"Č�	�w�l�ۼ+"�y�i��������5Ҫ/������!h�;#�Q��>���*=�Tc����!z	��o�ڭ�۱>L0'��U+u��/r��#UM�V����խگ��.,,���gC�Rn{�:����0�;�!���
�*��Z(��x�� )ڵ�&`W�Ѥ{��S�D�����V�G����gUpR�%���H�i��2^�~@;�H�P'|1�[f�����e@�����LlAS4�4lY��̰��<㿌��6���s�r�u��`�C�6���Pe�]��\D̑�����VE�纕�R��	������ �4+Ke�(�}k�[�R(A7���(stV�d(��.t��1C��7.A�w���qFO8��Uȅ[��z*�J��H�@xR����I�G�}�l�_3���m�5{�zQY|�%�kIz�6k>#[�Rc����dJb�_����I�7OehP��<qt�뎦�3�P �l.i�>ɜ���x�3���"������:"5]:П�H���D.�ͻ��,�����R���ie��y�&?j��Oj�U�<E.�a?9g�^Bk0e�;��K*����V���;�O
����%z�t!D����3� ����D��Rmk���O��掌$S T? [}.F��D�Ȣ9\6�oO�[�k�"�7Tͪ���j�2)����aq��_/�+�+1}�x�䂑K���h��L�����}�,oK�VuiD[���i}Ԯvr9����$k���j�r��@��th�O�D��?y1M�׶��������P�s�O�qL�:N�B���i �����u������N� �:�[ԛ��ⶺ���x�By��_����zĒ�b�D{i��ao<2�~��gQd�Yrdn_j)�s)vH���I$Y� �#_�Mћ���حTf.�82���L�9\���7���Z~�Z$�f#��%��]Ho�af���S#-x~�cSP־\���k��#ͬx���c`&���t1�N`��t�H�3��4ϱ���Ev��<�`��<�z�&�e9���66����ЄwА/>�
�̏Y���L?�7�Rҟ��ѯ�
"�jT�3���wi��E_p�zR��N��n��H������N�'êH��߷ȋ�Ra��V�;�1W�x��k��,P�"��ix�zx� �C����;&�!(�>���[e���.����f����}�ݛG��v�$�2���:4�V��O���|��%�����8��'�2,��%,6��V�:C�`C���$$���I�e�b�N�)��!k��^���jQ��[�2���oIe}3ߚA�h쭈�͵�zh��C)�7�
�l=���E�D�i�,�8�:��$�u�e�Bia�
��.9%o��6���8obƯ1���f9��څ��g�M�����2��Hqr�G��vR��<둦ɲ�u!s����U(ݣ����|�������L�nչ����K�FJ��K �bK�\�΋S$� -O�������ֽ�����U	U6�Hn+*v�<��p,����\�BqP�+?��|a(��Qg��MN���zP�i�柅HO���xчÏ�������
��/��yW�r�̷NOV�~=&Г�"i��$c�W�9�_�[��+��zP�D��O��%fZ�"�h�g��Z�.[�k�/���xq�M{��m���C������X�2db1�3���d�,���̲�BN	�Yb��43��ߥ� $�uc{�s,�����qP���a�Y�}��Mk�Q"�����~�~a�t�[��>�n�U�_�v�(� ی�@Ɛ���2��������Z@h�:y2��u��������ъ9p%�d�¼���(�Ϸ�m������u]�O_d��~�Eٟ�j73�!%r;��;ح8ɛXK�Eg��u��jP�`.�o��@�V@���e̓�_9y3T�(q����,L� �?y�-p^�l��,�D��rV��Vh�Kqa�J��VI��Gнvc�R�xN�6a����3򺞮�I��ۗ�Q������ӡEl�7R�Կ\>���¯p�-�?��MK�p�u���[�$�;�:���+%袛f����Ӣ\G����ԐYE���Uo���ac�&�/U.�lS�"?�W��:+�xa��D��2늛̥;frU��>j�(P�f4��7��>���Xq�N@�*p�˷���0�6&�����G�����9�=�����~�|4A��`����]ڦn��c�'&f����E��'6�����V�&��6�-gӰy.@}i)@�R���^�x�@��A�-�SE3�`��#�ˌV�r�qo�8�����L���]�+��DUE.\AMV��M���W�2X�ȼ�o@�:�H�O�M���S��ڢUr�r
fd��RQ����[)�2��ݯ�L���԰��Q'�x�F}�%,1�m=�����a/Y҄4V���=^�Dؔ��TQ�9���V�#R��Wی��	(ռ0��%)�E��������ނ$ ��o�ՒkM����5���6TA��I���>I�ף��h R��,p�c��)q
��nB�a��M�7��t��f�G,���ZE)z-��T�У�.��j�i��7/���r�Ac�jjy��.B��r���V�&���4��
is�M���U�\���i=A\ﱿ�X�]�����c�H����yTu�7�e�F)K�v
�l^�D\چsI�BcaR� Z��k�D[ę� ��N��G��-�,�Ґ���B��"�� �C5��)/b��щ�X��-Wn�	͌��'��:��@�i���D;:.���s$U�ګBk�u��%?�@8���}�'r�/X��v_M��!�%1I�U�q�?1}18Ф��-~�[���+�F�:�Ng1N�����l�I��5������&)jڠ]'`��	�n?��i�gt��H�����ַd�@�+*,;�\��n�[��ם�^�>���<LmNRUn�_�YX�Ւ�|Pɔm�F9�:�?mN=��@�03�o�1�}o|����>ߚ� �\�ֶ���������z	B 2A�i��KĂ�B�|��%o0�ӁF�!�,axv[���(�>!���<vl�af.�f,�BJ��G/"�	�$�k	T�{�}�E�5x��HV�s�%S5��ů�ý��V��5'���k�Ý14hO��p���TMR'���fJ�"u���W���'v =�Y�ن�)�p���\�̝��� �FRl8�7�c_i�h�4\亪�Mr�D�\\�0�	�I�giD�S��/��N�[r#�ա�d�X�bx����	芒3��`}��+_�
 �?���U�����xgdy/���pC
��}������>�/>�����a��N���)!�O%0�ʷ|��m�������߮-��5i���_f�!��-[�nc��/.#���q��"����aW"P)���Sr*�����'�]�5�>S��Y�f�;��s�;�)q=C���,��t��+�ň�ڲI����ݾ�]+W�6ph��	��z�g�[d�'�d�T�`��PV��lO
.��2^�*ޏ��x���W)^�Rm\.u�
\�,�ex&%5�&�")�Ȇ*[5q�'�W;Ă;��Xu��ȴ��2��E3E�8VB��A��p=���:z^dW+��Wo�?ZiA��,�Zwp���JOs#�H_I^�i~������o2�Z��'�K����d�	zA;vi��V�_��y�[ƙ�4�V�D���9��1i;!B� �-	:gn"Jر��\���8]��l��&���|��[��f2i P��>A)� [��G�hE�?�,(��+u���o�.�[CT��Y=|��4��5�e�zE�za@���;�9���xk�^�k�U�'6}��j$�]>d��:��0!��C�7�v��e�����c}~��.��d)_��;fYE^7�h���^���0�	]����)"���\�߱qz�'f�����x�X�+p$|3X��UL�i킐��,EO�R�ƌi{w�3�Yh�6�B\�4�d�+E��]4�x���غ�=��XCs�~j�F��n�չ�h���N��5^5��׌��ė���� ^xhd��o3<�h=w~�Q	�O�� ����gY\N�^���<�~�.��� ��Ho;
�qc*T��._f[Wc��B��sX�Lc�{FϪ&As� 6X�?Q]��+����Q5f�����@`��Y��!d�gp��ow�t���?`�L��/i=��4��0��O:�$�D_b��	�n�j��M,�7g.Î�M?��<m*4[p��_�\�lkD(�N�����dLo@Q��i'w��L�kO(�猊u�]y\� �ad�l�W�0���E<"���/�7�(3��4}~�g�˺SLҞ���E�a��B�Es�Iv��L:�5n����\9\��q��p^z�c�t�;��
�)��h�������3�2�!8f��\�6��6�ARͰ!��	4T��Dft�o��!J~b��|.-V	C#7��U,���x�?L�,o��1������z����4��������y5��E�v��:�� q���y5�ݘ�=�g�[���[�Z"Yh�ψN�"g�*��wR]y�wƊV�Y�M����ˉ�=�K{s\7;��zˇb�D?�ڼyWQC���Y�^�!*A�(.1F �V;���~��Me��0��Y�5����`Vd����Hdː�[��I��[M�G�H��="��^1c�p�\��ƍGu����������~�·�3t�����	4��9&I� �lu�T�'ӿ�[b!���c����w9�RM�	�v��(oP �T�W�n��/\.�꥽������m[�lj&L��2"�w��
���P���b��S6֤�ٮ�������\�m�{I��]b�dC���Z�+��5�xx�U/QSܽ�1秏7i.%��\{Fy��T��ЄFbȯ��$� >�<��&�EPfd,�{@t,lW_�y�ᮅ��8 ���{o��Q����O���Q�#�t@hJs,�KJ�����ϯv9��Y�c��z����u�es`����3[a�kBB��2v'�*Z��^hҀx:���۶�@��aO"gB|��cz�F9tq	�l�k�����9�����%E����
˜?t�N��7��U�>A�a�6��ߍ�z���KT�ҵN�>��ٹ�۳SJ ��3�p�\�.�S����w���U��~m*�X
�fbp)O>=��YUE�d�&P�{mU�����u��oAAX���&I_҃��iˢ������������D�FW�?y�)2Iˡ!l�&�k�深m��=��^�yw"7��I�+�[�<�æ&vp�G��ĵ_���^	�ᗹK����_Hc<n�� |C���R5�|�@s�@��.#%<`�Jh�Þ��?�uҷ��j,������y��6�	+r�7���!rk��0����%xof��hM�e[��0����;5��{�q�Vȭ�ݬ1@o���^�řs�|\}@Oi��V������&���(�����'�B�����%�!ٜ��<�:j�����3f�~ס��PtP�!�A*<�q��/ �iw2,/�� �_�4T�8�b�Z�s{k�.�\,r��
�9��}��W���CN�Q�k���{����!�&�'t�&ǡ?��w�\Ǡ����?�J'E>MK���A����${TMw�_F��	{ڪ+ ��Zh���AڴJ`֣�Gmo2ƸZ��WI�>�Y�$z�ޛ���ٵ��I���	 ��Z�+a�jS�Yp���EP�28Jģ��/��s��4�SՑ�	��^ӭ�> �JN�����>��@<>��$V�M'��=)k�����ǒj�T�Hk�؇cA�v1]Y&[5n�xc��-N s�m9�L��_3ST�7����N�����������N@��� /=��t�RD�o>�͕n[�Z�[q��lg/�gF Jh�����ӥ2G��c��>"_�0�W9w������l��B�c؁N.r���C�.���L����a����{�et�e�Β~��2I.��4�����e	����i~��	�W�Q�д�k���؅�;g�І�x�����Q��]�A]d������u���p�u�z'U�'�5q�r�ڬ��w�`�N�*��V[CNQ�&�̽�ap���}��ٶUYś�[B��e��8�T�F4�� g8�Z�O{�Ww�-������4{^�����ص�"��˯�����5V;�q^�A|�T�Tռ�V�+��t�#W��2�YF���EAo{����]7�-/eI5%��ۊlObY賤N�3z��]DD���TS�T~jP�+`���32;����.N���L`�N�U�|L@6��0�=�W��#����1��������&���_��ޟ��KTlq��?���e|f�'aK_Ӓr�����Y�%u��Jzr��E�)�P ��,�K�cMՏ I�/U�QS���h@F*�ap|E���b���t�"Yq?3�1xW�_<Ä��^�J[� K���v��}�De��b�(�z)3�q�T).�yX��c���6�7{�KmՁ�ԕ3�5�jHx��:�Nʳ?o�]d��ds̐�f�jKBcT(�P)/�Dj4�����>�|���%�������!��kܹѾ&6�	������m�J��o9s�4/�����!�v�0>q<��?�L�lV���|�n�������b0a�<.!�����F����˻{��w�HPȅ �:��u�m��vV9�0jE�Μ�P��̍��06ToA����^i1��r�>z���b�H2��S!�TP!Cҹ!��x,��Ʋ=ƫ�|���EiW�_�D|��R���c_��ʣ�>�>xا�����"6����l�_S %L;��K���H�Z���9�,�D@\�\���]'$,��(jJ,�Nl���G���H�G�;ژ�?�}6���o���R9)E�N���yx���-��G�ɂkV����zkХ~���r�0�U���Ӊyg����C�,��OÈN��<�~�������ʒ*��y��{Ԣ#7�ԠL�?���>J�v|,������]��83%����ȶC���<ml�s������#R3r���&��o>}N��i,��E�-z�Ȋ�>�~zj��SX(���xRG������A�,�]ā�Ä�k
D�՚��5s�r�ߏ�	�9�R��8�w�b"��wE #aS���+�A=aW!`���1+"8Dm	�[��B�kI��Uљ)�d�t��샀ѵ���<��6������v��i�#��g�\�r|(۴��z~yl�Z�h�R�6����^��GY��9SY�HV��_����CѾ�����_�j�=T�%(��[9�{>�)d���F,��`�n��E+`�o^�D�Qc�;Qt?���ۍD���K+e�Ԯ�ڮ�|o�)X�M���o9���ֻ�ͻ�9�)�.BEF��N:x[.s�E1��
�[ZGU�c�w!<A7����3���6ۊ�`K�f�'����Soӡ-��b�$�G]嗰�h��B*h�HL���%at�X�r	[|�u)��jHY;�tP�.�c&��:�E���V���q![9܍�n��&QN��dȹÒ7�G����ƞ[�n���t��#;�Ϥ[�`�S������k�}��d��۹SͶnn��� �4
":wZA3ޥ�6�����Ӥ�B} \Z(Da����eI�@'��ROe	#��o�
%�Q�H�y_�v��,��▭{�I�2/�ak�B��������w0�_�w,1����bҡx��@��ϙ4����8�$|�o�,����Zm�����:בB`�W����\���t�B�����H�po-��&����+�7A���"ү����2Ym"��^��	?����O\��J)��u��/�ptmi:=�2P��Ɛ9��uA�c�`aްs�7� ��1H��e���=}�\����x!��5K�sE."yF���Q�>�N��|�q��H#�$�g��>(�샿@��Oha�9��W�����ֵ�$q]Ie��v[V���.�!�����L�L��|鑮������,�E����Ą,,������?�4�}�j1Xh�iyď8J�:QC�,�>����3e�7л�.^C�7��a�r��U��һ��xn�D<Z���G.�n����?'�������n� ���oȨ��Ͼ2W�R~
720w$S1�7�fC����J�y@�����+��Y	�T��]�r�n-�8-��� )��P���Z��T�ӌ��`G�I�5Bב	Q/�>����Rѓ�~<���n�sOt��g�S�W��3�l�g�.h�S$D~����j��ܴ@��D���3�rZ���S�kRQ��Cq�%#z�����r�f1�Za}5�xq�*��c*3��CcB7�'����9|L#�a3����]��>��ɨ�t�5Whʑȷ��J6��p��@I�I���'��bY`q��L�tA��#]�7����4M����� z�襓�@�
�Rx�F6��3�@N�F��7,�Ni	���K�P��j���b�P��3~�]�8ݺ��L8X�;
��d�RC�ڎ��W1{<�R��N�~�?����M%�b�_�C?�y�d��,$+�(������L�2<�����ێTo"��6�<�����o�m�������k.��x�뉌��(Z,����i�9@�%-3i�g�.ۙ[@���(Q��S�v�� @Qf����/gc��� �|��Υx]���L9���	ћ�n�x�&�/}]�`�U�䤜�̬�c?>�$J<p��ؘV�04�ėQ� �[h� z��+w�5{{��R�\�Ħ�t������v�ޯ+A������}i���LC�8��j 0�����3]�Ro:vv�P~1_2ج�dV���d��e���z ��xj�I�4g������aXa_t)7�罅wqZQ��t#:w'Ɣ�m�o�)�(D��\���t2�$5�<t�ǝiWk��ZR$�(}>P"�U���ӣ�3ԂѷvW�@�e ����G��l�ߋ�}��x�3�x#2��H���	�+�uR���{��*4_��1�=�)� �Pғ�\��%�7��<�"�y��
��m�Sf�_ґ������z�%�P ����՟/�1]� ��Q��t�1j ���4�V�+������ �r�}�7�.�'���D�w<�6M��<i�x�zHmͨ�U�w�h���D�=a��Vx�'L�o&1�t<u��݂�t豓��ky�qG�C�K�p��D�n���d��g�`��� �sONӐ�RP�J^�j���X�J�g�4h��KaC��>[K�Wa'�j�2�%>F���8�Y�+F@/��=B���ܭ`K���{��� �쾓F�Ŕǹ�M��'e��b�.ؼ �#�X�� 6�X����]�&��F�{��Ѓ��=;�^�2Q����0Hcȁ�#'){�Q��d�:
����9W��O��	�)L�4d%Y@�:>�%IۢzaW���`,T��E]�Ȕ��5w�/����a������
u�f��"�.:#ѥ\���4��i��zg����D�e0U���]k���
�'�˟���m	 Yb�k�����(w4W���*Ӓ<o�r�!]5N�b����8���i��#�yPw�F1v���wZ�k��Ec�2� �q8�
��
~2��&�B�`�|A1��3,�Xg�0�#VZ<MJŲȥ��	�OA�n��_]�P�����������5�P:e`!� S��I��^�ӆUW�9?�kEY/穑5[&�bAhB�( ��\f��i}H۳���(N�����/�?�~-�d�}�F��"<�Κ��2�֗��8E�'�C.ҕA�9�4ĕ�f)��B�<�F��}0�����Cs�@	e��_{3|��݄�l��\����}sL|��z�~䇞�;,'i�)b���d	�OP�KY�*@���!����Ƣ���5�O~m�Kǥ��謮�^%��t��AۄCZ�g���GwCn}��4�'�B�d�^[��,{/FnUd�Ꭼ|X+XЃ��N��m�w�V?�����p�>������^���G`{L�]
�[nC\������vkګK٪b����?㫶��*�ݡ�.J`��o����h���t�����SR�-�&$L��T�#��	����*_no�-7;udK�����O"	�=M��:L��7y"�R¿�`YoDY�-p�[�1uvw��A|��B�PTS`�^��ǡ�S��k��5;�(�L�^d�H�y��p���q�Mpj;�*�ڦl���;��tu��Ųm�Cm� �f���/���/2/��m�G]��Cp�d;�عF*�5�,X���������VkE�CE���гPQ�gԄ0��&v ���TV�����w��h�����F�O��; w,�B^Cv��Њ���]e��X��_����X��'�Ҭ��Q�[�~�����=��j4���n��ՠ�_�A$V�p��t���`j����)Ǣ�[�W���Α*_,��t�,6!��1b-����<#��I��5��
����a-��݄:�X��&a�K֠�� :�T�1X2lJ6�}���}�" \����q�1��� �MB5�4 �d��|����������s�9�>ac��.�A���Lհ*�6�b���[�+FkW	y|�8�e����S����.2#�7��u��֮O�[�YdZE/���NAd`+�rl���@�F�傫�
.�Uu­�rI��	���c{hl�E(z`�B�$&����T-��bT%�4��@̸e�&|���F�!�F~��G���R2|��UhE�=Kq����0�2_��vJD+�i�Լ���因u���O�C�q�"@�ĵg�܁��Ӊ��,�
KF�V�d����-�P�Q�o5ݯD���h_���$��ݖp�/x����Z�eS�R�e[��^��/@�
0͕�`�u�Ժ��J�@pT���e�0g��wځ�sj����~+I>���p��h�}'k��z�z��Z)��팭��:T��e�d>ɟJv�g��G�08�}A�$NX��C�!�H�ٯ()�
{���ԁ�����fB�6F`|]r�҉�%�~�\�s��*�X�_���T�C����.y1aIʏks! �X�6s�W��PKQ��Dg�����i��>E�<*}���:��"|�	�
�G�V�I � �Z�7{���� 9=�,�t;랦��L���ˮ;�Z��<�R\$�d�	�'a��Y;��p�W�3�}T�Ǭ�m��Bl,���<$+����`U��Cqߌ^��E����ͶT����/a�˱���k��6;ᔋ;g�L 3A��T챶���n�'s%�ƒ()�7�`��@���iJ��8�PD��>J����!�0;~y/ !�<��m�B]�&�i��l�����.Z�)��M�1���t>�ձ��7Є�*���g0�����϶�X�{�zd`Ynx�m��IקY���)�Ic��z�9�sW[�
`u��lֹ�:��q1��>J�=��������3�5�>��fb�&���T�,(��%ޑZ�Ҽ�	]�,(v*���U�W���p��9eߞL��[>�XJ�UQa�S[A�{_�2���(F���H��,�-�'o�o�t� �����d�C6><A@I�(�DD�Qc��Uw>g�W��|�˽���N�pp��SopP���G���n�9P�VB�˛"1��1�Q1�wJ%�g��8~S�`��5n�Ո�.X�lfX�j3�[]/����"똦�o��0��}�S�}��hi�<��Z=���{��[ڛq�s�l{W�Q�<eZ$f9�2�.ˣ���	�u���j>�����5�v�5@�a����D+���	>Tq�%�qC�}��ju��l������`
�#1�BJ�Uc�U����;����x�Ȝze�����n�9$T4c7�9��y}�<sx;�@j_KZ�P�}�O�EI �'�&����>��vf�s��6��F��3�J���C�N�����\�O���z0���%�������Պ^���O}�``��nT@���^���e@O�3ܧ��`��]����7���:Xq+����s�v�?�%�"2Y��g�_��gͦ�:�EK=������l?/cl"c��uw�_��1B`��]#[q�?�"��	�m��j��:���r��c*2@�C�p�7W�X��tpK���T�f��K���2/�xD��X�Bsa�������qq	J�J���=1�Rb�<XD4�I��n�cޘ��:��L{N^�"JHŇ�ձ���zͦ�>=��&"/ցu;�����άtB�O�>j��$�U������f���.ԕ#���ʻ�ͤ+���uZƼ����Sr(��"}�R2�?t0�چ��ՙ��J�9B��33Q�#<F:�~��-��Ҏ8>���Z|��6�����n�;6�Ph̅F�-r��k��?yZ�H��	�=�f�Jq
�G����Fi}f��g+hT�>��sb.����r����Ŋѵܻ��>h���ln����c��x�܄��R2�=	٫ʇjY;��؂5p�
 ��<�[K)U�9�]hG\B�^�$Xx����ꃎ�m6"H�).����O�� %��Yn���za���/;7䤨�P�瓓�y�a�5������ޥ+�{úQY��8uk���a�7#ډ'���p���q���vu?d�@5���̪TO�Q��c�}����f;�nv���v9�_�Pqa֐����H��r(�]��͏�{� �D��q�G�# 8�N�l�@!�`fѲͣ� I����X_��T-�G�r�`����d(�8��:�ؘ�М*���]� �
�v*�t�Z��w���\YQnj� ��U"��Hz�[�9P�DӁ�~q��=	����׻�kN;F`F�'&/wP]�
�>��S����<=�H���r�]G�'d�$��)�A�l+˂D�����I���w4��U.�D1�'YTJd"�=ms)�
x��E�8�Ȯ�1�Dm�c�^i�k~'��wD.��5m�\���~#x�C?j���+߾�8�����_[9�r�bZa.�����q�&�|/=�Ԫ�e�9��d%�F	����-�CM���Z ���\U��ud������;`�4��Nj��"����09/��qJ�9;{Ò��ޅ�����,���-�����7����f'�CΫ�W�K����u�˟]�IT�1-v'�DHqe�0�(Ht�D/�B�S�ͶN.�+� :��P	꽃���@�Hf;#I�^���z�(w�n ��!��^���E�P0���P���N׳,�_5o�'�%4=�Ve �� ԏ�c�H�RNYCK�tqS�;����Wi!>�8�>KT�/��5�`(P��vl5T2VT���t!���T��0^C�X$g@gv�.�r^q�>R6J9��x����6m���2W5eC�hg���>��Yν�оs ��ɀ�U�S�������DNS!$��"X�G��<M��X~@~"�t���ד#_�-���v �F"�}�)m�N*��}��j�;y*?v�fF��d�h�����o��Cb� �0�
�aLR�5�`�IQ�jG�(���Hߓ>��NE��^�ڥ?H4�#ֹ�R8��j̇�-4망|�:P��gV��X�Pfs=�H�t]RJ=!'�\&s��F$W�N�ĔMu]�5oO��L�:�	��h��P�*v����:��N�\�[8����A.�wq̻�Z*��I�"l���~�f�^��<��mU�W0Q��	�	�����(d���8 �$X[�~�k���ջ�9����³bh���Gd����0]ӊT��_�%���|� \���((U�U�v�(:B��0<�xz ��d"[>���f"9m*=5����*�,�;П��M��v��rAOϸ�R>5���-^����z�L���ce�,H�&H&?�r�B�rX����u-T��Z �����n�-�Q}/�;e�ב-�ݖ~R�Pu�ԔE�
�J6ܡ!���n&�W�D���