��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U��S
��Q�$�#�̓�tk`����!/����Gʁ��C�����Ez�h�v��a0@����Ù+�*�a�t��w�E�t'�����\��i��V�
H��(�����SǊ�},�gd~�Z��VXR3!q��3s5*P��A�2H�8d�]����k��S��=bт=�ҭ��&�V���)�Eܛ7���ؕ.8��2 Yի[��;pts�S��a��RgO"$0���+E���.��٢*�R֝�8�E��s�,�¼���=��Y�Ks龇V�ؽɢs]3�/O/��������s�,?n��$x�,*��=v�IjF�4�z�P���`����`,��w$� �M642B:H��q��b�F�8<���MQ.5�5M~D���� UO�yt{ӲL�/��
V����\HeG��m�=�C�8"��G�����Zh������ӣ�7��>�mf��z,���SH��/�q��kS�_���t�)c�RE;M,�������������o���Y����'�P?����O�%��%B��./Y�$%H�i{9uS��(,��g�*\r+	'��uQG�K�җ�����D���7w�\�LY$�Aݨ�ͺ5d�a{���e�t�5�f�K6K�`PE���e�G�O�������CS]�ϥh�I��A dDR��|)&��Ui�L!?�.TD+{�/"����V!bu�R3����=g� :f3c�7IA�>|����K�����eMX2eV�l�Q��j�UE}T	 ���w"��������N��:^�_۟����z��&��vʞU�fC7�h���bJ��&X��:|�o m̷����E;��L�6.˗Ǿpɥ�Rg'U��|��5�q��%Z����
P��Y�u��4p8��.}a��c~s��a�k\��<��!�d7!�U8�R>"�������j�w�MQ�Iq�O��R�I�e�}�Ug���N�k%�?���ݕ1L
��zS�+x��gAl[N=t�g��9���yu�qK��<�Iߌ�}9�c���XsWM�P��c4H=)2
 �p/w�y�P���^�BG������r]���r��簥�V.��Lv��Ϙ���x�ƕ�2�kg����o�Rڔ��k&өKnO��(tl!p���O���|���l�fإb�m�	hĔO���Hj��ġ�'��[ؤm�*��,h� ���۷N��S+���H�=�SJ�x	Og��5�BD^��}|$:�6M��;�����{�7�Lqʘ��x�k�md�X�$D�K����+�k�%��@�|j���2�]eey���
v)Q��-f�y�<	k98�a\"�[�aX�P�V�.\j7�c�#Y�m�-��z�O=+��8Ħ�e��o�bo�G��W�r?4� ����{A͹�v�n��M���%�^i �L6u�1���!0�&��,W��f�:��n�X��ɘ[�MD��:���$�{Z+'�tVw���CC�K��Ґ9��R��cS�W����E�EqF���MG/ܸ����=����	dS�������E��r��r��Z��%(j�LJ�f���Z�s���A0�Lp
��ݛ
x�
��s�YLf���s!��Z��f.Bw*��Q.w)�#-��W	>*n�಻��ʞz�����Q1��u\���9}�*.��S�m�ԝ�'�	C�*��ȾَBG�aB��p��#ѕ��W�ގ6r}�I��o_������<*���{Tb��rn��u��0�cW)ѕ�Ï��_'��V�xB:��v���-Y����\�+N�;W�c�P�ӆ�w�8�!�r�C�U����r�����i�0�i�o,�k��	Mq�'�x�S�i�1�,�a@3!s���\j{�`#EX���m3�C9�ٛ�����8��~w�3�@fZ6�b<��m6��׹�,j@�F��婭�'���`^�w[V���r,�%���t;(�k�k
2�Bg��Q:��m=Y+��R[$��뎰|:�c�tW��G1;���p���_ѻkm����n�U��? m��}Z��O
P������;�!LNl���Ij�Y� �Nq��!b�)���]�p`��T��m\a��P��P�6�~l��H<N\�,�h�3��mJ�w_�ׁx����؉���<�j����bZٝ��=&��:Å�xD�x@������nܐ�'3��z%ҙ҂�7� ��z5��=�Sc���S1��&������iNj��t�l�Y#H����b}��Z���$|φ����"4�e�Ye��#�!�^����̕�o��7�g�� ��{K�j� rՒmn�eyjI؜g��l����4�ajO�_�DXb����� =�k��A}���Æ1���5@�J=B�M:(J_�����;x�4l��J4��o�q^ ��=�,`��W:c��q���[�9�N~��'ژ�_l��.��/�A����|xPh�.(d�]�(�ݞ+͐����u��t��ٴ>jr���ұ��G�1�\kvȎ��
Ů9��V�Ckۺ�W��!��ɮ�*�9 �?����S�04���ӣ7j'�4�U6��W�X;��Q��c|�{Ϡ)�����5<��D��5	}�2���VBf�?���ԥ��ƨ�Á�=t����┓��@�l��_B����t�v)�N�.-���X�����48�*�i�A�7�iX���2\Q�~�L�v�Zح�^�.z��b-xN�'���	$��"��l�Y�{����JȺD]2^�ٌu����%vh �Eu�7c�"�2�MOB����#��.狭r�`��	e��?oib��9)��i�~�����j���F���	�-�7�3 O9PseϤע�c���f��s���dq�$c6~<�i ��ד�(�܀M�VǄ�X�Vc�fp��x�%��W�]6��?�>��N-YM!*���L��4�J)U���[�"qR��Q����ױx����=x8X;�ni�wp�<�� >p�>\�H���Lv��GJM�l@�##!Q՗�ڳ
آ1[%2�>���׉�[ko{7T�D�(��s�</��-��јs�R��^j�����:�.�x��,���"N��Ka��T9~0��H��U�f<}b��A���ч����H.��#���;������oS���+���o��K4PԬ��d�<���\[�s�\�����N�����e�b�$B��(�Ub�n=�t3��|-�
��~�W�ԌBB����.�+n?���g�-��OC�@�փ��i4ǎݬ\z"���Ҳr��F�Q�K�H��p�Y��bM��-�[��0��N�)���P��5��}xg�la⼺r��Q��K���F�[�g�t^�z>�L"��v��a�	�R@� �Z���옖���T]l�0E�%���Zy�Z��D�3��]�����t^l���qI �"��+�=,Ck�*��î�V��l�S��MW��s@�ݔ>��r|ܚy�\-N
k�2-Ãğ�s��ٶ�/�+�o���l�XF?�Ue�?G� ;�t�z�o����TM������V�t��{���1h���N��)�faѺ����8�c�0��k�eC�i���H�����Q}^��r�W����0��2�,��}t���]��j������f��#�P��"��W�5b_��E�
+K�+:��e�t��eU���^�+��~�%~@�̔!;z���|��\��XC�j}�Wi�'�� ��/"R��x?��멯��nt^�3�*=�w��2)�Q�{kof�lgF}�W
"��A���n%�*�������Q�%%�k5"坞��+�6�(VI�OO�ϖ@|��q��-����U��Ѱ=�,���t��M �� ��z2����{�#��ڶo�s.��;�|a��R�˷���m�m+`a��6�v'�R�䵣����s�rsMZ������ N!|����$��%�m �sq9��c�u�� ��{[���l�y�-���'��*h�<�0��z�ܣ�7&�Fn?�{�	o��I���naZ�:���79�3 �G =�}���`�C8
N�´��$��9��Q��au���\i�:!���Y�n�k�d�܆wލ���U�j�ճ�F9��=�'��z�z�3%�ɣ�G�a�hnMs\���+�W�0�d"�9B��*Ds�ے�Zt���p 8�_�M���'c���g�]'�.@��)�b:p��xR ��!FC_�]�F��DDYx�Y��RY���	���B�M�`2S�4u���EQD`���ֶ0`_���sm��tmW�{R\��*L�O%Bj�[�����AQ	Ab�B )��l�OǬz�������}�5+�V�
�7ߣ
�������W�B#`�-(�$��ޓ
���WF�,��������V-�i&Z�nI�T|G%��C��l;��e�9��B6z!À���� mGT�Xvy���i��9�y�GQ�B���$��A��I��]��Vne.�/��x�V�tH�H`C�q>��0�3Zhwv�kz�HP�k�{��x���J&Fg�vd���7ѐ��r�,TǛ���O�y���(!\f�=�Gi�qLW�R�� �c��\����|8�y�d)p���7!�������K�ի:j�aL�-~���x��H��bX�����k-�e�{��N"�)�8�����J������._~�`���"�ĺr�aX�e'6G :�u�邶gm��y`\��V�Mמ���k����Q���6���vVf�D�b®�F�;%%m�x�E��ZǛ$>`��	�
L(Uvj>+^1�4�K9��)�+�ޞ���o{[J�����W�5罈 6���&���{���Uz�}�������\S��{���䶞4D';���!��5��fTj�n��v�	\u�)*Gs���Z����O�����Cy��n�d+�o�O:1�@@��}�$}*ÝX^�q ���<(A�#�MCR0D���B!�eŞ;"'�&����(р���?B�>��3�·Ow������x��9���By��t�(��`�q�f��V�Bw��2�tc��Ar�=׆%��T�:���֝��g;w~id��=��h�(�F�vC"Nҵi�'�w���5����R��<'(|O�T��J����UYo�����[D�kmr����9�
D�Yf����Z&I�w�}x��'}�'�t�­
�r&a��vs�����]�T��1���C(ms(iZ��;��7YO�x�|V�f~8��ZM����J���S|��~}�U:�mGUIJ6)$��1�Dl �Ф�"7�,���/�T`q���QOc�n�-	b/2]�Wn��]y��i�����,�KEr��-l���'�m�=�絴� e)Z"�� �>��H�G�n0gr���������/�I�T��[*�fL۩������� �^q����B�G9,�.���Z���[��7�!��I�vI5�e�N1W��1�X���>D��˽h1xAz�q�=��L��"���Uz-{Y�_g�xR0V&Ją��u-���x�)hzGڷ� &�Vj;����ãdC�j$���|���J}ԧjO���nRoDe�6[P�g9׀=�<ꄥ��<����%���TB ���	���������.?�Ό�V���)>��:w�,�x��{�����Qe%��B�ͷ`-2ˍ�FY"���Zc��������%{.j��j�ͦCN��ݔ{Ȼ�03 Q�����~�b�~n~(O�4C�M
C�^B�90`��ګ�5���#�ff?�CުF�A,��D01}�QZnc��jkhsd�q�ٯ�!	?դ��G��z�����Y�� �5�⁜�o`��͵=�-��S��JG��f�~֬�p�L��0�Y)�kZڜD�=8͓��i	�F��3��>sDQm��c[�,���w�Q<zl�g0o ��;����x���YߺP�Vk
���!b�� n`g˳�O��m#�ٸ(viE��qr��D��V�o�1g�E�p~���@�'wfJX���W ���������n�M�Æ� k�׭C�4�VT�C�ΊQ� �^�흱��KWJ���}��1�7�=4>��%�%1�m�Ys�q�ad`��ˤ:�̮B?OP�4f��'X�	�C�lz1�rud���̒p�-/���[�傞�f(�F�Kf'���Xi{�4<3��.��?�i'L��L��U1[��Nכ��!�nA��S'%Ʌ&m�Vz襴��[��Y�����0�)�ʬ�OIO�N����ڇ�c�Bg�~بb!޻H�=U�C��O��CZIC� Q}�$�!W%DsHH �d���1���Q�5."2@�)�o�h������K'�ָÿ���(����2�F8E�;s0�w3���EF�L�*�ϚN��|�� K�ޙ������M���H/��;�f����Z�����*.���v�Y;e��:���*���޳��)���ZҞy���<9�.��˭��������Wڋ��Ws��6�G|�Kx*U9�,��R������ mz�9�����k��;v��0`o���x����j��|���'(��#�
�$ǣ��V���s⮝Ͳ�����_#��M��*e}���$��e� ����Uy>yu�9vM����{��C�MAԨ8�i>u��1ϕ�Fm�\ڻ!Z�C��pήa�^�Y!����lʲ_>��^�,V� U��YO�q��K=e���-��� ����Br�4�o^]
�8a&t�m�.w'�"ڇ����X��R£4���$�=��z J�(�J�z�������Ճ{�B��Ao2vϾ�"�H���<��N�!"C>*�j`�3n��'rw@���HC1`-=V���Q!�4�4����)��gS�{�SD�U��yH�)�y�$��^:}s�}H;ȉf���V/RP6�j(�Z ������mDA��l�,6��yYUE_("_�䔃w��TP3�	�X�b��W��E Hٰ��;��?}�@�/����p{��Bi�w7�Է�ݲ�S���2�T=�5��#ݱ<��v�ttsܲUz��	Gͱ�6���0�J�M�&[IB�`<NG�K��?�	z-���hƘ���q0��^lш#��Ǜy_�G"����uw�f�eb5#E���9�6[�n�:�hlR�<�A�i�_U���d��~�6�B9�SS��,�,��,D�8���$�����T�v��17/�jo���;'u��k,�j�=e5j�	N8)$#��V�?���O���Z��f�(�h��N�g;�W��l��s-_g�������P�$��ͮ�_+�f�����
Ё�>�*��v@z����8z�vfpa!�Ǽ+6T;s��D�_��@�K�0�t��6�,e��~FRS����|���c���o��,-�qg�u�����7��u�C&�E����&��߬K8��s�١6[Q%�g��r��s{vCN�h��;8x�!Ii����)lrl0�H�f�\*k��W�3�)�o�� ���� ��(��Ep��vx�0��C�[��/
YZ\g�V8%||.=3�����k#Vʘ�ǅp�xq��s�[�f}�t���JJ��K�;���M���� �5{��(kt�3��������1�0�,�m�/q
�G-<���W+P����$a5-�o޿�kpd�4ﱛ�
�6!�C�V��Q�wj�Ih���r��IaZ�OcQ��j��;�r���D%�_��.cj�� U.v��O+$��^sB�*�Ȥqg�|���<���w��)o�㜹[��^-��:d�;�<Iԩ�ɋ��Q��&����2^���q�35�4�G��j=o�Dc��Ocr^�V�%)��$�D�#��Е-���`�SM�|~U�Dw%B,�ﭜ'�	��Z2��{�%iN�'c�6�n�\�C���6��X"�=y8;�,K��)=_�l7�J�p��5�bm`�H���d:���be(�P��e�4s�GAQm)���A�Z�
���2�K�FKǊ�e�p���#E��ܞ�= ՉR��x�t���:4���,�d��g�E��}�����4�����d��W�U0�?��7M0���)�l�C�����f0vSy�N]}�bk�t
vb \#�����d�Y��z��5����j[����D�������ƞ)��ߙ�Ý�o������6\�\߲����4F�DůK����(;��ŗ_eL*���Y��k����ʙ ��%K�l�Fސ�qS�޸�>.�O)���s�9�������du%�*��>��k��Q�)�p��T���V��˨�����İ2��=�$\�#)m�h��vT�"��yÁ�B��ٰU�����	�(B���0-xԒ۵�)�%}�o`,r��xv46b҅7�&d���h�,�)#%�xq�{�~9��-�H3����b�"ߥ��-v�bE�(k�v����ohdvwuQ�D�$�K���λ�/�?�����,�aY/V�0s[P��N�_�*a���X���̬Ȭ����.��sK��fy�S�������E�M��HSs���5`������6�zc�Kic�ۖ�������P9Wg�=�CKu��^_���.�� &����[�u�_M��j�X��K�Ha�9�aX�T��_��h��n��u�u
�SDhǟ�^�6��R�~N�Sʿ�����6��]���Ԝ����ǭ^_��hZ�m
aM��Jj��'�l���vЍ���%��xs�������r+~���#�b��~�H$���	��OV`]wxcJ�a{$�դ��MF��=׃�� F
� �����S&�T�Q	E}�
�_��b����m���F.�����n���� ��
��2�I8ON���AM�3����%�R����-�\?ǀ~ �I9����,U�_dZ��eU���З�g:殎y�i���)��Q���v'�t�%���먏bӥ���[V�>�[d���"�u�Q�hh����bm�yAj�4�yBE��ϖ6��G0�ₛQ��`��9��++�#"I��Wέ�U���
�^d� 2ޜIv ���z��/'8FhQ#��x�����M@Z����59��dWu3���NE`0-r5�FK8�Y`�Ȼ,w�
��+�h�����I���4��6��O��¯2	z� ͨ~�������~ґ}���\�D��G�S`�S�=�����[<�������S��1�Вp��O|��#�EUp�}.	�؂���U?��@n*��$�H8�fR��=@r6����༹GMA�<�6�vlo�:8tV�t��Ǧ�MmӖ,,�ل���Ss���Ӹχʴ�<A��_�j�j�°������ku"B��Ƣ�|;���Ԣ��ެ�	�����Qd��7���?�+s0K�J�5ٸ��o�����n"�mU�������)0<�Q�Ù'?��Wk���b�}��
�"��[)p/�DX�W^na������������|��^�7����ʦ�_�jq*�w~ޝ��D-�48L��"���ufQ����G����B��$� �i�Y�����I�0W����Y���L�Кg���y�/����t��I��� �����j���D���GdY��_Jl�g��l�`�J��(�P�j��ͰJ���e@T=�M*�m�&����w&�Z���Q�	�o|��P�=:MS;d�|����N��-�)���6���
�lY��I���.UG���u��h��Ua]h���$����I�E��ݖ��q)~�pz�'aDBtI��\1����K�\MܟR7�M�2��`GF,����g�0��:M��Xo�2������j<X�W��d��V�"����Z���f��tN�F�oC�������*�	��D W���T��~���!��9 MF��%�X�G���m)o�4\˪V;�g��(��'	J�7b�Ctnh�,����L#Qs�؋�o��A�qQ�����P]�Urg�_�D1����%OA��T
F�$�Y͌��ɐ�-���X,�ӷH =��ٓ��L��M@�1Č=���'�����-��\Ӈ�
�����}�5Q|���ȷeLS{_!q?A�[�����L	�B~U:���Vf��۔c��R���N�/@'����4[2lE���f��2�oZV�$^!��T:�I�^�ƠAvjmfk|q�cFUK�'�X�<F�t���R�f�6�6O(�P�٤E_�~���_#�ߤ��w
$K㶥��� �@�K$kT�5pG���gSj�;<��?G"ް�����4�R���˰���2%��v�2��0��?#!��K�P
>���h[��Z���1�<��uđ9E�lHo��0�I�|:���U'�&k�L5D����-�yN�BQ��@��X
�]�g�v޹d���Ƽ>ߤQbN�r�-~g�p�՜���h�LFuÂ'�B{x_�Cy߳�Wr�/K�/�£���o3�[�ϥ�W�1���;���{������d��U�zˢ%4۷��s��{'fp��&_�of�i�B�z�4on�^�-R�����������ru�Ҥ�Q`iwQ�󣻂9c�p�_�_<�5�5����]E!!:Ҹy�Wi�A�WH�B��<�H��#�����nє���h�d�"���7��5�<�n��àŭ���{vY/ҕw�g�Ӣ��y~�tuԼ�T��p�������=�q�Լ�	���0R���x���ΟN�AO��������`֟>������eFt�\�@|��޼�8�o� jkSF����ǋ/j���!/�q�>�`�,b��z�閲#(��f� �R�<�<����9����s��oʪ0H݈�EM�w|��?aEn����plB�*���jo��9�0A�W���.�߀[q��Y�#����vF�`�~�Hy��A19�����}��[�|��s<a_�h�2,����M��Oǩ�#�����V�!�(BI�B�٭��$�V�B<\�-�����]��v��rHK&{؊۶4��<��`1
4%V��_䕗�K��-�����#���h[*`�v]�2��'Af/3~�FJ2�K?�"�l$�}ca��D�*|��Rω<�I�2E$�/�)��lؔ
�p�(�Ve�B����h�ÃA}T�w{Y���Ǿ}z} 'J.�k���0��S�1A�u�,i��G��TP��PE3��t��g�w�zF�*_,��Ol"�T]H�	ɪ�FH��a�D(
O��q��/)ۧƜ�gמ+u/��. ơ��v͖�Zڹ����<�hQi���A��DF�QR��:��%�D�3L<��"���M6}���\*��o	�Lu���_�3)���)�C��IO����g3r{����� �|�Ȩ*���䎤�Y�d�	"������Q�=��Oۙ�m�ԋ(�n_��Mխz�s����<u1)��Q�ێ�D����E��X��]��7(��"��J��c�y����b��j{3l��<Ŵ�xyBh1�ђ\%����V��j[�KBN=Y��j���Q���S�%_�5�j��yz�t&�J����1�X
6��+���R�P9����.���ڇ~G6���e������ͺ��f�oT��`���	�L���-ڎ����i�p>�0'%zJ�Z�^��:ـ.�?}�]Őa�����ɮ�e�?h�|Bi��aAFD����Z��a��h:(��puq�@� ^,�;d��_y6��Wt��Lԝi���8����A�P���!��b8Zq�;>�#���V{�0�ki!����~�K�m'0�:q���Fޙi�dͩ\��o�#�N[	?���m^9:��1�-n]�'��P^����k&ѓ)���K���n����h�n?���/����~3� �ߔcF��v9��T�fq��L�y�6��lI�� �?�hzg��,8�u"�~�]�&��	��(���OH���	��6Z��,
�"�؜�n�U����t(PG׷P�o��E=
�r�y�״���yI���T��: ��q�C}eQ�J;��8,���y�V%�ZVF &�3�Q�)%i��goT'��`�5�"��Q>�'xZD�*,6���Os��f������#Q�_.z��{��Dd��ז�u�j�Fr�����Q&&3�����(-�	���8j	_�R*�����ΰ'�;un��/<��|;���/��u�'awU;G��n9֗�Z��fL:-�<�4z�K1�����Z�o�9	*.���������^~����b���LJ#��C�>�p�8�>i�<�1�����gU������ ��}癔�� �s�}e$�96@�,�+g;؍SQ�w#d���n�]U���°/�}���:����Wߒ����h����ӻ���_n��ŉ5s�xN@?4�{����|�<�?)9-����6���Xb�P���j�ma���m�^t~���a���܍�`�ӑ0�N�j�L��Jy!�r�%����`��_fI���awyw,Ap)r�s�:a���(��ʑi�WÈ"RF�h� �Kޭ7�'�G��� X�2�� ��:L�R{Y���i����؍�)G(/�?���v���.Ed�a�g�}��:�_�sY�Ђ�V�1��i'qWmf{oO2��ق.	���0�P����܌h_�9W��Z����.N�{�0�� ѭЊ �m���+�nCQ��P�*���x��Rj/�<\�� Ƴ�U�df�tw��c �r�G� ����ʔ�b^�o�*w%�����(�ѥZ&���xy
�([��3���p��쾉%�^@�-)s�=����0�tZ�;Oͧ6t%h@0�����e�hqG��"�ge���u�n�E!p7��qȾ� �x/���*�ޫ!3k�����p�j�N���ڭ��)Е��]�)�U�(�_x��Lk��U@�s�4�:�1v�;u��������3��:�J3dְ�aM��,<�M��g�I�a����{~_o�9��l�~����h��U  ̸W`F��o����3���Nǥ�M�?�-J5PjA�<��L:�t����x�M�Ҥk�s'��ttB7$��TVS�z�D>8�����*5���4]#f�}��d���x�8�<�am b�泘�'�8�����T 	l�A����u.���en�1����6b�����v���&���rf��!���9����,��	8è҄��>����/�,�B��,aIO��Ζ��E���@�r�١������և�oc��������/����soQO蔵�����������k����-����/��I�*�ArdE�I.G&w��1�E���	�?5N^z6WK������ڛlj��v�t�n`6(������)�5.%�ڀz5�QXU��ehd�������T(�M��RTro@��ŭ��HU��BZ�T��ʶ�X갎�c��?u�M���mH�q�o��83g^�{��N݉�*�B5}7�;�Sڪ�ˮ�)>��%�i@�o?���j��Z���2z�W\2�@����-gQ�z9u�&�#K/V���_�!���?�?�=��}����y1H�]�7��?L#'�	A���5J�d����p_[鍞�������+�Py(��S�]j�?�B�"��V����U�i3Ĉ:_K���W��}���U����S��9���j/��&�B2؝����0B��Eġ#o �{f.�I�ޅ�Κ�k��+Q;Ι���jk�0��t�[ܤ��i�
I�ps��}�)����Ϯ	�4T��<PadOo��"�*�V�F��:0�Tx|�K���x��r�W� ��14��B������h�;
G_�j��Q��nK���y��ZW��f�jf�e��x[CR��c��J]9fDl9��W�X3��\�+�ā[�S.W�#Z1ݞ����o<2bN"5> �M�V�J�����H�x΂�E�����>�]왒��cX5�2��n�BZ��ѐ����U���o8!��%�tfY�a�� ��`��]G�)4�h4	w`{�܁��e��9���^Y��ɥ#�LӱYS�M�Ʊ������S|*6�QYp��/�.n�Rx�T)��K����1z���B�C6�|� �����B��w
H}aЄ?u.U��qi�i@��oSf��o֠�w�d�զ���dNd5�
C�;0��+��01�Q:�U��h�Yc�Il~v���U�
�T91j� B��Z&"��џ%ʼ��h�����j��&���$c��Sd_�3��J�X��~ԅ��Sh�1-��E�	�﹖dL9���sK���q�żH=�N�D`�	�x s�AE��5�!F2n�Ӂo�.�\�yt1�&�&��
���ܭ��`}C-����H�\�n���*��`/����M�����VXv1�>�w�&Y\�� :�a!BL($Rgg�\�O�Mu� �&|�jNA7�΃U��)7�VE�P��-ҔF���>6:��s$��1
HIkyQ8�6��;?$�@���3|� �'���bgꩻ*Vv�lr��m=	P!�����2��*fU���a��75���JlJ� ��>�������k'���N���{y��&�N�����f{;p{5y-��������*�-¢sC*��A��~��ޙ��O��qɼa��X��Ŏ���^P=�S�j1���/����p$��e�e�1:�����KM�(���M��N+�E�����
>,:ݞsKg٠,(;����Ig�zDS�L~��-�������! �kdf�� gX�i�ii����r��@f��� �A�,�W:5�����z&5�֋�,��ۺ����x�6����dբ��_�M��8�e�*O�$�����Aw��W�)%��^s�I��M3J!���S�Z��c�4K��c!�K�n5H��a��)l�	_����}i&<����5䀕�T�S������)�څ ��رs!�@Ǧ����"��w��e:���%�u�6?#��:�u9v_�0
�碞����������hzêr�h���W4���JS%\�!�y!8����]���Z;7c�����՜N����q�:�+.@�C^`Ej7\ޞ+J?�{�@e$���:(�0��w�a�$�^A
���Y�ǅ�M�������3F�ia-�e�ʲ���O���u�#�J���c�xۇ��,#�,�3X�_\ea���[��1��r[$h���`GYm�b︱�I6o��`��t�S�8͠�ρ�᳗�G<�4h_,���02YL�6�z��j��U|fOb��6�G��Cx�[3�Z��ٲdM�����n`�0�$����0D}�A�S�W~ ���eo��qB��>�A��F�R��HѮ�fα�?5׍!��������[��3�}�)�i�T8�,�bT)����1�����}:7`<��x��@=��2��4"�8�7x����'����f<�hg���u|���4��D���[.�T#wC����yQ��Z7o9�{�ٰ�qT$��U�N�D��9���c��F6��fL�&��
\>���ci��f�7W�N=@��rz��CJRS�T�k�b�:�b�2)���8kZ�Tu��ޤH������񏯶/){�g1㱅��S�ݷr��������u<.ip5@e�<���h]@vq�_m��J芹���-ER�z�����6w��s������(*�D��{}i�酊���%�Ses��4���� ��!c�4�ػh:s"�T�7P86#dDO�GnSa��jm���i��ɵV
AS��cŧ��v���4���J���	ځg:._� �-��Wu�I^��US��W�[��5'��L:i��4"�t�sa☿E^2�f��wK@�!A����w�������gV��)THЀ��PF(-�q��
�c^�1A�n
3#��hK�����d�$��|Px�bH���faO�Z�/��.Z͸��%G�hI�(���� �M���lfN�$x�_($���_Y�(UH�Fn�K���v��0>������e	��4C9��n���Ң�_�U�`�b���GW�"�{��s8���#��D!�h�N�-��'8�+#���}Z[�:ܹ{���Y���:���.b�����8j�DA���7o��>;��f��X�w^���[�F���/�3a^�ÀIZv�n2�4X5(:�����[�L���ڮ��p{_!|�A�z]��w*f��wJ�h��Z9tkgDU�5Y�RE��	���X��2º��Iރ�U�e�w�;�4t1�T�g����ӌ��r7=X�ls0���A��	d�4�	�\<��\yo�ޒ|ZP����:�����r�{��V��;MX����n�B�.��~�\G��-���+xª�kQ>1����p��%��qlR=��☋զ&a��Ԩk�t�W�������<��>�IX�(S�����H���v��;��v���I�b�C�ݰ�QA�W� ���F0�����2�uֱ0`~�XN��	$��S�����&���,����d����Rj�<��t/W�u�pL�yptysA}+��1���R&9��d��|�Ȫ9ӐG�Y��d��=2.V����ZR9�^���M�O����S[����⼳߁bq�ٛٿ?����q�ߞ�p6�bAߤD�Z)�㒽�iʳ��.�/@���x}�K�$TR�Ȗ�k\\G��x�DuU���Ҥ��És(�h"�Ԁ^u�?�譣�wF���c��!w�H�V��o��y�ј�Jr�;с� ��<�cPAײ�+����@]��F~� 1i��"��0o�r�Ө��s��˕-�N,%�?D�Z(9l��q�?�ol�>���y�3}6���^�[g�P��6d�z���7��I���ʒ���s5s��9F ��&l�kQa���h�CΠ���"
��7IM.�;U�I���.G�z��t[E���n��w&Q<���ޜ����y�'�#
�ݓ\lN���_�3g��S�������$R([d��ƪ"�+��6�It�Q;P�R���u��DB����=>��7��7���8`T�=�>��z�O��he��`�􌩒�&-�&F��$q[z�n�Ad*!p;~ˆ�[�u�|C1��7b���e�~�:V+c���w���	e��u7�b?�M E;�e�rL�c/<=��]S�ʍ`f�h6Ԁ�����L_���@,ߞgP�!���O�2P#� ?����E����Z���N.��y�>8!�nxhS��ٱ�Թ��x���p1�)s{Q�<� ҄�g�i�ĥ����.Nt$y#�$յ�t�b�6�;����T�׏���ɐ,�7]�q�K]et�����k����7M��<��}��+�~�+�$�;#{�y�K��N;��!wp^*�C�<F#-P���V�������He�!K�Լ�{8]�y� ���p�nd��q�S�ю�~;��"J;Iz:4�ʋ��-?��(w8�����\Z�Wқ޾�����hH�9������L�?��	��B��p��G���׏^�95��9T9��c�T��Xۉ��a!&���9w֪Y���H�d��ێ�=�ۊ��eHo��(e��"��/p5�]-��-�O�+��a��5�Sti�Wh�3�(W�_I��H03�ah��?��\uF� �o"�tL8�k5�8 i��p���2�s��Y��U6�ƪ�o��Pbk��v�ڛZ�h��F���9�y3�,%SБ��TKi�� e�	rZ�|��1�	��n��a�cGTIv`R��kݢ^�U	��<w/_�}�~��$�G�x���D+τ��Bz�দw3*S�+���Tݶ����N��|`�}���E;el�m%[�5L{��[i�zL��<?���%M��U�ʇl��S��xf�Le�epO�;�eO�҇YU�@�'�Z3ܲ
�;.˦,,6CW�� ߏ��:��v��j߅xk�FLOem:�h8V��(���Wh!�_�r�y�����
����'v+mib郼�בn�$6�ڗB�j>�\�aco�) |
ep[GQ��A���� C��@{�s��?k�R�9�8Ù����wQ�̉#�x��\�t��s2ge�S������9�q��z��bUA�鎽>�2�ٙf���$
����>-g����y�'�'*��6��l�ܽL�F��/h�*�"$��ĵ�t�n5�!�&RD��B��}T~������]��j��.$�ɾT;^U�Ƙ����J<\����ưq�ɛ���X��~�����ѷ�[������[�s�W��8 D���V�D��6�G7�
��Φ]�.�ިw??�߳����q@-��R{���X!hB�����e$��\�v�$Q��g6*abK���&-����j�ɸ-�~����
��>�,h^��e�\<#�m\$�|`0���i�t��ՠ�Q��	�(X��RNL�u� 	��\R��CW��#ԏ~�f���0{�����0�Y�k~q�.ύ�>��0&/��&C���#��q�Q����%"BS;%Ğ���Wl նE� z���,ܐk4��T�z���
����_gv�tNe�|�a̸κR���~� N;`9�:% �܀b���:t����k/%lyO��f���ź�7���7GJ�����$|�����)��)v�-z�ˈ�)�2�Y.��i0�,(w�G�g��e�BdNI	�0U稘O��<ȿ�n�AR�I~���4�MX�=j��ߧ��pڊe.�A'��9�NnП�O3\����
 �]|��)k�+C�q^�(l5�12�V�ι8���F+D3�a�����g����TJ�8�S�M��l�Y�/�2�)rK�)�o�Z+,Բ�v�)3I�6��.n;e��u�Ԥ/��@g��3�|�M&�9%$ST㶖�dIr�H�_B��m�,<T�+b��<vu��!��1�Dv.u�\8�^��]����E��$��w�#)�!x|�!6����^��%Y��g�k��R��͖Q<�sd��?��t�3��(�KT�{B���T\���s F�����}}���ú%��%ʻ����^���.�<a�'�jT=�Tm�c(����蕕�*D��LÓ�;:�/��:��^�'�є@��+���JV'�$T[h�Q�ZE��?�!c�o\�EoK9ƼO�A��\�Yl�v���2z�Wd�v��94�.����Ĕ&�(�+MjE��d�};!��Rx��2W��p�B��=F� �dc?j�xr�	��Y��*��aUv����.�:�5b:�C�@G/�Ď���#�ۉ��p6H�]��n���?�u��+�fc�(�6ã���T��_�8Fˇ����%��9�A�nTg��e��9�LON����cA	�-YI
^sM��֫'��a�y-���+�z5$��'�Û�ԋ��@#� 
1b
�/��Κ��췧n���U.��a.Zv����S�.�Jۂv:qWb����|\��a�ˇj+nE�q޶�w3�%~/��ae�ܫ$B�S� *�,��I�
m���k	"g��b��%3`i��������gǁn�l���'��ںFi��lϥ�J�"�,���L��\�L�����Uy�n���4S��CTN� �"��L�`B���J�[�����ҵ�gD,�]�!zr A� ��+��YX��%�����V�����En$!��#h����'a����"��GqK� �l�ƊJ��8���F��<Ե}m���{�U;B����s�����N���Ŷ�W=�L�"7~��4D`k���[[�	�z�R3���k'T��lqaNk��	t�h��.���#�V�sk�	��m -��K��y����G��;��E�c����p�xn����{��3C��tp�������m�~i � ТsX��e�PAh�|�+QF,����jj��<�׺L��2�-%86���{�/�je��xX��\6��im���f:do��s�)h5A2�|�!{�)��Zp�	w���H��AMbQĪ0�#�xb�T�!pS+����������k!��Ưr)��`�c�u&.� ���ק��FqG�e�g}o�6;4�z������_aJ��s�}R<%A�&^�>ʹ����GVH��yIj�E�w����'T[k�i���3
V�{���d{2<2�!G��&n}<)�qdm����� ��ݍ�����pm���)����Ȇ�V��&��L�D��s�Ǯ���9/{?�0����y��L*\@�`��ήﮠS��m|���h��� �ye��dNڡ,�CM�&����Ko�y�Of�l�V��"C��n&��EG(oa��>.ߨ��ct�������׺�w&X�O�*��-��{j�HH��~�&9*�2�n/�MQ=J��G�������,�'r��%���
�K��~���r����Z�EI�ߍ�-߸�-Y�5�!�Wȝ��[� ��J�%�V-)&kn��@{��M��j^I'e�J]䧮����jV���m�W������4����	�?����~����Ii�vq������5�!� ���Av_���w���O^Ha!���|���^9򃯶�����I4�����P%�����w�l"�~JĂ#�4��mQ�-Y�H�;>�XF�e�S�����f���@;px:g�~mn4أő:"��۵�{��Č�}�S�7��>W-����br���)��ߐU��d��[�|��w��~�q*�ϼ��ٔ���U�hx����A����gN���:�Yp[a"=�8�u�Kgn���
=4 kA?��ԝ��-�ҿ�yP�:����e�R>]��h���"
��#��&uT.��5�ԡ�d���@��X�&��i������Π�b�a{X��a#���=�������U�eT�H,�����$Dvh��/I��g�N\^׾�k�Nz����@=��SO�2��IH�sNK��r���U�b���Y�*)��)48�5*6�"!���{(����b�sL�˙w����]��n�G�_�[(,ƙ����w���Tܪ��?O+��q|�1�4 �T��t�7��4	m	lL����^�9��^zF�t&��C�֪�de�S�W^�}��-bV!E�K�}{O�� �u:�P7-Ey*7����i��|7|9F�{�!D[�3u)L���4�P(h���Y�Ō�m+���\I����ev���S����J\�盀<��UX�V���e��.��G�'�=&�mK��Eu��1�:��~����~��[:�5����px�����&οѱ�]���!�ȝ�Ϫ$c_�X��
 삕<.��d-��f`���P*�f��W&b��L�)�@�o�[+1��։n\�mr����Y�lF��K�
�WNӵ� �2*�&�(��� ��M��3�a�[甈���
��'��-A!��Ո���ĤM�s�˃�{b�+� ����v�e�I��2�69��cDщ;�`d;LХ�|^��2M���4ݿ�-�Zfk�7h`kn�a�1��R���	P�all�c��oJ��|��t?�BGY��-n���6��?���pad��BR!���rP���\���`����|�H[�N5����w��<�p�|=��8������Z�w!�rP�l&���nby�qaST�L������(����S?����^eȄ��[���mm�=�Ot�����;�w�|o�o(Ki�/���3��t������d���7R�撫w�O_a� �yu�lɬ$ݓ����hA�Ր����|y���r����mH<������D�@�!̉!3%����-��)�Kh�aD�K���+��`l��I�P��
p�W�I�_�~t�	5��Pֺ)Q-ܵQȢ`>Z���W���nb�gC)tȐ�!#��gU���B����y�.v���ԛ��d�K:�OZ�b���& z%ׁ)��a��!���y�Bs�yN�9��moj"����M��S~~�z����0��E�n"��e>�q5�з�w��D�q@-N7���'��,�4%��I��K5�#���P�-�z����T*_��܎z��w(]Qʱ���+'m&�s�Z�!�����~P��4��gz&�1R`ABe}_��qO�`oZ��A���hםH��'��^�Y�gKC=I	 �C/9},ߙ��!o Z)�I4�������i0W`.�R��0��By�!��y����&��I[�G����xV���Z*�1ao�o������ԁDZ�����zYYp.N_V��%�p~�X�^��)9hq��4q
ǉQ�-o�Bҵ����	ې�i���H6��cT7�"s������m��׊�S9g���u���oNT'[��l��:{�#g�	e^J��`�wTh�)8�鶆9��fP��:��p��P��,��a���
;(2ю1�J�Wp��RU |[�+#�P��8ڰ�����.�7�I�*�ei����)�չ�F�i�,������i�	S�������UdK)��S�$�2Õ3_�Ҝ�䑢Zn�o<�#y�ʖ}�?�[��,^s�*�����J�Ά'��\��#�,_�`��Bm]�UNI���1���(���;#, �m6��w��_���}�1/D�:��3�C��m��s^~Q$�%��w&hL�*��Z�J��=�E�;�oʝOK��R�>B97!�q'`H5��?�o �͈�'��f+6cSR���.J�?$Q�B��߂�f{���=�f��;��%����xq�jU��
��jN�2,�q�6�����R	��T�(Ђ˄����д��ΌY}��d!�MR'sl�'J�\�n%��iC�����,�`|�-����(�wAas���&���$��O�Zӑԡ!��ig������+"�X80�������̟н���&�\�7XXzÏ�(QV������kc�_�A�� q�$�=G�-���Hf�e~���,�*����	�;s�g����y,U,���!�P�Ԏ�z砤ٳ��,��?P֢������Q�La��Pg��R�$Ȿ����y<���?�_���ㆠ{0��ǈ����*�MN������K��w�th�"j�i{��jRaz�� R�'4�)&�~:��J�Q�/$�>��i4�%�v*0�^mC[W��� �D����C ����.�ַ��u�+�t��w����[C�ϥ��}��K�U�7SOr�[m�����\��Ȋ!��H;�w��t�M�/�3<���M~�+��k��A̜��Q�M�7o�)wWl�"�����%}�ɾȥ�8w�JIS��D����o;\�