��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#��y�#-����H\rD����5�/m���%�ȳ�Drn��K�� �:����WIEr��YsL۫�f��O=ϳKR�2j�]\QZ<���B����	:���>K�D�%����������"ٜ��iLG�w4������Mm�R�m~6$m�*Dd�b�k���� &s���r�}�+0�?|�.m���b%��?L�J�t��ݥ� 05h����Pz�����􊮏�UNXp��	�:cG���Mu�~)����%x����/��M���	�	�Pb��0�~d}y#�+�c"�p�Y4�ޜa+��}m���4�0Pá��E'��A<��V��m�0r��w�Tj�? �+^�vj7�÷�g�#�}Z�P����,��̧7B^��2�t�+I�<�MU�7�e���R��4\u�¼3^���]�6��i&?4&��d\�f'���0�m�5i_>kN}� �.r���چ�A>-�l�֣�X�Y{a�Ij�\�3�38P��ϸ���
����M���04s�рM�� ��[�JC1Cg���jZ�G����wvd>���n���?�:�l�� �;��
��b0m���������2�E����4��_9y_&!�O0!�r�Хh]ea|�IY����h�UDu⍑��}U�S2�u����>Le���2���x�(Y��ʮ0����E���E���l�~���Q$�����T';v]U��"T�J��ȟ&_��0G� Ș?��tcQ�I�kӎ����+"x�1UC�`�E?��p3Q�i��Jɳ��2ٱQ-�'0�[l��$z��)D��L�*w�*�R��r�o�Vc��.'DTJ_M�+��}s)�V?�.���,Q�cQ^;���K�#j�d>�_����]��>MO��@5�d�)�g�L�{C����1!#����}�h�k,A�t����7��1}�f݌��'Dô[��OCu�� �~h��uo<��㪆�/>0�
z�`�P��XǛ'���3gvi5��l�L�L��_���E<�7��B�'��0�B�zI�mս�qJ���v��/e�џ|ҳ�}.��7��@��6�}�o^ ����]�c�r桝��U5��1�D��%Ė�JB�w97:���*v�Lk�L���땦#u2�%Hv`�5��s��v7�^��nN���-���@^���;ҍ��?z��P�b����<��k,����/�ˡiH�[K���{-�0J��,�C�M>��k�	P���@	4&��q?��������4 /��j��}�*)�}iKYUwR ��k�kg'��W��UF��\Y���z\�!&
�!��m�rbt7���2��c�|$LXqb�[
X������9�~>�9�u�{��j]��z�`hf��%a�,�<3�o���+4R�;������˟�%��^�/��eƷ�Q�>��g	��=�Z�����h;s
����kx̎V�@���kPtH�x�YFX���@p�DsΗ�a��}0�Ie�g�E�9�+�)�'�_��1�L�S�c�S�Ŋ��mA˙ϥr� �ϸ'�+>�i��j^��Qè��B��V�E<�����M?���{}�tEX�l7�K�Z�t�<o �4��,'v���D塳�7�_3�!�jp~�Ev4}=p���!H{�����vS_p6�I��mN�1Q��D�Ʃ��s51~Գ���VO���2���^V_:�b���ꠖvd���E�H��J��,`'�+4bp�D�tև���V�{D<���=P$��PJz��ۣ�����x�H�I���?@���[A�b�ĶD�	�I��_pb'`�C�_=n��>�D�M9��3.Y��2�(�i�A��W�$E����;�3�(6�	>���K��D�yժ�I��:���7��5wt��m}�Ѵ�^�{��+�������ю׶W�9y\���]�NN�j�7�)�,�]�z/�b{6(^�h��3��)I`����Q���`C�P=�10x��6��a����{H�.��Շ�3IS-EU,���g�Q���c[?K�h��x������5+]
���qA��U7g�"`�3o�2��	�kK8^H��V�mjm��4ڮ �=�ۖ�$	/�i�NHX���UYRv@�nUJK�N}�|6x?�%���D4>����eI ��.�2����=A�o���R�m&��g�q�l9��^1�e����bIw���\� �ꭕ].֜q�U^O��ٍ����}�X÷�3�%�K��l.o��C�.~��f�?�*����f����$�&u�Q�����Au�{���e�W��v1��ץ�aE5�����|r�A&����M���;���c��9$6f�g` �m�8�(�:u�~�FÇaȥ1���:���V"vD "��ٖ�*�g`I �8��/Lx�j>�k�ջy��*�؎é��w��ˌ�k��;�Lq�q�|���Cb�5|	�&Q��N+�;#U'A�}��|�0��;ضv^��ڋ�<���%�|�g����[v�j�ᅄ��4yO���/egJ���$�;�O��3��u}��6�t�\�7,,x4��E=p�hnˡ�H�N5�b3�92
��k@jT�n^����"��7����x�x�ա�8��=�u���p���ҽ��|��`? �菀����<\\w�7��Z֍f/^#A���u��&��+L��#���&3S�E��.�����M��!u�U�ʿ^���fP�IK+�j$��j���9�+����p8����r��i���n�|�����E�:�%fX�7Q�2m�s���䷜�'��r~6jeM�{�tU儀�%/ݷ[���e�A[/Q�B�����X��WWp\����-�:��H
w�`�xk�17�8F{X��Ր:�Zm�����N:Y۲�P��ZL��V}h�F�/�P&O-��Yi?�j�sup�Ǿ�9N��W�i6/ɍ�k���R�W�`�:�ζ�[\u�7�B"�4jt��[�l��aS�Q�{���ȫ!��	Ku�~%��ؠ��І�'Ju�k�u?�K��������{R�C1�ڨ1�d������
 ��B�ɴ����x9�M���L��.�� &�`,��Z�@(�9���Ea�����ƈv�3_��H�Ҭbص�X<�h�)Ջ�����fL1l��_���̓j0�s�I�L�?9VG>
�V�]}�b�,���$Ѝ���̺�5�R������<�,:r#���'��)Q�7�>��	J�2�嚮jWPЫQC�58�H���)�..��7���gU1�d��jE���
����xs�F撿��Ӊ>-pX$b�G��ӛ��s[�Vbm����8��N!���-�4W)*@X�8�r'RҶ��oc����)r� ւZ�l Y�v�w�RRc9�F��u#�BG�M���N�o��
U���\�w�¡G�':�x����?	�o6Vv�_�&��x(��Lv��W�*8�P�؅'
ޣ��7��+zY.*3#���C5&Mԁ�_�������%`i��Ӫ�9�&�hfs�K5X@�R�<�Z�����K;��x�"b\��.V�c��=da�PGw�M륕{�Gb��X�E֕�,'�}������Lʈ;>Q�v%ϤlB�|����Y�ְ��k�d��U��J�һ��� ��y-sZkd�(�R�z�m��TQ˸���c���=����.s��v�Y�9��;�'�Py�ƴ�yl�C�g���$Qq��| 3Ĉ8��3�̾UE-���2�"n�+z�er-�iū;ٔ|��Khg�-�_��쇾�jdI� ���Q�Z,I����+�w����6��4��G�v7L��;�Fe��pg ��������9���8j�Ɣ�[�p
\��x㹸�Fj�5�U�%���w��o��1x	��!��<&�T ��b��E�O	Gv(����U��>��(��]ۍ��{Lu�1nu=�k�Ԝb� 3�����©^�
�B9O�����.�
�k�Dph�ݐb�Ƽ�0H�N.�? ~��դ�i���߷�@����;>F��c��w��䖄�{�E�>=����f�����ѧ~�C��Yj��M�y������>�Ogo�50~���RT,���8Y�$[�M���L	����>)R"4�O�����HnF�6Y��~�Nb��3rX��D��Ǆ�t�e�<,��$T�D��O�K̓�Pnp�p+�:�*j����؂� ������qBHOW�#S�gr�n9�f�F��ۓi�cDR��ZH�Ϳk��o���Y�������'��w�A�1��� \=e4g�gv3\�[ظ7�i'�U��� �x�~0hg�Xxk�o&�P��ʅ�t*�+,=����22&)Hg���Pj����F=��9������Wj+�������&!��l�$�U?��"��N���t�f���ă���K�w;B�f�N� ���Bo��*����,fɌ���������%�?
Ѐ���Q;������dM����a���H�~�����Y\=�f�:���(����'{R�w������� ��6��~9\Q�8�� E�ſ�����B��*���n_)��R��|{�6��`�⻰`k���c���ֽ7�����U�Nv�J�����������AT���eg���$\_�f�=m�mXFV٦;$P�m��	�qBuh�w5���ʣ�Zqm.�\W7�:I}ǫ=�|؎ZfJ��T�����CG���K���rg�k��7k�����w`y�\+��z�%�a�A70�U��y��`E/������B�ퟵ�~�����3�U"������(5�Yr����5�%��ڮ���(�g�)�W�ʙ���j�:E����>_�R�=t+�tL���)Pt�P�\��_Ls�� �b3(w��Н�'X
�B�w�d9��>�Ҡ��ӇO�>��#F������Ւ��M9�Acs���$�<buN�`1���_���G�8�&-R���Ƚb&2�1,��_[;#�H�t!�1|��[����Js�����X|:$8A��޵�"r�b9� tW/���Gu&䁣R��=pY5�Č��qڀ�����sUa!����*����}�cT���Z�'�Y���f����Q2���� ��+&Ax�,GX�9&��1��e+@)Ӡi��[��;���EV�B��YSk%R�L�����ؖ���k=�8�xR�(F�X9�j���\���Ged�;�j���ʇY�F��UA�����W�4G��z$�\IL5w���˺҂��~c��(��rg|~J��7��O�;Ҭ`��]8enW}:���z�߸�t�W����QL�¸q��RG�ŋ�Zh�6���"1��(Ҙ�=US耖}3��&�c�ߡ��w)�ٷ9�ۧ�#+Wz=��Dn-^��Sff!�zQT��� Je��E�͵p��>��z�)�^��K	�}K�i�5잒�fM:;;�y�f/�[�7��QQK[�d�p��B��e��:�XAcR]&�1;I��@q��6��i�*����C�4X�����ع���ͮ��a����Y����r�h��`��e��Nn'3�<�^r�,-�T�����yצW\(a���=i�B��2Y��TB-�ewﲃ����
���&p�; �WF��CR}$��6��c���	!!�I7y�K��7��6[8���V-�Z	
)��&p��'��]�"����n�{}�'i���ȸ��^C`�3�8��W1���;:�*`�g��m������w�5E�h�
e���%�k���Q��-�]����#�ÞaG�'��s��z9�,����s�J�`��g�19�M��"����"�u��s8�h�"�r��d!�m��un	�_�҂Z-2���$��n��{#SnzE�!I���-p+p����0�)�T��_�Z�5VZ��3*��[xq�gV�ѮU��o�Jv}��j��(-�X�R`���y+�L���;u�D����f@��9tf|�c2\��ߊy���-K�;�yM���z�$�c��CnL��^~z���1aQ6V+�г����Y��BPS�wPK�Z�m}Ho=�E�Xj#M��N�)^9c<��] �ChuNg��V�U�O����U�<]S�x���?K���(dg�c)��D��Y�ž"Pl�1�+�ԙ�?D����dM_fN-*�X�$��>������@�*@6���E�ŕ�c��Pr_�o��~�w�=#1�c+J�YM��V�7vZ��Gsc_I�C��ʃ�{f�ա��ɛ��9�J� Y]�M�O£���n�՗����O�٥�g�Jk�?>9����{��C��^���Uq�C�*@�۵�Y�1�(�{��h�~�bS���E,(�#��}�SYJ���Uv�w�t3�m��6j�������qA��U}̳�� ���l����ݛ���)7>��XQ˽�ȟ�OR�@}֑\}�2��j2с�
�.Ё�c��	�8K+Y�q�Q�0��3G*�Rs��ē�#�0W��(�
��_��҄I��+�"���ȓ�w �Ώ�o	�i�&)�8!M�
�t޳Im����cڂsGn9�彏��� ��}~Į��*�)w��"���6�h(H�Pԏ�[�./���!m-�e&��wk�>����#v�@	��s����q���|$h �[�Ԏ��fW�iԸJu���Fvn-�x����o� �G�3wB��!V�F#oK>�@=�n'}��?~���d����۫|���z�F����^�&��o5���d!�8j8��%�W{S�Āน����/\��w��}���e����gM�C�\�׳M��Ґ\���烼D��(!��w�t�����&� ��ܤkx|m�$�2�G�*�bL����E";eJ�_A/R���k[ ��M����}���|���¾&>�sz��t�����o���2-�p.Ps?��
����󘨘�krX����Ƴ�Ona:�h�v?YM�R�8��ظM����<H�wFc�'U��t��X�/(G𑠋�Qj	�gL����S42�%r)�I_i{��(^`+X���z���S&��s�6Ƿ���k�TU���}?%'�Q����h#�~ܓ����܄�~��N�7����Ǫ��{��\����Z���ko�E���(J;|	��{��G0��n��g��!Z~]��o�"��<��S��ٖB��(�;�c���h4��+�{� t#��|o������D�
"`�;?�w��2����B���Z�ԨFI
�'	��r��:�x"��^{߮}<mQ���D*��EUTP�"���З7��:?Dםd+7)�:s�s[�oO�w�jd�����H~� ��/W�&�|@�-6������Kh������i<:���t�ꁞ��/F-�����(M�(�@�u�Sa�	��;*f�V�πZM�ANh����nh��b&p{�S��KF$o�'� O���GSŞ��m"��B�����ۄҠH�S�t�5����	�n��\ث���\�&ig���e�gj�Ry�v�t2w��:"�iɠ� \�.���k+�  J�$t��p�:�Oa}�*�y㚋��*6���Ɓc3����'Z5?��à��$5l��Z ��u��� Mԝ�v���k�xTG����:�ǯ��l������N�$ə�ط���Su����u��-�nU��|����[9�u�>/�"���b�ŪPf��<QE�	���O3s�G����v�t��X�����s��Q�bv��<��.�f5���;Oki�e��U��/�!q:����x�S��������O��n���5�傸��04�Q������Ŧ�Xhr�+�=�bm��r�R8$��X�j�R�E#�Բ�6�r�J�� �TY��a�lO�D���ܸ$��zv����
�Q�Ύ���9�M#�B���Ct��V�S���2����<Q��g�����<��mo�05��ɰ��2�v��xۣJj�e]�"�Py��0��֜��f/m:������콬Z�v�tBTIZ��j_���$>�u7�%K6�r����LK���ӓ�*��y�ͯ����5K���ܟH�;���ķ^��<.z�i�}���ä��t/W]��>֥����~L��F��j�ۍ}s�G��۳W���ˮ3r�D����q��qԬ�1=V'�C�/�DqIpu��99��{�Z�ɏz��#� w��S������a��}�ҿrR�p�n�`~A�jkqmK���ř��G.ڋ^���`��i`q]���A?��̈�އԴ��?)y40�p8¬��}�!����m����f���E��k�9���}�k���߾�����*Vp �H�J�EzV�*M��ZW�ȟ��""�7�K�.uu��I��-|	 �/���'�85$��6(���;4L�s~Z�Z�u?R2Ua���=jܳ� [E�􈑋���3��P��}Q�O$�ѥ�7M@��Bm�I*b�ğ2Gz��`�?�d�@������&^2�Vx ���(��m�L�R���$�B���i�C$wf��p��$)pew�ނEqsz����@��P[��5�z��~�f-��)�_g���Z��� Ĭҏ������N�c2�4�Js��z�����k��d)F1X�2xK8밿G@Og�C�֜uo��@2�7!3>�Rm/�W�A`�R�����-z4t|��ʣ�-sʅ`
��_�	)�Kr|�e�{W���:epLC�#<�<�V߅����Yj�yͽl�5��~N��i 7���SI,n~L�H�1��߷پ�C~���>��hJ|=�����������5��2�����f��HG��6b�t����&�ruKk��eC�Z�8���c�c�ϭ�i�������a	 �'��"��*g�g�@������e�{A:���(}��^��Fظ�b:�5�I]Ҩ�Ec`Y��M��E���X3	L���)2�����ۗ��Mᵂ'�>�p�Jg/��=D�6B;�qTt �K_���A~��Fe��k,@���<C��B�`v룤[u�TS��	�$yOI���x�X��S{a�S�R�(Bɧ+p3���/~�򵜾�!vx���z�v�q1%���t6g��vn��7������#v��dE-hp	!a�����'�Di,x@b��b��p�s���|�W���-s�_VZ+m?5<H���˟ 	�Zy�CB&��H�F��dJDP�����e�@����[4��D�LI�.��K%�V�r:��V��
�@f��Ꝟ�N5�!��Ïf~m��OS�ۗ(Lj~��`�ɗ��8e����[�:o�ٜUk��������8�V��ɦ*���I�
ݯy���rV ����1A�.�pF�{���8��'$"j���@1�7�k�/��{����z���x�v/L�G��9�g�*e�S�}�B)i�h	��i��fu$�.��!�42\��b۷�[F7lQ#R6�x���Aw<ô�#n��jp�F�ޱw����H�WA׃K�]	0a�=�4=��s�!�y�O� �GF/N��o�"�[tH{-����ez0��KJ��p��p����j�A[�
7 �U��2���u���2{u/�s�:�7uT�#V���4,`F��A�b�qB��� �Hg���/|���f�3s��=}�	dh�^G�6�3o��%ٞG��2dT�B`�oc�i��*�M�jI�PU��aT{���.E��u�~�%����&,���ٯ)����Y��c�2��k������n�Q��8�$����� s�� ���;:m�R���-7��\�hbXSi��4�3������ŪMb�Hu �1g�\�0/>����I�~�cT�׺�1��p�G�WM�fs��ڱo�Z�m5߂~6�_吱��/�̟��"��l�X�I[7����$�?g���}����
��o��>%-M�/�$՞���A�HZ��+� >��HI�Yf��8��R�zv��E*5щ��|M,�)A���������L���;��W�8����/��،�n a^��	í,��OP��\�ь!��31����?MÑ�-��y���@��&�,��� 4@�Q,�JFP�o:����Z��T���m��+�Ɩ/TS�O��r@�`�	aP$��@v�"�n�V�͗�[
ڊ���]d�k-6-Y���s�e���H@$U�l���GS�\��a�s(��# 2Bl~�"#1����C;,X�bΧ�LYe��ψ���=�&a�Iߤ�NK���LhQy���/����tay��[�M���uN��T��A����8�/eQ݌�ǃKk�$H��m~tv�����Z�ɕ���(�M"|s��5��$��G*�6��$ ��ҳLR �\��:�'��[?��/�m��:���M�.&�"2�l^���g"����-)*�f�|�Ć&�)'���'�f����'� i4~��GVI6�4#OT�#�r.85��2�8������e��8��+�)8]v��i�����ɼ���qcyr�,���?��Q9�������=�&�yE�}[�߃����j�ɲ��iR.>��OA�Dg��j��VD��W)��e�f<u�����j�dAj�5nuLf;Fqylc�tl��0+h�3��G�ת
N�(�����|8����W���|/H[
���Hp�q8���G�5 �����~*��D�"��#K�����g8��ϊ�� �Ӧ�Ho�LG5��a@�	 3�@.�!N!EjQiH����@8�"r���z�x��A���ٱ���@�a(��+��΅"]�~�^�:��9[��f�=���:�"�}ۡ��Qb�9�F�:��q�ñ'|!����'Ri4����N���9�{�u m�aK�w~Wn��0�k�}O��� q��L��/�� װ��q���//�9�o���n��u����]����w���)tf�bTcd7�7���X�C�����E�(��V-PqV>�:��l�t#�O���7�Ʋ��YN��?����w�^ZHlާ�ҡl�>��1P�"�O��'��&���Ιg����1��c�Ocxٍr Ĳ�I{y��]������C��d��U	�Th�7�F2	q��{�B�X+�;�r����=.x&��&;�Ȳ��#K�4$w�u-�J�+�����KE���7p:ЍY���>�z��A�	[�-zF]���/D�f��� �����>�EF���Qb5���.����#�o�IG��r�h���;�+K�<Җv3�mS�%NTO_��hn@�8�<ⲩN.es0E��N��k�V<f|�J7`:Ҍ� O'�A�/���8���լ;wlBRފ�2�M�5�{¤�Sc��bA�Yi%n|q޶����Һ�/�^~ܝ���#�P�x0�/]?��0��t��D��7�4��X���%j�V��8OS"J�̏4�w�����;�osqy�BTg<?]���t�b����m���Ӂ�������ow&!����q{S���j�����&;��y�Vo똙6�/U�0��u<��8n�{G��4�ٱ��3d�7i�I�11�{�eS��qGggϡ{�:���*Gm�I��h&��l���S־�������i�!���a�q���A�eV�7bO0��A{����_/F'F���N��e�O�m�RÿD���/+���&7z��a;X[��I5c`X+����@����I5��	g̍�j�5MNsw��H�Z�y!w���$���O;��M�}[���.$f��$c7e�-����I!Hn��"=�iM��H�X���*]7��p��q�٬�W/�S5����vr�0�s���J^9H�3w�4ǥ�l/�E�d-�����ا����:G3�EZ��"�1<[�}^\��쵼�R�*���c��&}��r����Habf��W�%� �QcA�p��I1 ��^�QZ~��׭��~R�Ctz'�ǲ8ֽU=��YV �}F��,�yq�Ԭ��cU�D�Zꇗ��)�|}+��D�I�
_�9��«�V���#�]��]l�ԜEN����|-�<�c��������1_\<�hc'v�͍D���edVW2���rt��MN.k���xe�q������CW��J�=�g\�ֳY��WgR��~C� ?��j�����j�.��\b́������j�Ƣ𚹎��9���]-��~�Ts�`;���_r����b�c��&t����6�q�t�<(}'!�j,Y'���k��ƤXS�&��S�!A��ץ��isj�������b �x�8{E:�lE��~~A�3�����+��z�z+������l�p ���L�FM�&`�ޕ��(�՘{�:�"5����� �����%��Af���&�9(
q���Y�g�qL��r[���e�����zڼ����٬�#����;�bRç�q*I��y�8�6u�Uq�?Qb
4[�z�rP��=5w��υ@l���R�	~'��/x�J�bSN�m�ë4q���T��:�HG�M�i���,(�ċ�*Bw��m�P�е�9ڝ�ŉ+H5���~�~��M�X�ԗ��S!�g��6P��-rkΈ�al|���<mN��6�ν�Z�Ya�X�V4װo�n��?S���=��=����O/h� �]��#I*xA���*͇����}�-�b�x�TQrԱ����R+�U ������p����;�.1���Tr���[�Ъ� ��xMV�R�xA�y&F>���"�"���e� @�'4
�������"O�yH�姷5Y:�$\���x�樅*Ts2Bl��l@���K�AA-x��/מ�3ѵ�I��D�9¼�٣ͤW�2��Y\�$�Y�1�\q��1�}Ң7�u:�j���91O�av
�������\���D=�BpE,�&�q��V�cjXd�x�W���I�s�u.5�ޓ6\�I9��_�ϫ�ڨ�'�s>wmd��s��q������3�8R�#l1�\�� I1�	��n��u���>�i���#:�����"��ɕ��Q�<	Lsl*�Z�?��1qs*;$�3����^ ���" w�I�T�#�ɹ���S�fL4�2Ӂ`��ܝ�6�����E@·T�B
���L3�:� p����ՙ
J^(k�gna�%�:𥃄��9���rL���)���H �a��1��Y��HNn�������
�`�d�1Z��놟@�QĦ��:�#Y���"�+G�@k�Xz`��E3u-��u���	�{�|�����3�"�=%^N� �U����R��wTxmh�_L�F�����S�ә2�T��Z#!8M8|k(��B{F�P{�i|nu�쩸xU���ώ�@�Qf��"*/6U1미���o1~�����U�� ��St� �w��Ê�dd�*3�/嘈� ���S�c'kLa8rk7)��Q�[\��Ts������W��Z
��8�ܨ-��)��#����1�t�779;��bU+�#o6Q�8�"J�݋|f+@Z�V7!�E�6�� ��n�UÔr^��A�<ڠvS��M��>�Z���2��'v/T��dA�p�,��H�{A���T�2h�[))����7=а����B�)��6��(
j\���V���RL��� ��d���d��So��Y�Ě��} tn��ɾ�=_�=gP�5QϘ��L�ZՃ6�<�i
<���V{���2�O���m9���L�L[��|2rS�]���J���k�{Г��My�f�I��\�3y�v�q��\l
�-S��]�����%�߆��̪��f���~�}�jI�0&�����ۘܭm���Z�x�����k{�1�!]a��b)q�n�
 �q���)��&}4���� k���7א�M��������^PJvEГȇwu�]�8VN�0�@�iK{
ǻ�;�����,I�N?ꊦZ�������9�h�����}a�#��De:�ֶ����<�	�o����	v�*݉paQ�E��Hd�r����I��ِfP��0 ��9 ��*���V�]V�a���K+�X������=���O�0��VM��-.!j��P���i-Q+\벌�\Z�q�U�
���tKl�0�1�6W�q	҈҆V�Q�J�]�
\�u�6k��@9�k�	�$b�r@�$�O�șɫ���Ԡ��QQ�'DH��-K�HF}�+۵lo�ܛY>��N�JrK�]�bZV�|��Lk(�k��GѮ�C�^��l�N��)�d5�]��-3��P<��p��pcuz>���V��XO�p��iyp��k�J���H���G"4t�l��J�&Ʊ)����2�g�_�YA	��_��/��O�Y�]
��#T*E:1��<��G [߿��XlE<���ZVٟ�Ìi����q��2�	�qŦ��0�|]�)rK�Њ��4��֖�il�����4�C)�w[@Ԧ����y9S񦷻_�y���\jD�r�D�}/q��^�UA�O��UG�^��4䅯[��V[������A�F�=��_�}>H�ej���I�z�:�B��jh���/B�N%5t���D�'�dY#�2>r��gqI�wdog#7?�>�(ʮ�Q��:F0�"A��{H��7�]��=L�����3��n� ��>�p��L� "�g5l;I�dP��Z���$�|ք��� /Y�M��y�u��A7X��h����R�oQ���L/�|��W�K89�8@�ޔ	y�B;d�6i�Dno|�_DIv^ɛk@C�*U�'5Tϙ�x+ �s=���g�������K����O��9����[�.��2UQI�����)6��l(�|��ؗ���=��߽�P�,�F���B\�	���kP4�[p� jؓ8��'�*w��L�b"�l�����Е�'(dR�����%qD��k�_G~��3g�h�W�J�{A�Qt�($�ٮՌ%�����oV�cjҦ�x^��z~~�\�n	��𑹴�n�l�>6d��U��������|l3�fLX�bhO�݆�%S��_��T/Ot�)Οh�Q��j��Q ���Ǟ���x�H'���Dakt��2�=�����h�4�X��S� � PbS)�~7�V�eg�dj(����e���"ڸ4
��_ܚX#A�����,�~���� [��\7��W~�������T��k��hn���|���?=�%C6����� �=�X�|��q��>��M����X)U����~�� �0�~=� "�Pa��?%Hڐx0�9�U���\L��g)��_�n���o�I?p����!p��b.i,� l�na����	xV?��[<Q`x�ݹ] f~C?i�@2��`q"�qh� �U�b�S�k�+��sp�I�L1��u_��Iy8f��-r�K\�?>��U�4�� ?��G�K?�ivJŕ�M
;��M��31qGj�e�#�����|aS�"�����ڼ�2GL廐y���A�a|��	�@����M#ƣw�W�1����� �
�W�K�'�Znί�R(Li$�z@0�-�W�ze�'uP>�~ǜ�.إ��dD��D�ΘT����i�E�Y�W�2H��7��p�sh�&�
>ȸ��M=2yKƝ�A���w(�`��%n/9���bt�����ɯ9f��80��j���1@�?1��&X-�+l�q,�2�-���+"�]Ͳ���.*�#�P\��L����E1D�tgf��9�4��@��k��ݍ���K��D�$�z��{9�l8H�b�V"ɊW՟�xG���.�'wE��ܩ���9��Mh� 8�*��k����j��Cm�ʚ�q�n5���싡;�9q�<dz>k�gV�Bbs��c�Y1V�/���5��&���q�Prф��O�dH��h�;_Λ#ɱ�38�!����x0��+I���[Ji�`6��7^F�?P����J� �����՘�O#?�u(�������|[!������������·L�Mira�$>99R�&���[�[_s�F[ؾ 
_��k�����E�t��:��k�w�T���e�G?坡aP�a%�M�&Z7
�8�f�θ��
?-����\h��Z�s��(�Y��th���Ŋ]���Q+WM�[�f�͊Oעpq��%:d��r	6�8�qb�ED�,��8G׷�h�'��R����v��_���r��$����հ:�� Nr�/���w�3n��ބ��Wl�c��࿫6��봌��2��,�q[8Xnc�8�Z�m&�;���C)��@8'k�J��g/va�BT1�Hd^�{Є����]��2)
��f���(=}.T�=t.-a�kLCe����[dhM�]xh�e���0x`,���5���W�
?����$f�HOU�\$We�v�U��CSB�8���0m�r��{ �����A�+Ø	��ƅc?Sn���CD�']�1���uHe!��j43���e ��Mj
��aRu���ܹ��2咡6!�Y��a45����α>b4�ݔfCsT(�z���oj�kh��)��/PGo�XAh05�}�E+��`=�XEٺ,�`��!����A�4��U���#Η^��xY�9U��J�t@���O�ݹՠ�Fh���Y�!K�^�6�����p���i�Lv�Š��B�C� �H�u�;�P$`�����"n��	$���x�>�}+�b�6��^VJˁ���P;�g\�ʡFëQ[�h	�iNx�|e+R�]��mNxoĭ���o� ���.�ܕf��&��X��+����V�3 �p�Aˈ���>W������6Liy��Hpl���PE�%]]۵� �c��9��G��M����9c�ȶďio���-��dK�N%���� A��F�gc6�mT?��[��n)�ob�c$՝�EX���6���dm���0��m� ���'�&ML�@j�Vm.n���-����a���ȪW���8���� -Ed'��z��b�{Z�e�P���t�^*qC�]T���%y�˽5�!Ǿ_��.�b�XG��B�5�4�)�,d!�' �[�+F�v(�7�I��,1Z��%�	,8v �<���V#��]wo�op���"v�x���V@W�t�D��}���!����o�2r���璉����T{�ʓ���L�A�haNlt�B�j�ծ����k���b��=Vgr�E�~�\���F�z�%i�+pȴ��I66졳���%g4v�� ˪�h$&�BE �d���q����m�S4{ƿ��]���#�8�C��w*�(��8���6�B7�YnY�P+����ad�nȘ-g� �#B�$߼�`ep��}�G��
x9��kƳ���KQ�����K�b�_�w����{v��Zn��V�qx��4j`���겈G7K8�TS0�~HiHŪí�����鲱� ����)�Jx��������v�jƋ�c¢��	o#
0P����h��jSZ��R��aZ<�ʜcռ��P�����Ֆz��A饺d��5���ܸ�J�0�~��g����u�a9������HJ� `^@	��}� o�(�|dTNL�)+���"@:�����|e��D��1�2]�}���������0��/��w���E��--$IS����܇�68�96<�Yr��q�����W�6�VƏ�=�"6|
���r�l 7��EA�̵��Q�Ϸ�����h�!V�����%|����;�k�n��;pl��!>i]�����^���R��,2!<����\�ˮ|�O}C8���;ݼ��d�2>��C���k�vHg�IO��'���R���9�RVԌOg�H#�Xnl*�t8:~���}��Z��I�>9�. ��0��m �;���N��)_ c����T�L �|_WN	�
�TCp�>[�����a2��敖��`�oZP��U��2���3��nB�l��/åL>d"���;��SO���d>L��{O�WF0�p��*jA՘#��*���5ټ�3vl�����Ux-5�`�Oga�_�tF!��i(:�>����q�� ���9�Y��{�Ug��<t�[��&�����w5�?
z�>�^�QRKՅ��Ck��܎z拙�I�UR���T�����\�-̹������<�uG�6Z�6�n���e�L�kO���r.������҂"�j(9HS?H�X!,i�Dgz��g����m+'��J�"�q����C]�?n��G4ׯ����3O�L)��U�U� �O����,NԴt�g|U��_.��2*����,����Ջq�7S��S"���m۷�����@G��X�>��)������D�2 _�tX T�����K�d�GC�al�mYA�R��U��:Guծn�a�dط�����|	��@�E��w�qª�<pVW��ݽ�LJ�W�4�T4�i>A�[9P��K�U�w'�y����?��Q��V�q/�2!N7�~� q'w���T�^�/�`���s�_}_����yƋw��%Wl.q�W�X�֙%u��94�*�s�P庋����~���/i���E�V����c�W XF�&x�_Q��z|
b�<D�SĞ�!~͵�|�X7w�Mz��~q�t��mO����u#�$K��)�83��lsIsM��������N`/%ne�Ҩ�� ��g�����iϩ��s���O"� ]Jlp��m�!m;�U�|S��=s�`�!l޼��{�NI[�����woCS��`�L��w���f��R�zz=�LȖ��Bӕ��UF\��O���2I����k� R�!M͎ƞ_-�o�p/9�^j;p+a�YZoh�K������<P�������oK:�����S+T�`�R�"�)���"�dl������e�9� �w$��G�i���.T)�%^v�yܦ��:e�Y�I�@
G�t$"���O&U�ρA��5W��������Ý�`�ώ�!������&�+��e�,�f�~@U���h
���؃�3�>���A�(���3)�"��o�X�9�d�����"��A�w�x�V'K<���X��l8���'��m��|!��=V�8'G7���u�����q�L�!�:��r��Lz�B\J�6��/S��{O9�Kv�a|��V��t0D�� )e�W!�kz.�ks���NB-��nL?���3�*:�B;Q��*'ȍa��S����ڂz�sS��������{-���
 ���K�P�}{�Q��U9���i� �V'��g�t:���3��9y�݈�
W���e�JY�VY�t�`U)V(�&�ec��|;�BO#���� 'f��v�B�i��Q����+}�YZ�
0���~i{���`�[��r��ZV��P�f�j�>�W���8+�0��ҁ=h�:�aY�\mx$0�%��U��fs����ۢ>4��Ɨp��B�]!�ِ�J��G��!��\T|Y��xm��X�L _!���&��3l['������S����}��?åڙ	���b���'�2��*��P
 R"ô�-�x�(V7tt�K5#���+_%�>�8����2��cg]	$�b@�
�g�ou&��W�M�����̯��W2ij�(q�'�"��,��uy�gn0tD��4S8�v�Gs`񊔄*��/���$Wc��*k��8�������r�D����2Vr����C�R_�	�e�\7&��W ů���I��n���B�!�a1~�)d�_���\>�7��"��Ѓŭ8���u����akެT�+8rC�CT�Ψ����Co*���y���4x����i��ߩH3Il�1�E�B߽�w�5�f_ڕ}u���,`,&���^�!�|�N�x�n�_���[|!y+d&g��`v���D �.B�֛�i?v������a�͠����M"����TZp@6��ڦ�ٗ��^J�a%�ӡ��s)Lr�T�;����Ic�)$;~>Ę	��_���`��$�E�x�dm���'�N��[�В�0v2�;��X��5x�8�i~���ث%��%�3꫅(L�����<�1��cP���e�I�����Y�7/u;NJ�� )�ߚGhT�P�R,���;>��( a�:ĔڹS���n�4����XB2���{��h�?,���M3>�	Z���<��@�C�\i�������H��}%#5[t��$`���l�^E`qV�	Cv��k@o�H�m�Wt#�뉏�;�9����U�Y�\қ���Y8׾L7~�c9��U�Ӆ57�!Rn���c���c%	�9�c�DX�Ŀ'��T��P�|E����U^�A��:�+��ӱ�*;�џ�uO�WAς���� ����w^�z��范��K�T���CC���^<��[c��>��T�k@p�,։���2ǝ��Wƈ�h��4�@�	�^�]��r	���e��KW������"��2�M���R����]�~A�#�(�V�������,=�L1��/���(�����s�n��i��6�	�|-�?�3������g��X��.+Le��;�ɜR�ڡ*L�73���~B���Ƚz�ɳ]��s�9��'!���@�F4�bp����������ZA�C*�g&'��(�~"a3�ͻ3� ��떥��l�'��Hy�e�9|�`�3r�Yi�˚��?�� (�iD�bi�Vlfm�Q��i�.�FzJGȼٚ�F��^��C���k�srW��W֧g%^p�o�*�-�n3H!���)͙��}����A���^T��S ��ԉJ��(@�$�=r$l� ���xj>O���"��M�1b�P�%�t�0�~��D����̋"=l�ہ��2�x1�bOK����L����[n|L+�z��ϐ4N+%���Sr�u����\ZrcDg7ϓku{���"[0Z-'�
��ݐR��>�������[�)�
brm��;�ӄbɸ�'����7Q��7�۔уp�S�xB����󄺌N�����(��K��S�T�z�K���]ώ'.�ad7:|���x�AA��酧��U�B��|������*�rǒ�:8�F�)���ը%�(���1��m'0��+��Bb���@���)`��?�W�z�"�E�Uo��˥���y\�<�t�R)�_��B��Znvӓ��Ԁ�:���pǥ��{����.�5�K��p�#�X,4����8�-�*,�a��Bh}K���ݛ�T~��N�E�>� �:V 5�>��[y����o+�b����*�6w�P/�v�Y�+��L��3�KU������^����6r|-
��d8��B^�7`�� �[GTNG�5�_u��:
̔���+`�jm	��b{4/7�۝O��A�ؠC�<~�r��Ñ(W%L*D�WO�]�Yl�x��<]�!��1�%>��[�����Q�)�����u���M�[�]v�+�2�!E1ֈ0\�N~cX>�Q ��Ӛ=I�zUwku��K}*#j���ɵ.3��J:,�O���w���2;�,Kbf�ɯt6�|��u�u(��I�쯄�S�bVL�"��Vל�.7�D>�A�ڐ
�B3Β�k�U��k��q��u���O��YS��g�َ��xB�h9��@�F�����TxT�I�bi�[��*��A3?T"��T��.�?"b&��Qn�f&(�ږn
�9�T��7�(�8�c"0`Լ�Q��?2����oRe똂G�YLX�E��־_�C�bN#�#�v��|yl.a=�$�a䶝ƕ���γ]A�A��2��i��!A��~k%��~K�Q�٨�% ���Rع�KHP��͈���� 5�;'�^k6U�["qSɢC�m�<�~�Q�Y�,�}��q~Z�] �*V��!�Q��Í*�to�䑺O@��>�O��<Mv�y�.<�����^�y8�z���VU���/�H�z�<a�?�ܫ#c�@��G_K�2��%:5PL!<`L}�a�pX����a��<ȧr��sf���'���~��3+�}t+���t�7��L`G��hP�ّ\�_�� �&��t��w�m��=�~1fi��)7S����T)Y�F���ʒ3�NԳch��x�ŕ�oT������-P�y�4/1T;��2�s@vxAT��Pc�`mJ)JL��(y��|z�(�׏0뱚�5-�� ?9��L)��r�j�@g��l�%?�'�L���o��3%	��z<,���od�A0˲�.�ohn��F��̔�~2`�Q���:J�0v?=�juC��p)�n"^��҉��vF<��-�*=�Pf	k?j��pe��2v�k��2t<���IbSZ�Y��˰�U2U�������EV/a��H��^^;��J�F�N��q��*=�nᝠ�`j��6�{cF�4 b4�Ԃ��_BP��¾j(1�5�*��'����i��뎺JQ2�~<�5�3 �I�k��A��D�/�/)�2��q���(0A�v�N������8G7�N���x{5.�:� ��&��I��I��y��*8����vF��+4?Ҥv��� ���q�����C��rO�G*u���O'I�L+mW%k@p�[��Mam��+)�VVy��k+���}g�"���M���������A�eEStnG�%8���6����G��$6ـ@�Ͷ�ǚ|�*ʉFv'�o�G(��ϵr�]fr��Z��sl	~g4���������fT�u�ͼ�g���b�0+�y�>��y�� ^��X�2��$<����.w�����VO������w���>�����|��6ɤ�9���5�噳ȟ�@Y<�J�*��2�/�'^�f �O���8��1,B췝�'z����a�CT4�6h��W	�k��3�<4m��8'��[F�!? ӈu�Q���������+{L�*��V�qԹ��t֪C���]\�=W)� �&=��3�:���x"�l�O-�49�g��� 9�'Ě��?���(�p���jG�6�Al��Q��fk�n��J߫����#��T���85#�G�Ws�^���I'��R��ߕte��Y����/\ϴ���/~dKї�kGdX��(rY�f�j�<�"���
�(���:1��ۘ�TK��{����j��5AB�-c���[����R#%n��=J@^��y�O����[���ɓ�t#7��A��ĬB$k��>�4�ttX���U6���\d�=,c@" q	D���3嬮({EO�����Q-����U�P@<���"�UvDs���������u(��{�jl
܀X+�=���uU!Elq(��6��L�',�7�ŴHJ�a�c
�5Oa���%�x�"B�]T�|yj�+�l�&��*gՠZfױoa�[���{��졖�[���j��J�{�E |e>�W��:�Iֿ#�����{8�E�${�@Д����_K#'/����4l��t_-��e���uOK�vG����n<����9F�T�9o�oN�zaB�A��#����ʼ&>��t�����2�Hm�`�
�d���@{�x� ���7M۱YhQvL����Bm_J��I�! ӹ�ц�Ӷ���x�.Bg%�HG:ݣ!���]�s�E"�]`u�u��2���rML'�bv����"�%�y�15p�9���EL�,2u�"��|�bYc����/�f���S ]�q�1ׁ2��"�c�t��@)�!�i�S�@�D�"��ƅ��~�	%]Y��K,�[��1�c'������#A��Qܒ��6j�n�@�'+.�5���4� H�-�jPF��[�򕈟��W��D,��!�T�?�R=R�M׭xm$�7r:�r<]�����N%=��`�<Cq���B�]�:�-�9��BSU� ��<O��3��KZ� ���tv�d�.��#������,���
1d�[��u���*�9����ﭞ?��I�о����z琧�	ߵ4<*�M�[i�X��,E�g�|$\��*���+�	�AKQ!4���y���#�q��'��u�� 0kW`r���� ���'	~Uq��c0j	��P�ѭ�I.�-���o����5���V��� Nh���p�{�o-��� �8n��>'鬽�<dۊY")����f���t�P��%��Y��CӚ���|m�(A(��U�S��'��[������}��P�7�a�b>�o�Q�B�,n9�T�{Cvs��o����IW��r>l����~�o���h�4���Z�M\�$�CV��L����X�$���7}(��$���u;�]���F�l���'StZB��:1�d��_�!{�a�0�S�<�uOI��E�����k��O �M;��z|TZ�+�6��2!ʼ*��6��L!�ɪ�Նlx̅�b�� �I���L����;�@��(}����:6�At֚h���s��cs:M�0-����/�v*�G���S��Ӿ:���tF�2�<�9�����=%�3�{Y�O�!�PC2C'�00�=�k��a6�<�+�yPk.X�^�Z���e��Nծ���=P��N����?oM:[V������)��<��iƱ�\,���eV��fC�	|�
���E��^��qCGp	|�������K���8�(�
	mT�'1�t��ܾ���29�ߵ8�ĝ2�q���jg �bܪ��P{7��A�\|J�����b�,�6��b1O��
[�=֖"�\���&�3=��-=&,�"b=�5�ؘs��A��i����}X81;��&�����9y@�����w�d.�p�\h\8x�'Q�	<-�ȧiS���-�V�C1��__@�c3����[;R�;��/�S���%��\�r�#Ql�ӳ����4O1�3�_�5?����s�Ab���p�V6���q��J� �nqjN0�_V�-,�v�"�ݜц{��?�����A!t�+V9��I��%Efy�����t8\c�_�8�tR\���fG���z��ȑ��i6�7�?<}$��a��}b(Y���dv�����"�y�-��?���̠�j��r ��e����p�~� 0����w��&-�Ci"�����&�^��8��J������*}n�)�!�'���+�
9΁�jǈ��:/����|�|��G�c�&����TH��f�\��1�Z	��K}wa|<|q4�l�s�b�w�o�G՞5q�Ẇ�WBH�#�ߛ['�I1�B5�ee�	*ћ��3r���6!)�]K�9��5��l	
Y�;l}7������C�}1��=�JA��wx��Rp��=K/W�$J����0�8��&���Z�Ė��UD���oL��Ǌ�Zp��ӕk��p�@�'\�J]�%�gf�������e${X��s�ڢ|�;�A���ZQ'S�����p΢w�6�_�~]�A$�${<>N�L�L����n���D�)8mp�G�$�����4֕Q{��]�·(��CQ-3�����\~F%?�K��(y�OQ;���\�3_:�&��p@�-�\+&�/��B::yr�g}�n��ە��o�:�Gh���q,�'G�m2<4fvb&J�x(�v+�gn�71��g(e�h�r��蒷P����+Gv�5�����:�l %���m�I�5��S�u� (]�W?";,��Y♟��&�y2�8���9r�z6z�����ڎ�U.��]���|��"kYP�����N{,�G�Hy�2(3�0mC��<&8!�rff8�2B�Z�zS��ܽo�g%�f�p`�.Cf�T7�_���	H���*1��;��}zg̛ۡ�hV?�>����ǜ�[�VKH�9�:U
�(mW.Y�%��:�'{�m$m��&�z�h���[X�����o]��ͭUkk�f^�
�������Zf+�S�
�bc]PWZ�L��H�_���|0W��jt��3t�̸��?M�U�aj`u����lѵ%��EG�.]q���"t�k<{1�:��z��e����
��5#�%;���8�] �Z��,�(��P��R�40j����qoV�y*C��[QW�l���Y #͂��S�|E��S�T2�xt�h�T��ͺF�#N�Q���ٚ�)4	Վ�#��\D1Q�ON**5t����~JK������#џ����}�mP��5#�l\[d�us��k�^�'Z�Ͷ���R�~��NxGº�� ����He
3ϣ��s�� 	���H�O��:�	b�2����/����Ƭ&��}��[ٯ�Bڿ�$�$���D��#���1 <�v�b���S��;�D���?��i/(��!'�A��!�}�P̚���X�N�����*.7d&?t�t�S*ǘG	<���]������v��Τ���7@bg�{7�Hl,�|u�����i~"d*]T��T�M ɣO%kP�C�n�3po���/a3�*O��gL�d�[�o(��R-/�ws��}�U��m3�Md�q�������}�5P�=��Wa"��9�i�G ���q�&����9y]I������Q��[E��;��sȴw���γ��s��#촲�)���=$�"��>���v!&��h���,ߏ�f/Y�n<�ZW���NY�+�O~+�RR~���df}m��B��pi�)���4{�O���k��{O���f��rU��Fg��o�W���5�6�>�a�}�^":�s�ɌG�@�&�f\��m̈t)!��4�j���tj('�!_O�{�W`��.j��K<�WL� �a`f� B��3�f�gN�3��9�s7Q���Q����s/;H6_Z���}j�G��`ߤ�H<�!%V-��̾��GP�Ѣ�-�n���}o#Kz|�0
�מ�'�f6���ׁ#/���I>��m�/3WX�d0�c���G§!&V�]պ�������՛`ޮ�u������_+3�ZML��l�XڈlO%pN3��ً�w[M�ӵ��!b��Wl� �b�N�(�
j����� &�scZ~j�����-ላ5=�G5��;]�T��'�F���:��}-�ݘ�U�3������{N rb�_)�O�u�����1�C6W��?a�HqJ��d*�^�*��oӾ��;����;�Ii��ھ��x�j#�����]�y�rW�H��0�����aH�g�M�mi-��)�0���+�*����� ��'r" �#
g��gt�Bn^��A����յ���kD`�n��q9����P,����<�I������/%��UO�fd��.:��Qh��k}�QNu-�lqq'c�F�$����.����4����̵c�����,/�vz�k�5z6�m_��VY �im��WW����r2��D��u�ʪ�:W���6-��Vv��$XAE�M�=�GO7' �dw�"�Z#����:S�x�}���R���ǈ�ӥ���>&�����j��%��qoy��N�I�8�#K-��Y�b��˧<b�P�gYod6fq��`�k�R��:ä�
��/л<(O��u�2�>k��UC@���b�*��<�)��|X&����z:�"�X�\�aBP��)ޟL��c��D�)2���k�bL��ђY��~�6�E�G�p�t�b� ���*��$E$i�v���r�N�ex�.���&����
�0���_ww�|x���ϣ5�Ej�t�����(Zjr��KQ������"1j��/!���|��a�D��:X���N�nE�042�蜝���ު6l1����m=~�����E�0Y>h��%��x�F�k𧭍0W�oLգ��T�1��__�Eɟ��̡l��y���au�x��{����zaM��[�.�չ�4�E�dr���ZP�D�aB���TJh�u�u��%���b'�.��+N.���&u��b��>8�D	�$ߜ�4lq/A�Bn�� �����!6*:��+M0Z&rp�k�R ���t�?#X���,���0��FW����1�.��J/�{���[ڹZm�N�$ ��c(��`�ԃZ�	ZC*J-�\�����F�K��xͥ*��� ��Ν���1���~�{�>Y�=����n�"4fV���E��Ae�m�~=M�9;7d��(n�9��N*����`��1ۑQn�\�����#)������+���5����mW��}�XdE�B�������l�CDrӨ����m%�&��`t���t�K�f�5�/\�wt)�$�:?T2z�tTa�{������'��-�nR��.8�v���^���9É:s���qUY� j�ꚫ�	)h������mЁc�[�+��z���ѻ<� ��Dj�C'Vq�>s)��5�9�k��6[�P�@��^"Q�����{�կ���Ez���Sb�R�pwl1�(ф�A4&��I��=�t��!�ʷN	��"1����#����������N�΄{ɯ����^�kX ��{��딧��U�|^�V��D�����ԨB��,ܳ�m�v+w�E$�����m�;���jM���ra"��'����l�|��^ )N�)��L�?�b<0h-�7<��4�����~u�ڧ���^5����QrY�����*K��9sc�ۜh^@}K+���c�F����6�AEe��R�er�l!�����/i��V���^%��0�
֢Ҕ��W����a�-�꺫�h>�~�46���ҠPnwH��PŮ�j!S�X� ���Vt��O�<��vD�3�3� ����>u˱+����\īwP�2����}��з��+�W� �m0���聭r��VSa�'��%<>gԹ<��;���[��:E��o�X��B���Y/v��/�ã�F��	��'k��<�?x���\:yS!E~�&�`��ca���A�$+��IC9w3��d��n��Q��m���Y���'Xa��w�qK�f��xN���ѯ�v�'=ґ�D��:[�aj�(�����d�q�H�}qu#HiԷ'�5���pR)[3ʷ��^b#\	����n��,G�M��ϳ72��l�5��_������^�w�'�ie>Pģ��vv�B���X���C�!�F���#�o�2�D�攧P	��ϒ��*'�r���C��L[�������3
��@�^	sImr���봼��L�ֆ���TL,�Jo������w\��z��{�N��˱�U�o�3��,�N��H��b��#��3K��DW�#�=Bٖk<�l����p�V�J��޾��!�C�̦ D�"��<�Ӗ�c�9MN�@��TU
��/��Nڳ:�S4B�? �="�%l;~�k�^�-y��a����Q'iM�|�L�5*��$�h���
2���&UB��e�,��s���0�� ��cW.P^9O��P�Ƭ��H����د*��6$��`�Ƴ`�sŴ�lNq���I r�';���V��譺�Q����t"0���+.�"�ꥋ�N%Ċ7�mׇ��*4Zt�l�«�e �3��i��-c��9�A�c�灥�cj�Du�nͯF��y'.)���|msw4R�0��X��̳6���m���YqOU�mq��XT�J���Buj6�v7�f��� ��� }q�H�ՉDIQ��mS��I��ͬ-���РaW�P�4m��~!��B�S�4^��3�Y��L��ػ�_��}�&�YR���D�c�Oа
��x�@e5�.h�3��ލg4�Ɋ�dO�#`�,�����E�����^,����1��+(	
��L����-Uu�X�S�¦ �ᕗ'ce��IMW:�j���n�����묞�v�	c����2��Q�"oñ���N�m�hp�$�7���s}<P��k�'��S�*>O���d�+�n����6\�J��T��qU�a�Y�:����=&H��1>���h�2�+�֐D���bqM�V���������>8i���cv0��B����m��"�A�q.��g��b>&����x7K ��_F?(/��2�تh4ޠ�g�E�_�ʌ��"��t���Ɵ.�<c�[�\4�� =i#i�nT�Qy/j�-�B��W+JY�4��-�������#�/�ϵ��D=��7��L1p@ޏ~_�lYď�ޞ��'hz�gP�{߆*;�[X�M(}���sC-B0�0�����'�n��ӗ�AE��U�F5�Vh/v�A�*#�i��K�/�76�v>�ʺ�w�:�.ƀ��+2J�g]<}^I�u��2ڲ ����^a�yG�uQ�i�ǈ�ro��Z�Y!���Hx �W�਀i�
�)-ީݮ^T XX�F�v��($��c����ƛ��7�w�$�*��6T�� �\��sP`��~'V�v���<Y{y��B��>��>pvX�!AqM�xU�<*���D������j��*���B�n7���E�s|n��T��-�g����$�\{�K��
I�j}$�I�����I*�@���������	i�\@<M���ET��_ۈ;�p�w bkk���,�{�`�� �(��]�A5U���k�U�K��N8�t��l�L|��&*n��i�[o��a���'V��?9�����M6���z�;j(N13�O
bT3M[�i�#�Y3�1��:0r=�w��\�J�,%�Q���v4�F=��ψ��D��~�E�4hC�1�_���c�_�M���(�JUz�w�+B����J�C�\���m��A3��<�������Vq ��_�W�E$�d��t��Sb�3y�r� ��+�kI��_81��{���3�05�J>6���7������3� *��	�H���։���KG�����c��3���2\ͽ��|�f/��7b���n��+�� �Q��G?uŽ��k����=1f�m��,3��!�Q0�T�&���?����?~nt&���=	���Xޢ	�f����:'�1{h]xu���d	�6)��1+���F[��@��/%�	f���@�0��%l��~fi���[��_�����Љc]:!t'�-�����"XXXVb���߯|T�d׊W��I��� >�ˢ�W-Ё��d��6-\�\{�s�L5hd���с4z��c��ߦ��K0+������.���Z��&j.I���:�&�[e3z/g���R���!7Nn�~gミ.=y׭>C���z�J���ڃ�=5��9�biM����� f�V�ۢ%��85	�ʨO���9\y�i���z)��K��<61�T�y�gex1Q�E�o@��β��\m�2c+a�;�QP1?wg0C�B�%�cJ]>�F�e���c�I2�"���G�1h�?bĺ�M.N'�U��cɘ�&b��=�s��3V�Ū�m,�@L���1���E3�zK����f�+�� K���>���6��II�Ò,֕m"�p���;n�����&+.@�`(�:=w���{��\�X����'�ų&�a�T͚�y��f'�]�L����5#ۦ�Ԧ	�X��b
7����+$6A���0^��C�;5h�:�I��<�K�nJ����I�i���/��6�"/IWW��N(Ya3�-�y[�N6�Wc�Մ��m$�u6��"[��qZ�c ��'��t�^��s,�q��֊c~7g�˨	>��"9%����泮Ou�BT?���R�֠N�1�)vF�#���	��&#�@��%:�뷚c2&"��a�R������,!�[LN�Z�yS� t�Iˎyo���&D�m��_pU~"�	+��6ل��p�PY�Ԙ*�y���Q_͇ O�)ܑ�\��i�E�%����b;�x�o��9��٧f�C������[r`r�c`}��u��*ˮ�z��zB��3��=�#�_��ϼ��hg}���p���,ė��<�6�2s�
W$�X�Գ/]g\%�s�M��H��DM�e`��y�1oH$��qB/��p?��Mp+�Y�`TI�g��b�6E����+1K��h��&��ו�UG&ǟ�y� W�D�q�h0sA�ֿAVN�T'�18�M��>t������M��g��D���]�=���f|R�p�`��h�>Z��b&X|<?>X�5���2e6#��O,��-�`:I�0p���~�n"QI����Z��ɜ�D��|�,ȵ�� ���K����BcH\�F�W>�>���W�U�.�r���䰩��;��BE��𽔛#��=]:���N�6I+BZ���y�^�[d
�h_��e���$ʉe�^���(u� ϒ���ŀ}�d�Nyr�vҴNS�-!��@���7����k��y*p��q���m�Ք�gௌM�7"B<�07��$��**�e�gk�Ѕ�Z˛,��K��	<�KͲ���a�p���9"��+�Cr9Y̜�hT�s׆�c!��gTO����/������Jڮ�.�B�ϵ]�OW �����<�����#!��T��$Z:�P���[`�����>�5:�q��4|�ڛ۝='t��|h~�f^��@(8Nw�E�RˤV�6~܆֭5�s���S��,���3Á0A���9Ed��ֿs��m��"���@:�h�]���(h*R�J.� 7�xZ�x�Z(�L��%hV��aMq6jy)�'���V�nA�H5.����������n'XV�i�#��j6�ע���X�� �pc�X!�Kh�f�
�����@ m��e�mP��T�(���0K�wzr�D�:��Xݹ�KG��湁��`���H��`���\_p
,8s�ѳ�y�Ww�7��5ׯL�P���@�3�e���ce�:�#���Oh�4.���|��c�ɕ�ꚷ�nV˝�YB�=�y=�k}W�}狨�p3��;)��^���H�u�z�ݺQ�-G���%.��_���� �Ni���A���7·p!���9�2)�~΋�Q�ˠ����-3>������i�����/��'3$��@��:l%�O�s�i�wS�Z}!:�#7��ﯵ�]o� �Mˊ���W$ܹ*���,k|w��1zk����_jvpԫ���y2���(e��bk.�ȫ���Z��&t��*�{W~�	EQB��W�=j���d��0�=bg��"�U��)M*K����(x�?�Q����Ѥ��6��m�y� ��ʎ����G���Ϫ��.���r�?�΀�\��G_��
/�j�Z[=(�nza��DD��������XA|(m��W݃Y����psZXB$zt>D��.� ��ڊ9�w+O3d�t��� ԶW�������&/�	��o�]$��Z�@^7M�b���������\~a�mI�*�K���
�p|�+���u�j��:Px�W�-���� %��'fI��3a���F�v���Y�]��<W�A�h9��'2S�?���]vH,���o�W�����5�b�^)�`�jG��B�Ͷ�s�����e҉�VM���5�*@�����ڈ�����DS�m+���mUX���_`�Tw���v]7�d5�6�?"x��h�e��a�^��t��"|����^�_�m}_-�TҌ���,p��M�AӁ��ڝ�DcR�%Z�����l���� ���Mwy!xВ_�Q�^�p��$�e���Y:h>�2�p:E�LE���}�(Ƈ�x ��j.r�����u%�RY���%�����HY��,��	�ڤ����� �g�(��Q<��C�=IX�m9k��X���s�cR$X�uD�̏"��[�>��+hݫ!�ԙshI�N��V����DR�o���\O�8}:����1y�:b��uY�$��5�hʸ:�\�C��+������Q8�A����_w����� ��9
�IX���j'��u	��Ǜ��
�?�e������l�K�@�}�.���k�SJ�e��\Tr����4��$�Iw�ɜ�h�3]3�dBcu��,J�`w�g<KJ7K�(>Ŗ��lZ�����I�(�T1Zr���iӔ��tkXb���#h��J��<��E��2[0���R��It[	�9}�q��QD S���tl/rpBm�%N�R����/C�	�>�uϠ���Ƚ�"����i�û�RJc�2f�MV^�m)n�f޿���WC�@�e�rh�7���R�yr~�����Y��(�������=���oy�axn�7��s9'��n�,��ZYL\%���hB�Hj*��M,#(��6P��jVT�F���'d8t�?����:,���ɻ~�}����{�R�o7��8�Ɍc(BG1_Bq�����?$����+�Q��P��!����7Q]0ɑn���\Ov�I�����E&���W�N��(���O��W��F�@ʑ�#��BZ�鑁2<YF�(��W�����M[	�|��y�� �Q�����	:=�[Pb���i�� ��[�*�Rlf#@�:���^��U�J��rw�D2�4E�}�+ZK�n����>����;^/ c,�!�
CQ�����Ɗ���>�A�lIS��/����}1�H�CF��`�����qjy!<3�lT�8j
�Ɖ
�:�R���2˻چo��j�yV�W�ݤ�n��:�I[�����0���Ơ'��F��HlY�m�x���c��p�dy�O����]��oZY�$f$��F��+'�d"r��YR9���Xt"� ���@�����D��u�V���OQC��M�D��=�ݓ�#ȅ��ۗ�	MM|@�j�p��'S�}�������QM���D2����;��APV����m�1{2d��0 9��B�M`y�A��p%�ID�8��>�mW+��ݾJr_:V� 3<��%�w�~�fJ�l;&� P?.���5��a9�h����&�VsB�-�{�B�׋���pG)1z���Ru�}�/�ڪ�*P����`Q�^��hV�]�#��v���F)�+��
�� ��Iw�u֟03~������-�7:��ʕ� ��v�|�W�Ӓ�����R�n�鏰&�0+�Q�σ�ƨw�IK���� ��/`�l�ٽy���l8TS�O�
���iٞ2�w��Jx� <�����e�`���ϴ1��/�y4���k"��75��']��:�)z�c��o����B�>���3t�ߴ�1q:L�"��˗AY:��_�$�3Z��"�i	��vk�Y��Z�-&_Ou�������m�d{y&'��z��&�~p|��gQ֧�L�tگ��c�����?�h08����؅�Xɤ��0�Z�@�4b+�~�cM�1Te-I�}{�f�p02�bˣ��\���Cа������~?:+�:�D�n�<��Iq�������E9�N���0ԙ��9w>�u{�*���)��o����4��h�C��S�^d�Z$9v^�Ã�٥�=��]�P`dv���R��xZ[�>K䄔$)��<R������ڡ������~'t�b�[`��K�D0>t�I�7�6o�2[U�`A�ə�ꎐ]�/"R��ä�����7y�U��,�NgVTm��g� ���Mu"W�fBtL��o��V3�[��Jƶ�?&�񜰰%A�\6ٔȘV�~ˣe�C�<6C(!���lG��Ϋ%_̑1��F����8�_����z���'ƣ]�ǳ篲�k��X/o&п@/|��g��L�����튳F��&�:ث��#�D��㮛�9Լ{%����3���Q

�Ǫ�Fe{w���4��.�?eUQ�坊�/v*a6�M�a��a͉_R���;��d���]Ѷ^�`VV��>z����@O�Q)��T�QS޳rF�:��b:� I�u��'��|��G+.��s\�F��f&�ɛ�zTB�<QWt���V��	'��^�]�\@�j5�?n
◾�̫���7�/�ђ�B�'w����Qn7}�� ���D 
J�jt�q���>{�I0觾�&�MW<�L7k--�t�*��'mk��R_9(�֦�RIV�k!@Z�>h�U(�DP��9t�8�M�r��J����M���^�7S���7��T�T���Q�4��1ӵB������͞LT�H����{�{$�Y\"�8��L;0x�w���hO����ayݡ�C��]������n�	0"ev\�H�8�*F�x ��N�-P�$ <�!��soY��@�t
��f���`a�m~ݝ�QQi��7�U�k�V��nr@��e<]�0wkf��8����@��%}�׭U�+�ڡ.N���.�^e�e�B] '��x�=��r4��ǉ�o�����W��d������-]NH[E0�	�%���8 �9�h�Pg�5��jC�/��9�G8)��>4SV�����о�ۮ����:$��A4MdKv��t���V~t$?8h3�K�P���Z�Sf�ړK'��I��A��X���N��BiT�`+���g�������BN����惴��6��~���`��ߎ��ZA�'E/#/�k�E�����Ϛ�7";�3~bro
���&�3�u�:�M=��O�<��ǒ|�*I��e�/�qr��1Rn��&�'��[��ᨧj��y��|��v8�)�cK���s�MT�=��qt��T�l|T��[��Z|�5��G�Y��H���|/&*������gY��b*=y(V$zr5�b�nWqO���d��i�V8�0|��Ԏ�*Qo3;t[�I�b�M��<�w-)�3������8y�	a����
�x�AK�	���?���{+#;yRAC���R���&X)7���B���T�IWp��_F�z��� �:��;l����&C5��Ԅ�����
���9�0�,C�����la�B��z U��a�ab_)��ZE�����7���ϋ��r���n�&|�@�͒�@��<��6:[��*�q)몱 �{�N��%w�HQ�L	�T�˵f�<�τ��?J"��h	�<�i��/�p�=>�E�v.P5�B�QM݌c�ߌc�5�W�$b���HE^��ش��@���7��l]��_�����3���#;�(3D7�0��2�1|�Ek��|����d�v�p&蓱�xgS����~��VY[S G����-�Z��gC��LH���y�K��ϫ�}2��G-R�tEQ���o�ˌڌN�O)Ƿ={m66l�¶
���	�=��=ga�_JP�UeL��BX�j��ȥ���Gy��h&�K���z���%���"c��En-]�2���M4:�E<�hnJ���������]>X&2�N1���/- �Y���'b77��UHء��}�n1Mۇψ54��
�	Qo����d؛� /#�\m���CFK�]�z7�����2>#캯s Vf���!+Jo�d����4"߈�w`������kQ�Z�H]�oc/<[!`�r�7�9ȁ�#'ȉ�W�7�~T��ȃ����&�BS;cR�q7� ['���mX���8BN�������
Ϲ���[
��5�b����(�9pP��>�Y�R%�B��ْ�u$0����e|w��Q����s���W+�B� {�`е�W��^���`�97�L �Uk�����\L���ԣx��D�5Eޡ;��g�X[$���Q������)Ex#l����A�;O��s��&l����·��!gC#s���a/ޯ.��S�v��ԏ��u��m�&�p�905O�h�!�$$� S8�dF���%�XISŽ1A�q,3�A�@�ã����* j��ar�zO{uٱ+�jҼ���ӄ��rY��@�Vq{w��
���$9i_��vvp�P{�I�ۍ{�Vɦ#Ki���یxiX2�(*9�!_f����p��z�Tc��6�G�K�ߎ�:��NJv"���M�@�c�SB`�l2���G-d<7����� ��� �y�'=�䨬�b���CT����!��|/&_i��"5��f��@�Hph�"���@�	&ԍ�}mЩ����e��υi�_�in���l���IW]�����d�w�A.���#�V:�����_J�D�\�𮙎8������M��8���-�x���6�z��nLE�kDy�&ǐz���མ�t�?�ߕ����*'`���<��)|���c����?������)ȁi�DX7/��33.%�|�1݈l��F���1���?��q�C8�@��5a�R�tB�����q�x�{�1�����5pn�ArY���5�1������y��)��Ѽ�`�{�����M��GL	�]�,(�'x����_9}O�.�S��<1�I���;�F������nؿ��s�݁�#��'|��G�(�`1�0q��U�f͂<�i���8:s��)m��s�nllz �AE���ك��x�����M�.��7gԸ|y�@.�rS7����̂@<�j4�q�K���73�W�t̀3,�a�Y�z|?]:�˾��8>����d�{��^M�O�t6U~��|��d�'�y!��]��+��r��3�o�5�
�g=tpt��v�L��Q�cLx*�Å�`�=����Y=�j�3��hT(U�!�}�"�x�r�s^�#L����ܫ����8��W���\ ��`c3�q�;�aᬔ|F�R�>�!���
0\&y���J�`�i�<�7�	�lS�HC�£�K�Y����79O}��e�g����G���9�I�#�n�c����[^�SI�?����-�!������x��(�2����5��������`k�]d�&��^�aV5�t"׻��,N�T2fZYac�a@)w�;��,��yV_��LQ�#����S
ƺ�`���>�W����,1P��8�ǧݺk��BRY��O�I4�z�'L8�.:�}�v���JȐ�:B]K�����"&��ʇ���/�RX3߰��\�̍���(����O5V���}D `�'��]�70���s��W��k�2���&�(E��@AKi��5�8���(�(F(ifj�9
ӃZ��ϡ��K!���O���
x��ц=zc��GB�'�k���Z:�/y���$ե��l���R� ����O�vD`G���Q������Nڈ�
z�z��f��S�྘�v���Q��T��
���HخM|d�"%C�Sb���uo��V��D��ړS;/��_B��pE\}��7AJ���V,5q���<�)6����I���YQ��P�����p|�Z��0�r3\K ʹF"'��ߴ�|h�=XsDN54V�}@��xL-���s}���I�PЫ�f�W�6�q��O�[i8��Գ+�;쟛v��N:/f�v�A0Į�*=�e3;^|�,M����D�K��!��1��'�L�'w��U�$z���[���3�{�_������s���$���qܺ<[���Z��h�+f���L��@�,M^�($4\����-�$ Պ��W!#4Ty��-�mO�r��Fë{�j��i��?������F���z�j�N>æg�����Y���bac_I�`��y�3b۱'���82�ڵ�Ia\�uH�mI�0it-ÞwFϱג�"���d0t}J�<��^�6ա>i��"��I&x�4��?�����ٖ�g�4u���b3;��o5^���9Q�����dP�&O�YP���j�uZg�T@$�r{7��
;�E
��}s�mI͘5�rK��Xp��ۛ+�c@ɰߎ}����!�7�}Xoz/˶n%��<���Ə��*,��I�)3�;�ȩ7���a�u^^��j�50����6�.���غ��\q�rHÉkUtg�7�#h�\��Y"_�IG+��u�T o�����1�˖Ąݣr���B�ZO�ϕ��M���Z�AN��y-�M)�j)���L5?��߃A�v�e��x���_�f�D	�L�uP�����>�S�4��<8�?]�i*�D�*��\B�sA����v��^֧��9�oDkP*��ߠoy�q隝wH	���I���ף$���k�  ���l!���PY�wo5E�&���aV�s심yK��a:XY� �n+�?T{7�|�!H,�y�^�8��p!5�� U�n6%?�f1A{�
Pܴ��5/�%�ۘ`����2V��i�`��!ʙ�W���^<���¤�&����n��t78�hD�TSB�`��.�y̮�U���5� ���-�y!��M�P��l�������Y�Q�Y}k�zAP�+9���
5��2����l��@>���J���nZ�V��WI`���	ͦPԤ�M!i��]鷆 �%G��S��z'���;U�N�� ²�b�jx;k��=ϗ���Hʻ�Lg.w����U���L�Z�~�Z�X�p�$S�D�aS���E�����,dE�H��[�����C!u S��qWMwZB�
��@�>jhO�c`,�M������:�!?r���S�]��u돐@�~��I�p[|��.w���#>1ѳ����77�w����*ح.`xZr-��D�(y�B�\�?�7]3û�^O����~e]9&Z&�GZ[��<m��g?p]�8#_�a�6Ǫ�����l�����ϲ�I�1�Ǵ�T���y9���)�;�Q����(�-�|
J�ML��%�����ץx��^�3��Oyq4b;Ь|�6o%��d/�E�N�s(߯�ӳ�����Q��v�Kx*���U���	ӂ��B�6�v��8ޭ���~��+:Z�82�vi� ����D�Q�2��Z4��%�g����]���J�T���	m���T:���B<�Ϊ̾�9�.�-�wy<k�S�������m��q4U�v������@Mcd(�T}�[V��1��0b6�yh�{ �$��V�G�� |��X8�ʄ!��c�s>�����w�x��]�
8 ɛ�n&�\�v�k�#��ȧ:K��.���0�f�FJk��2JĊiH'�~`���|*��v<�M�7 �⒧[�x�ނu��>�:�! �����V-����Sd�`���-5��>�R4�&�N�)���u�b���,���/"�b�x��ҋ9?DJst%Ը���sT���PgG�mԏT��H3�K���;Z�Bj2���nb�I���hݝjJ�M�/
�>�7����jC���/�ja�����Q����7�h�G~V���1@��V��~M�4Y��I��D�Lۢ�60����I�/��V��hzӗ�x{N؆�hVi�G�j��c����$�q��!�5L��tR��tO�k*Z<���	��7���^tb#��,�?wF+�a(S8���|�#=�0��g����3���F��7N����s�7@�]i���[7=�Ε������,Y]O���N�xWE��[ƾW1�ߐeu���ew�R8�̘�?ت*��[��wo#{"�6��+�����:��n�+�.|��r��{0��󝆈�[�wF�\���i+�Y�mNVV����'q�ɡ���	��֚^Z��V�.I�F���5Z�E��wQƉ����x��`g�U�݀X�l�IǵR%�2)��zC��cҗ$����������u5�Щ�����0�����᠉aUR��[g�{7ӊ�H��K����-��þ������C#H�~��:���ع�����չ��R� nJ�\�A�w�7��.�H^�6��?�U�2�3�~ԕ���9B���sx`h�^�4Co��t���S�.4�*�:��Bn��'B���ϝ�$���#M��U�hŜ��>]������}�7�e� ���_2�Ay�ލS
nR3&�(C�)9Id�Vt��S?t�[+ Y��
�,T�J{k8��8/����o�s�5}Z�g�옦�(�I@&���k �	��~��j�N��݉vD�8;��w�.F��|��	�����)��4B�$�ժ���\�������0��f�ӱ�fU�N�C�CK�#y��m5mbBƔ�K�_#�b}�$��W�	R?U^�eT�T�2˫�)��aX���K�kN��@�]��-_T<�rX֝b�"�׉�3Ϡ�3<+b�ݮ��\��YA�+'�ρ�e$4ޅm� ��ӗ���"ڙUV�g�g�U���&jg�yskB,�]�m�]�(���WF�@����w�>�l�U��m<!��8s��vF!���Jyk���GsI�����硳��*�=�Ƶ5/�:P|����1�Pi���jb��J�᎟=ũ/]���_���"#By6ph�se�C=&��:������I�E����᠎�6���L�6So=z8�t\�����Y�����<sc�y�����������z�X���2�� i@����j��5gÉh��Y��5�	 �s�M'1ib�K��;�����S�9�`+[�z�N���
0�S�Wi�f!�C��*��VLjC�Z�=�P0�up��f�L-�K��g{@�M��`�"�������8ж���!�u8����Ο���bȏ��vW�x����ؙ�A�
�_FC�k<���7HuLS΍1;�
x���k�����| �g,�ht�؞3��c6��xSc��� 0��HU4r1&��M�����*������!�|QL�^�<�3���Ђt��rȲ��4�W~����`/�0vM����.�l�oN�r�Z��@����}f(ݺ�@ɿe:޾To�����iS^ja��i�"(���P�Rq��a�Ȑ@�n���*3�N�7�|V��� Ʈ�қ�D-u,8�Ȁ�=݂�/��r�`-�3OUh�#�ą�t�sa��~Sdb���WK����?o8��G,a���K	��W!F��jbX^ �F�AK]�v�
�
�'Q�41�{e8:c�9�~���`�r+=N�5��粶��SX'=�&�Q� 3{�~�RHN���
R͎X�q�ŭ� �A�\D������,cܷ��/��:������>�#?Jug��Du	r��=_��B?$^�������n��oKѢ�4�ɪ��J������Ge�E��� ��\�ߎV��OOF6�b���KG�����N�--�'��� ��<9����U��D�U�vf�>�Esd�FHҺʉ�$�Sʤ�F�Hl-oeΏiC��)N0,}��xkz��?G.�q��߀�B���"����*��8O(�y�mVx8�j	bô1	V����M�ݫA�T�Dڠ}��������S��^�]9�rGϨ��ݱ��o2�fm���$`LwÆ�̾�*߇;u����?�.��HA8*Wg15bC�����1�T@�hE�K;.�N�AW�h�]���E�W�06��Fe%�>�k�xH��r_;��Z�?�s�`�Ȱ����'P�j�'m<�ge�P��n�jds����,��`��$��e!D����t��HX��9���=����| ��$�u���e
��V�i8�m��[�d"�侟�'}�qR��Zg�f�1�ǻ���v!��=��^��j�JH:�wk0ǝ8�pq[ #�\��ty_� `����K�b�P�5K�O�A 9�}i���b�	+?"��eja����N��<��>�����k�`&��n�(���y�S��P����և%�A,���yi�Z���[[u�23�:��9rnɅO��B-E�Y�۪�����,Z���c�b!����;��}݁�sďm�2(2 ��^�Ņ�G;馟}��@|����A�f���%�Ap�l����g��Ղ�D>���:�?/|�c�A-�8ն'��k;��/�/��E-��刬5�`#�����C!g��~�����U��wn
�Q�\�h��7�.����A~D��%�}Nɉz���12Y�:�w-�|���Y�/����m���Zup�� ��;$�Ok��\~���n����-�IC�9x�
X/|�� ���٥�$���"i{и�u��m&��Uv�d��ߍP�e��?,�"�j�L?Oi*��D�I�I4)m_5�@r�S3����Wn`�|��!��:���E��̊A�W+]ce�؛A�����v�{VĤ��/�ZEq�َ��s�� 2�ߡW�`�ώ�\.+7�d�χ'B	DS���g���,l�0�M$Ri̙"�!kH%B��l�>�C�t�e�N�Q�+����Y�o&^9[��ϮuL-��"/[�\��	%Um��Н\��v����:�4{�G���<�_r!�8���8&+o�S7/
���.L�y��.f�²r�ژ�b���#��tQ�"'���UF�k��K��Zi�:�Z�����a<!>�"�L���1H���]YO�KR6�U�ܷ�&��j���J�?�"�����ث�9��_g���o%��>C�N����)GtEo4�ҿ�&��Ul��&�s!���2���O�/{1�sk���ƃc�7���q�p
*����P8`�؉Wգ���������e3��x���YR�[c=�2��;i�L(�ޕK}�����m)R9cKXnU��� 7��ϲr)EW�R�q�<Q�n%�����RC^����½oz_�H��@���7�����v��#Sq;K|رv�U��j�(�u�]��wIk�s���e?���\|
=��&��k���
��-bӏ���~o��3Z��'rS�#s��[JB���Y{�&�ƕ$�s�o���˶��j���X�"�~F�S,p�?������S�/�2���u#�� 3�;�G��6�Aǐ|�%2�o��U{�+��6����y��{R4�'�A�>��Q�U������klaF��A������������{�ю*S�^I��K5d��9I��UKa�%׵��{��9q��.��w�4Nv7C>��y�����eH��!�"��N��݋lu\eʺ�R�ͅi�9�Rp���sz.�?7^Wn�W����&B�z|4Y=���L��^�����
�N�}(^>�CB`����� �i��<�C���dZ����@�m��{�%�x\SF0�Z��˽�~���@$6��6��A�r������;�"Y�m"6�|.b��i�^� �$����)!�Yz�����M;jӉ�H�gU���̥G��G-� ����j�b�	-�$���Ϸ~�e������T�VSĊM���-]��'mD~���?�����_��3��-�6M)]zd� �|�Yr�,lf_�T�O��j���[�ߖ���%��$U�*�J�W9<d�Q�<y����2����P.���Ta�Pݗ.����:*�7_1J�9�����0,L�� �e����������ıV��3��Ş�O-N�u�(˥n�N�k|aMt�\�HpsvJ�,�/�WQ
���T�h��bhB��yrh��i�7���'jk(��g����RO�\^B���-A������DB�,4(�	I͂��^��aB��$�w����3���
���TB*`��	�/9Tشsє=��~����� bx6g�Ü�T��Ɋ�N��+ns�哀?ʉ�*�T'��InZ񊦆~pAQ^|�+ٙ�݇v��	���Q4P=�FU�ùHgQ�/�D���Pn�	`C��	ظU�v���7%���+�2)-�2������Y�0u���	�rNhPԺ�����R�L2�����K4��k�@nX�>�	�L�x]%��Z�KW�i�JV_|b{�D�3�H5��S������lɶ��)��6���6ѭ?Hv	�5～��kXY�F1%���sz ��/����&���'���d���TB]�	c�@Oe�;B���\L]A� �;�Ν�>�P�����n�y���R�6��q�C�8,��ce/LPA8��}�P�	7����"��M�9�����i`��m�*4���-ڷ�s�]��"V�E��J��xʴ\�F�� ȌuEG�¬�[^�x5�5�[���mc��`ޟ\�� ^�
�HL���w��~y�CR6P��b���|�n��i1�[�t�&��#�x >���^@�,���Z��O���/`�@��,�izA|`����E�N��q��"�W�^G8�9�ݲ�U#J�G�a�#üWs��>~��!TX���Ic�<B�Z�x�"��x�zV��H>�W�n�dE�417lвB���y��]�����Ù,�*���J�]	K�G>{!(��W$��k�>$���mӚ�ʉ�Y:]���#J�D��`2R��޻��Wܨ�����E�Z)4)����	 PӍ�m��ː|��05��w�vN'ϗC�!AL�fe�bҹ;�h�!3D[�y�� ��Y�)��i�j��8��E�`��.�h7��mKt���#V�*L[Ho�yȐ��z�ڡT;\c}f�N��_ S���`@�lku�]�� ��v;rs�?H �Ǉ��lC��x��C�A&`�>�?胄r��O�$'&�p.���Feևs����0��k��1;�7.q�-���Ӟ���$���Xn���R��{��r�vb�n}p��`��["QmV��B�������tM�g�;���T��-��<�w	�ujC�L�UM�QV&�D<����*@��̎�0��4�P���Y7��9e�����]�b9z,��ꄅ��2U��}��� #�<�R��I0�����8k����?oϭi�۔z��P��kg�����O�3��ZҬs��Aw3E*ʬ�m*�x��\F��Ln�B�ᗯ*H쬙�w�<M�{U�A4�p©�X@��6���R7�}LLs�M��f��-O �+�`L�L�X��_�	I��;x~V��0)������XΘ+wl�I���|�p��S����!]��*��Y��97,8�:O��V�t�0�Zdj�<��N��dS��1ՙOkU��,VQ�J�+��XǀZ.�Y�8�/�GA$��;��I���wR:�2�<B�u��K��E/�0�-�����*R�T'm��Q  ���"ө
P>�|�vM63K��$�N�N���婝D1��� ��pKGd	~�4(9��ٹ�w�q��RH�,*�R٤�����6��Ӊ���5h$hg1��2D*$?�U���PE���e�o���%Q��@���b���SJ5Y��Q���#�������Y��/E&�	�.�jw':t_��n@�$��<��#q������y���V�$�*�%�v��sx�s��ϴ$h��<R��K.��yf�����+2�6�~�S���|��x�ϣ����:j�,�!In���쒧Xcg\È<PZ4�;�<��?P=��h��\�܌��o�OJ�2s���ܤR飠x�TC;� Pe���"/1@�P*�+{.*�x鑡����}�]F�h4��0��kB��9\r���\邇I�����TT@�ڷ�W)-h�ra��ve~���aʇ�`�t�0΃�9bN��BN�>��Fٲ�::�������8e��Oܨ��G=-pJU��(�Y�Y%%���`P_ҿ�@ �b��X�Y������. H"F<�;��)��6��R�sv����
��8@���93�GX�`û�/��%��l��3�8p���A����\K}��|��C�m<7cd@;+R�^��K<"�>N�ӂ^ޭ���F�G�{>��"�̻�Y�! i�i�h��o�7 F��q�*���ڈt�M��˟��7=j�j�?o��-�^�:��G��L܇�鵨V��LFC����`<+�1@�_�0��>o���X���~�P��7j��	#54규��q5��~3�	Hv�0�R�\��r�b٣I��b��k�|� ����'����?t	�u��v��+0����Qd�]���BV�op��{���2ϻ���9�������"�a��:��r�k0��d=fm>򝞠�	�ٰ�P_���]̃D/T�jt������EȘ���u�����b���d W� Ł��\�Yi]���޲SA�x�#:҈�2 P�"Pt�=�S�95l0����q���W���X��f�ڙ ��r��1@e�$�4(�~��̣���*X�)͛�k��x�b;�$ 	 �E�kH�{+|G�'_�����#TN!�
�5@����?[9l�wT./o�$^�ڳRE������1�q������^?����iG�V������4C�ԠN���̵
_0�N},%�ŲO7�H�
��l��H�L���s������^38rr  ������U�}h##B����\RU9����0�i�[��c�"�J�R7��Z��`|r�.>�@'�1���>	����0e���!-ASmK�u])�'s��6�]�gy��=��~�i�|}���i$B�a�k�	G��kȓI*�yը��w�YRp�Un�:󦞈��p�\)(W�MJ?`vx�O��ݟ�1'�Е���)K�%���V(��[2F��e]�Dyz'�0*�{:-�2nc%}�;
�U�B��a�.�2*��iN0ͅ	�a�{�f5m���Q��g0�ܰeAg"���SR�==�-�Q���$�M�Ɣ��Bbb�<��Ir7�0��-V:4��o��̘���D|[N�����:15W*�`����n�`ZNN���!����لΆq�\5��$�&������W��x��Z���I�C��H����v�=�o��'$�,�!�G�}e����>����u&���߉-�_BAAyV��m�UA���,�4��u����$ۃL���Hb!{;;�H-�<�:?R���%P�,���\FDϝ?Y>��TB�yk1]�Әwˆ��a���
�W��m�g�
l�c�w��.I��i�[�'D�ˀ�(ZC�y&�S��Q�>+�(�k�V�i��bt*2�(p��>f��R�Vt#�)~��y��-6L�Աʙ����9=����K�Y[������%'��m��^��怱(Tܳ�`�a�]p��f�N���1��xGt�{P�(o�G�Î�L�7�Q|����\���u<W>������O]����5M�ް���
�*��7�Z�p����J�0A?1+����Ӈ5(�9��-��.��&QG'�����P�����YH�e7|��h���EX�Q�"bpݤ<G��8��q�垢~��f�1K�Q3�$������x'Gkdj��I/�6e+P�ՄzO`W30:v~��Mk���߃0�H/��d�wgף�
=bT�1�V,닰�K�d���ӮN7k�6Ro2�e3'8�ڲ���"͡�)�n��~��L�3���z�+)�]O�G�o��[9�fH��(�<V�u�IXտ?�����(�=�B��Uٳ�Ѱ���_����B0�)PZLs���H.�O�|��)�T��fSg�k,
=C��F�.u~	���[�~�g�)�v��]�V��S�T�{��|>�z��&�5V�ս�7E͜�KC�Zl.Y�n"x3��aC\GϐES��E�.����x��cCJ�,���
ڡ��;�n����Z��3�4�:�Oo�w��-�.^�/��{�%�{᠒�7<Hn����r�{���lE	K7נĤJ�Yǒx��f	d`��E�X��4M�y��a�A��2��O��5?�Y\B�!.�*��bo�o�����[@;y$�OQ�U��ך�s����Ѐo���r�!��������W�/R$B�6�!H�pU��#��2FB��"Ì�������<$�Uo���l�0ɑ%00������
����,dtL�J�����X6M�N�,M<?���"_�XM�q'=�޴�Rj��'\�+WW9l<v��-���	��१�p����$�q,�J�E��o�"��
�������I��@�A����(A
�;h�|I��m��7�z'���d�&��ԵL�Nù<��g.s�������܂��ԓq�}@7�q�B��<��2�1��'Tߙu��Fz��=��ԛah���{��%���υ+a_�����k�!mS]H:g�:{��JW�j���-�ʛ��t�²D1���F`S	4K
�C5T�:�Ջ��l�?5��x�JZKK�I��%�Ƥ�8B���n9�Kû�l�(�Koi�c���]+Pz���1�;��H�B��OX=?�Zɸp��bw��*C�����8��n:ը������D@ӽp+������ZI�,:bh��H�3��F���3��;ȫo-0/
���O�XSs<��T8����<��r�t�Ɣ�ƹxO09-�����F8|�P$��rٴB	���ܷV��2�#�FG�=�Ցz���G�s�&c����(�e,�w��9����Ϧ����㠨��$f?e��-oÏ��y4��|�b��_��7y��J/��p�sF���b��Ba>ftmZ�$>��j*+�;�ǧ�&T�z8�N������DM(�&O�� -��ޙ�F��:�����E�&���^�bޓl�?<9N��~�JYGk�� '�%�������q>$��i x���Ǻ�A���2p�����Xm��P�;�?S��,4�SM^Dz����֥�a��p��K�(7w�1�L�F�PF^kU�0��e_!9R��x��g]ڻ�8���5���Rݪ��E ����� �K+@ba�Ĳ42�#m�kL�u�Mp��-	�9P��g�ˀE��Ϣ~�eCph�{�T������=����Uq�	�*7Xƅ����N_X5R�����9Q��H�a)�=��xi#��#�2a6F�y�8lڔ�B0�3�>�3��Fb�R���1����c;��VZW��ʙ��'����Gڧ\0 ��'��am�LOr`�"����%�2�Qn�(v��*�'����m�aU����t`%'I[nC�x��2��0t�/'�<"��lE����Ϙy��#����5��|~���T���M!2��5ӌ�(�sR&���6��ӏ�J�
�>�3,az�i�>N9v��E������M��k�� }�q$u,Ț��;��g ~��d�.lM�y�ƞ-�vZo�k5r������,���q^�7�J*�=U��z|����y19`�u��folGx"/��H_x3����&��ѫ����J��m���E��%~+��暂�X
x���m:�x/�Xt�����
;�K� �W���! lz�&&�n�>����SA�ڱ��͞�LQl���W٧�D�<E�v�]�i��n��r9f���%2� �ӬK�����ʅ{<�G�J0�"�*�;�/����$�fq�.�N�~F�����\�ep�{�0�Sr<�d��|�LR$d�_�$���ך6G�0l6t,t"������γ��p��*�oN��j[<�*��� ��c�yH?r�X�GJ|8�
��}�7E�� w��V�)���C���{�O��a��/��͎��Q��P���e�@��<n��|n�zm *��ᘠ�3-GM�Ɛ(��ה,���i/���e��|��.'�M�XZƗ��	�u��p�*G�������J�L�(|���;r2�3���~����3+M�Cx��UAved"��8��K���Ľ7��O�7����
���"��1.�rv��cu��a�\cǷ|�����U�Rي�;,���>���s���ɺ`�Q�-�6�w[Ӄn�V�V�d�Q1#��>���6�h���[�H"�$���n��JM�꼭�{�cw��'ޝ����u�-��Aݷ��(\��|�<X�Bo�{^X�3#F͏#ǝ������IB7HhNuO��5����SM�;��;�|�y��:��z�[�)�k_hh_H	��b`'��8���H��ꅎ���nT�`�,ڣ��oW�&m��t�ʷN+�F͉�
}Iu��83����K�bK�8GNA�j�'|.�6<��YM{|�Q�۬y:������e�.���&Ε�p��;�_��"���k(2�3���r]g����2�Yy_p�/�u�e|�8�H6tF�X�!�s#�i�^��eޛ���J2{���Z�\�"d=��{S����Gϛ&�C�B��M�r�ˊ#D�e�	�E ��v��\�Ĳ��k��6�?NsGI�H����%i#��Dh�Bo)C�I�(��hX��-xS�+t7������NəmwM�d���ڗ;�/�>�9�pf��������=�������6��=��	?v�[u5�1G�ݢ~L�4�v�'��-
M��a��N�F��C3��e��V�8��;rQ}��:z#��� Le��|��ۺ|_�����,���*�.	�Lr�\5Rb���Dύ]����d n��o��+�Z��!�3��4�*�r�of��%�L�����TP�ُ)T���϶	������QO�������U�Ӷ�mh�c�JX�Qf���s�PFw�K���"�vY�q����u�Z���㮍3-�!��)G��&ϫ�';1Q�8�~���5�ǐ�B�5�&��B���&;��\�k_����)�@�:G�Z����u!r�DZ'�|�|?�4!�������*����o*�x�Ҽ�BO�z�RW؄���H�OG�`�%Nq�78�<�I�=���"sw ���lNO;U��(��k=����C�n߷Y�҈`��F��WQ���w�b���#��7W�A_���
�����fI��r� �x9Y��cZg�($�)��2��̔��D����!m)^�\)��tHR$xTz���B���a������_��s3f_(��h%���1�W"&Hj#��_`Q/w�:0��.�wn�E� X���p�/v�z�⡝T�V��0v4GJ�v�[��Mt�"�$�=�U̅�|f��m���hG(������s�5 ŪZ�l����(��,��jPlC�JU�X)��\��1��&���I!��50MT.�]a!0CLL�2�CV�֑�H!�2<�b�|�%eOS�c��s��K]��a��n5�5�h��嚑�ǀA	B�/!D2��Le��v���k3�]�; 3&1�[N�as��r�`�e��|"b��N�C��ɿM���2��0b�M��~���u�Rϒ�8(9f6^̝,g	n��i��Q�Y�ȏ�1'��2�<�������ANq]�a�ʧ
+�t�OG�|W��;I��7�,g�����&瓅�a����wG��<^Ѭ�ŷ2(�jl���K�����h��~���KA�
]��Eq�ă�eVl��p��/r�rIi4�!�̯e�>5����_F�QYC���u�{�>�=�"�ɑ�O��������o�W�',�;����%�+PΟ3g~n�lbq��{�AfP�ڬ�����xUq+1(��mN�+��{V+=��v�Bf%X�g���L���GB^���WG����p�ҁ��WIwD�q�I�{��5��:�<E�Y'�Ԛ#~��#���a�n�� ��*�1s_��h��9��s�d�|C �x�;�:���G�2k���as�%F0d�"�t�x�; �3yx�1�J��}�B����@r)Xa���W$+]�x�Z!fV�Nh�&~��r�����O�}nU=K��UG ���_����qI�#���:�� �b�]��-v�?<�������8�ң (D{���єPA0�����F9����{q�~�WlJ̶�F���dw��B��$�UU��������";���$�G���~yQH�<����CĞ���������nH��#�t�pWh���S��_����W���),)�`��L__�(�,Qa]'�B�{v��nn��R;LW�v̐֌�3�ST���w�Q��v�m͕v���F:]&4ӹ�h�G�6�t��	�߄�:[���0����r�7�W7����N���<^���ʭ��ĝs�A�nm�2ks.h|WK1@Tr����"0���ax���@k�-Z���1lt�ڰ���K�(E�@��T�Tݿ�1��ܗ���o}��ڊÓ&U�����X^����Փ5W`������&�e{L�c�L$ \��"MS�Դ1�K�#�����ڗu��/v�;⨎��|�� QH�1a��)��PwKs�y��$�I����{�:�r���H��J�v֋ۥ���$�?�o&$��z�<�q"�!z8T/E�����1�VD�'9Z#t��W@{&T�Ò���jlɋ
��7���=r@Y���-*�^%�u�����-_��a��s��X��*�㿱�[�,�F�о�r�	��A�%]��{:�I��Z��"�'E�A3wD�R���b�U����r������y���M�����=��H��c���9��"I ���w:��'
Ё{,�(�A��j.�7z_�ќ�m;��hS�'�0&��3݆+�}Ϻ�0�ʑٹ��u�_��@vT���;�Zv������['�`-�ݼ�4�Q�T�Z�h���ѭ����C�nk${LTK�ü7��(Q�_�Q7�.b�j�f�� �$y��?/��L�Q���?��D���{���.�v����0U)�x�H��ɱUਗ�(�M�����o!�"��.o�E�x��Lk��
�K�3��Ԣ��w��:�����R����I��B�I����i�ʯT����y������~�!E�;G��\bYne���1�y!|j�q��0E�o�Si�-��%��K�lY<���!-��B��_��ڶл#�)���S�_6�����i����^%�a}[�W��;'�MtZ䵱W֞�i	�/��o�֠'W���d��`��"�%�0)�W�n�X��j,�WT��s������ز.��L�L��PS_%���i�L����0�vʏ
"��ܰ�v�1=�]<֊��K9��̦����k>��n �#8:,�r�o�������-.vz���`�{#����p���,��������ݯ���-Dk~j���.�X�sy{+VNmi.#p�)���痣f��j���ݪҮ��W�-N�W����o�S��һ���CB��)�
q/NX՜�!޾V��m�L0cjE�<����u�a�s�ue2��VmO_ںhó99i���zEO~޸�}�������M;=�b�W��2�Ǌs&�|s�%���R�5�$ [�P_fH��F�I�U��p�8"���ui##������è7i�P3���:rgdG0h��8�½�_G��^�<��u�[{j�T����6a��x��vj��s,j�[�ߊu\cs��n�k@�EY���G�Q�1��-�v���Φ�χt�>0��Ϊ-z{{ɃM�kӇ&U�O/�֬D����m���>�^��-
7��̗�ި���[�M���{����0�1ߧ;{W��\�8p�䇍�oH��T8�{������|bz9�B.ȩ�u�G��d���#z�'�WY0ɭ���4H������|
��I��)����x�c�6iG5�Xp7���ߣ�֣�sSʫ�	�I��#��%c�SKS���'b���R�K��5��q5V�DRx�}*X�9#�*/�x���~z�"�XCS��4���ٌIߒ�,�^���Q��n}	o�/h$��Z*�ҳ���R{�k�3��Y�����$����\Oף��
�j��ף~�"��\fdx7F�!�Z�yb���D���,R�W�"�{ڞ���`��\�{/�EW�C��ǖ���ah6�%v��d�*��$ol5�$.���a�Ýy�š�,��!9������Ze��hmpM2���M�g#-�T�L�Ja->�T�����<
h�R�d��(��j�^��A�V��+8O��s����j806��&�WZ��V|;9y]I�<tpY�����ĵY����IJ������4�`��h?��[�B8*�e�B"�Nm�|�	�DxӺ�*�ng��Kz��SxR�K�qy�t��qHb�!\�1ZМ?~z�˷(�e��W���]�����z��gBj❏���Y�{��5Y���i
��������˝#=��}?�d�}2?.�ɸw���X��ߟ�~p �;bn'iE�u�R	\zJۦ$�3��.*;���}/��2�t��E��I[凶�m���!�|^g�[[��z�rp`:U��lx��OrO\7�|C
{�'�$g1����v`p]A�DN˲�4���2��˫]g��{w�l_�F �;K���3o<�1�Q��#��9�I�s����L�yNw,��%��k��XO6�����\Ҟӓ0�����D���F���Od�X򻉅�Dc[�ը��/s5ڦc�];��[ �/��^!M`�'P�9tȰ�������w�"g`.Z�ϼup� ѯ謴#����_M�5�A�%�ͮ�5�4v\Г&��N�Y<VlƁ-pЌ�aX�$���i�d�L�#R'NbKbD$á�rE���a�l���x��"�R��-y�������q�A���ILG����yN�u=G�sŞn�Y���p�?�{��ۥ	�����`���N���g�������Q�B�PN�+���M�I���ӥ�d�,�D���k�_�M}�"�BwWњ&�:u@j��`-�����-ʟ����v�Rx/�0
1��(�c��A/�	,-����	�|t��|l���/����e�?� O
�m�i��S��t�'�,���ˬ��T&���:9?���y���Y��p�:��	��^foE��v���5QO�=�(H@	�;�����I')�
/Y`j�����w��b������Ϩ�`=�.��Z-4��Ʈ�+�J��r2|��ɚ��i��N�-:�7_��~@SΗ�/�<�ji�>��<�����q(�ư���x�I�����8�̾��P�?��w��X�EDFx��\K�� T(��sӲ)[`��mC�Â����[a����+s���e5�ي{�c��}��n�}���NE��_l<��g_9�$k��m@̍LʋڔީTa
�mHz l�;�n��芖�����rh����<Q�a���x�X���\c���<�|l�����]I�X.�T��%c/�lX�ԧ� *n20�����z��jE��0eb����iD��f��7�`�@���0�x���sũ]�V��A��-M9i��ċ?�aG�<>��G����_�M�빟m&vIv39ZP}XXI�h����Kɹ��(�SW���˷T���/u���R��`�U"�����!/���t��"�O�4<�\%�S�(�~d�5��?�l�ҡ�V+�1��/OV=Q����/���4��1��g��l�F�#>o���1F�|�&q�29�H�H�`��z�OT�5��7VӇ䷑��E�n�f�]j�����ǀ���j������-��S�S^KA��1Z1o�OT�)!o&�:BdG�\��ԉ�)kO���q/WK�;޶�)ǮR����E�����C~������e8�l��8��$��Vёc�����L�C��I�M6%�(�&�)��V6v�6�jx�h��H,�kU[W�a5�3�W�4�:�\����O��T�l�BK��k�1�~$/�#�b�>��sJ[L���9v,�ǣMB���������B||Oi|�i�?u�@C~�@#B�p ���ٴc�g�)���]��g_IjP�3\	�}��N���X��M��Xo�GӤ�8|����T[l+�Ue�9��g]4�vxL�l�'�&�>b��Q }����N�`c��!D_R�-i/6��	;����/�~�_	��w�!�z�P9c�"�F>jR_{�5{D�>Рa*�A���î��L��j��	lw��6�:�K�� �ٕH=����j;�gs���������wF�)���/�7�!��"���E�o�Χ�,X��@�Ӏ�>]c�&F��p<�v4�M�����&��/��(�l�����X�E7�*=P�bv��Z�%ȷ,�ë=�>F�Џ2�#w�bq�uF��{�x�U� ���U����B�ܔ����h_+԰�Uј��,d�c�v�,@�]R�y��2Ь0[��$� ���v��m<6f��ut�&��e�TdA`�͚�'wxO#|�3w��L�"*N[Q#{���(�T>S�&��f3�~r	�ኧ���%1fۗjDv���1�0��;K�p��~�}_P���l��&}��)��w�"� ��5���ϊ���$�k�L��R͐E��ci��������ő�)��xh�i�uh3zV�fT�q�l�?�`��C���&�՞q���gS* �����ۑb۩�o��N��"W�k<��>��v��N�_v��`׮�F�J��y�}E��E���L�4t)i��(��ڳAO�c��t�K���C��%�9��r^��!��%�n�J�\�UH��
(Co"P7@�������w���:��UR�3�{�y��FbrΩ4׍�-�}�c����*P.,>ˑ�8�A^6mnx�X���-�^/���eR�N�N�!Il�hdz���N�h����t�Hb�޸Qr¥U��d���C�w��[-����^S�ʺ�i���zd�{挵O�UAE�'�b� 1$ �k�x�ǥkC_\�S��N���?�Z`߯Z�A�R�̶O���Ř����Qݐϓ��#QY��
�T�r����i�Ct�5�j�"1�-r	���C�
�5�d�"��EJ
���2�OQ�>�xퟀAۮj���f�f�*�M"]:hL�#C������U�� �$^kJ� �\���>���V�F��xL���6�����ρ��� ��:Q�R�n���P%�(U��)�������
_��D���@���|�>�2H7g6A�{�+�� � 36y��K�0����Ojf����+�[�����p�æ�k)�~��}�뉐EYE�OͯG���߳�΃%����-�����*8w��8�iK*#AO�_"-�  �^~/���yƛW��΂�%��"�ϩ��6j��2�5�≽a_��,�aKsY��B@ �Z�;ʂk�R���H`N�d� Lݦ�|�߫v�"�l��7��w�����a��X���G��ξt%0�9+�}P�,=u���Cu�t^^?� �A��)\C�"�5$��5~�'�����>R=ɏuN��:��V�]jGNmG;���˭�[D|�;�M��S H��A�dX�Y=BM����\a��M�0����~�����)�q�I�x�L���N?�D��kBχ�c@��X�,�}�wJ	k�:�A�ܱ`$1�w�$����d#6x��f_�t���&��"IP��[%]ߙ��f�B�r5$�� >���O.�*��#�y'����	������gz���ՐE��޵��iڌ���ƹ��!.��idZ+���~�O�x���bi�4�d/0�0ՠ3�h
>�X[ԺO��^�6�!axw���3%�����5�"������}`� ����n.2��#{�X�
"0�)�He�Q�*d��bmA�橯���Q7���v;�Vp�]�N*Y��6�NB�2�c�>cs�'c��T��Dj"F�
 ���6�_]��zr���G��gg�#M�
�w�﹀^~j+!�.������=G��]2XD�Sp���
8�Z^)XY�!x��<�"����k���x`a�\C��X��>�F�S�6��P}ȞlHg�=`5�^��/O_��;�JڑO�f��v��B2����_H��}����F��~�G�Yb��g�R���9���3"$�N���N2�eGE\BEo+D$���x<N/�N78h�-��X6x�wD-<N��*{��M�����B�y.p��Ů-�\K
nm|8j�����D���UuD~8ı��,z����YO�YT+�_J��ԘsI<,!`�;��bؐ����脲�������� ��Qt��і
���\�#*%�������y�:s~�R������-Ԝ��A]	A�M���;CT~K{�i��	1�(�#V��a�(��ln���x2��Wў��/Rj��4�N4@���Q�p�����=���N��t��&��������/z�To-���!D��74ީ:�ld{N�c�%ԇ�2`�`aC��)��u*���,i��#����A�'�(�2��`���S������4t�IJv� ��F�h�
�����Į�+��?�w�j7J�
��*���֤	�O���3��u��o8��'�fJ��F�.����}���/�Q�S��!�V��#�S��kǧ��܆��9�����V5�8���*�)��D,�y��#�����eW�ѿ��^��D���S~�I%��X5��X��y�����/��F�����D��H�i0��
�v��9�{�]�<�ӯ���6���Ȫ*WFp��Pm�]����C�Ai~�D�Ϲ�,_.��&�hr
�em����g�������Au ��#`����>�|���¯@܍�����IX�.+��k�&kΎ�bJ|��D�fj�VZ�aͬ{O	�� �`N��։�c�EB�C���+Ry�M{��Yٻ�8�
u��9b�܄����'�?���tf�����vF6��>�O�Q/}�A�#>�U����מ�'��z"��&Emj|-\���~�ydҵ�V	�]�U��
9�l�7��?#��Gq�X�p�����sY�(�f�Tv�U��W�)��p�'��r����� 1`�l�E� 	�_�nG���YP�M����� �񾓷��LK�w���e�ǾB�:\9B �+!m}�P����f����Ҙ�(]�,-�F.��Q�$�$w�T�hfR��wZ��䙴d��Q��<�^��5{v
p\���88:p��3���7�os��V�	�����&I����x��~�%?l��iQ�%���;,�	3cTF������xi ����h�`[��!�B�eO��d%g߻�E�'ϡ�@���7��$g"�J'`�[o˻%�-��������TPE�
"Ih��L��̶l��:��O�D��Z� �Z%�����AC�#~�-���� ��އ�(~[�:!,�~,	�X��.��`5腅[�|�<�0��P+��>�g:.6O���`l�{%V[?\�^�7P1I�Q7&Ήc��$K2-Dh��hLbj7���n{�ÊsG�v����L<$�֪.)>��K�d�M�Ֆ��2y�Jg�4�'�"������sn3.������{`h�ޯ�b*vD܎��B��}@ݸW��#Y4��s=|�2��=��w��N��Ğ��)R�����=�g#��t�������rv���9qe򭐪in���$��G�$m�U�gi��
=�������c�S��l4�w��*D�9%����� ��s���.=h] �	�ӄ�~lG:�������924����5[��q�U���`��r�����J<y`d
]�2kڬ���4�>o�C��1�ڳ�h~�h1@���Q�t�(}�`|-��=3b !q���ƺ���~Xs/�Y�B�Ȉg�9��o��3���s�&�'��3�1 6�j�Ѷ+�9޸��_=�u�8c�p�Y�o[�
k]�}¤�C֒j?[��+M��'��'���&) :�����I�#3��zN�;)Zhk
r�XNfd����eQ��i��V���9&��n����iΛq�n�1g������2-hm��%���X���g\t�Y�s]�@)��2��OT�_�X�Y�����5�O۞7��p~�v�����2�)RU7!I��H�2E�;s�sx��%�x{��3� L���A�j��c�������D&ȿLi������_F6������(����54l�u5g�0V����k��v@��&;Ix�PT�Ċ�ĲLo�g n(ĞsuVbY@��'���b�n6ƹ�K]���|Y�A����]�:ڝ�2�Q���gq���;��s��Ĵ^z��'Il����_�xJ2OԊ�
(��b�q��R_/��0u8���ޘ��Y�5Rm��� �qpe� $���2��ܠ�M�mH	�W�?��3�4���E&�k�G��E���AI���X�ؐ짳�Jm*�Q�/�d�->H�2T�R�ͮD�,��@T��}��E�zS��^d��'(n���H��������{� ^����DJ�>&�vyڥ�r_Y�����- �B�_Z�M�����Yk�mc��A�@���
r�a�c�[CW��ZS����ż�z�^��s�.�r�M�W. ���L�d_C��(oP��1f��/�?���;2)9�q,uo޻y��>��8Sr�*5p��6� j���z�K�֛t���\�P��tt�
�v�>!��B-���Q!�T� �;�[ђU3���	�0��>��,�����?��7��,�0�I�%��7����&�A�sG���,�P�C@�O�2ouXj���7*�?6����'���_aJ�S�}��!١��	����9/v�X���h�Z
�'�٨���eJ�V�>�B�>G��<l�`s(wT[����i��z;��8��l��St.�K3��8砃H�ދ�g�fJ,�ti��7�0��t���-g�~��s���6� ���+����&8��}�Ϳ� գ$����]=���V9p��� �1�f t����*e�ƮE�5�s�.�	��W��C%��}�U7I`u�yK�%���N!���ν��J0C����=�0Zޜ(��|��ڻ��ۻWŉ����ed-��z�d`��lLJB���t��K�R�9�wW�	���t�����@,8�>��^�y�M�rʥ	�L��j(v��i��^m��1 zDK:��H�Ud��<��X�W���B8�e��Q��Xϼ���[��åo�8]\ �m~b�!:c�����t�����Y���j��f���}��C���&�����ƈ����s�������Ķ8=9�}��:&|U�+ŋ��S�J��~�e���K��D[~�¤����%egPH�ۼ��G���
p� Մ@ԽK�ר�C]��^zD�,��.-�x#��[�6S�tݢ	7'��`���t��zB�����]~��� U��l�'��W��y(q�1��p�uW��_BP�'��;��K%��1h�m����k5 H��N#n��ɝ"�׊��#��2=���Re�sl���Ͽ�}�L��~"��5Y��6�r��bR���&����Ó:ܬ��L�:��Ш�t_)a����ج���HRe(���+kã��ٛsIl�ic�O�f�DPR���k���s��i@��"P��mir<��$4[6�C
.�V�Ae|�6)sl��:��7��}!G�;�%�aZi�ui�h��q���`Ȏ�!N��^�Z�C	��E�(��T���qq���������uq���0K i,i�u���U9�#y"�ף4:�.GQ�,xӺ�A�{���kb.g�>��$�����	�D��Û.�fP`�X%1]al�TBɳ����t�F�k�P�?`!D�0��"-\�S�D(���L�,g݊B*Z��UT���0�]��Њ�m�9);�Z�g,�����`9�:��'�\'�{��� ��9�������C9�"��q6���������JyW}��	�;x��LVr\G.{����J�����}�dl�)����� m�����ӌ��&)X?�!�zn#ue[l~r}��]{��T�A	�M�e��_��� w
�p�E��A��GK	|�+bH���Wk.�# D�*����.�"���X�G��M7$�+��O�Xs�vOъ�;�L��Cs*=�����?�p��5)���#���$�,���s�tr�2��J[��Q'Q�9��܌���t7 H���Ē���C�n���$�ٙ-�W�����+]��w�3���g�i Q��xeA5��|�Eʐ2��B��4� ���#+xNVN�ֹ��֩6}��K���y�Tr�V�!s4�#�k�-/| �hJ�**R��p��3y���q��Y�Y�\P"s��Ǒ!��A�i��ױs���`�8��3�j T�E�5�ܸ�hCN��/�%2��+D5c��"��Ow�� =�&���Թ�|�+7+�Sp����Y��K�T�9>Tȃ�'��cRNW)�C��#�P��:���vI ��#QI$�һ�-�����N����IK��Y3	B71F�)��-���@��b�̮-룴�B
@���͂/Ge�#�X��.���g�m4c���$^^<~j�z�fR7v�m�ݗotB��1M���ņ����O�!��� ���0�LUs�C�(�B$[E�!����'Z�ڼ�@�l�Q�@п	��������ot�&�AI�X[h);&��Z��;%3����C��5I~�g�Ġ`��H�H��k�����6�ek�-쉢�~#�o��P�w���i���l�~�;7���a�(�sY>_�C��&.�B�7pP�����Iu^!��sb� )3L��,�����*��o)\��΂/��'El�] ����f'Z���Q�BdFВ���SP���]�#�a�:D��͑���N�RԔ�l�e��$=�+�6]��L$O�4�S}���_e�I�R�Aũ���kfȠ$P�Q:?���Q�7�7(�s{���y�>�Z��WXU�}��m��!�Z{���LGNY"b�;6kM�J��ia�Iy�bMN���Hgp���"�B��<Vf:{�]�@P�J
���İ��f`��#z�_�p[�#[���?�j\��&0�q����_��r�0���B�:I,�C����'�uB���Z=�0��4x��!L#��������`��4���h _rI�0k��D��!;�K�}���)��f۶�x�d9�g�a�8���	��Oʨˢ� �Qv��q��DZF�fP�TFɨ��N���>��"N�unW2x����
��[�A�*��8so�|nk�W_��1�!T�Xm��H��!Eb �~Uj�ۗ}�	���*���+U�mh<��DА�%��9�%�<ݠe{�=�St@H֛)��DE�	#$z3TuP��N����D/�X�ٱ��*ܹ�c�I��a�0	O�`*����fg��W"���[���޳�wƠȉ.�G�rY�khe^E6�v��z�`�33��a�����Z��~� �|#�F=N�	"
i�"=~{a�w$k�]l��� �QV���E� J�;��`�K����(h

W��ef2��!���W��^��Ax�7r�,x%w_��*|^%�r���z��Fا��c���#.�e`�j��.�ӛ��=�Öv�V��;��s�_��1z�Q�G� q��b��.�k���{rzz+^�z(�@�G#:*M����<�wC8���]��t	�:���[��j	5���B�S�R��)˾!fR��-yS�)$�ΩLj%�}ut �Sؚɑ� g�N��	������h��Rk���^}�(����攱��Bi}�u�L�K���:$�C�+$�7��Tū���B�#�S�)�JK.�^�\����9f���|�̳����b�grH5���>Ⱦ�Ւ�n��V���h��f ��惚0ª���	���:����zd�6��ń����L��{�*3I��]D���^9���(S�˾�bk�`�??� �cO��{y=_��[߂��`is~��3�k��_B����N싖ii�&5�j]�pnY��W3~2:.#� ��8�1Dv���s�q�G��g+V?%�v�ÑW��d��G�N�'j@P�hͭx-�o�EZ<���;;ԙ��.��!��e��C�KQ)�����m >�x��j�K�CC��e��x�(������y*��*�3V���3vq� 吒���Cy�p��@b�& J5����^�B�X�:����B��9_/~����a���B�A7�3~5v&�����.j�������d���|r6a�k9��ME�#J/Ȟe'ڵM��p>���@<J�[���zU:��+�^��ts過���R-�2�Ս��)�ց�xb��9�|�r�^)�_�_�N$�7
�'����T8G��P>h������x4�}��@nC$k����E���������!j�:�/>'i�&�w�)����럸.���};��z7E�G3 �y�z�A�a1xH�&e��[|���ՒJ���#�	�����@��{���(�8�	H�Vl`e/�a"曓�8��s*�>Tz:"Z~���Ta	Z�R�)�_j	��d2 BS�jy�L�bX�P�2�Zr˭���[��A#P%�Vٞ8�͞�dJ% �Ms�(��$���ټX�Qb�Z���¡���?�j�������]V�w&�O=�EV:#p���s��7���$f^e�S[Fa�s�C�m��
��dOͥ�i���m�]=�&W�^��b۞v��\�'3>���dLR�	��(Ǟ�y$���������"���t��ȝ�Y�������/�b�t�y.���/�_m���D�bx6�r��v�\�cڞ[PM �	)���[����+66"�_S]L��ǧ�����j��
��DG���٠)֜/�[4���L&mf�dz�H�aő?�E6�}�xԗ���0G��/{~YCޝم�C��-1��GcL��f�<���!�E��x�C�xi�����0֠�=��꙱+|GۯmP3��S-d+�ɮ_ 8�a� ���?2;sų��	����^OI��{�jr��b"�+�D?�hɮ�b�}��%/ou��P��x>��m�f��\'/`Zۡ!QX�k�ʕ�8���;�������hk)�>��n��m}=R��G�abw&�{�s��y��:��N�.�풰��
m.�ɋ'D��ԟ�����ř�d��灼C���E\?�z�Q||�&#�!Z	�*�V̮��^@�l(���c�5q��9@��I{�����3{�U?������>�[\ ������Rϰ�4�<W}k?�X�K��P���.�LOj��ddW02@d�B��g�ڼ9�9/5�k�d;���+��#V/i;pv�VB�iD�O\A&c�O�A9�9>+H��m��#���L���ÝB�u�}~#'��-̽�|fpŷ�x��߳���B�8xT�j����u(�;9J�Z}m(��H�ND��]�����;Zq��E�;���
u�%���Ɛ�� ���V~�~��TF�k+��5(y+8Uu1��c�A9�"���(�+�<��>�#1-(��Zݠ(Z�.��0r�#��u�	D�QW ��Y�#��Luo&��b7�0�7�+p*����=�v�h@��Py��j����Dn���Sq޳Q�2.p����{�Wߊ{�Sm�v���[����l*pƄ*Ri"~E'�	!�w�sLKu�gY!Df�A�h�p�Ii<kk���9�#`6,%����s-�6��I漫�l�6�?d8�E7�C���~[T��A�2�Qm��^~�f��Y�h�e�x�B��;v���/�8�d���D�4J�0��S&�q�0�\<�����VIʖ.��m4U���_�ǁ�"���t��	�+��T'��_��Cbaҥ���B�r���s<�Z<�N��G�,��iʊ�Ő���<�8��}�J�m�#��,ɡ^��h�.�\��9���MgB����~�	�o(4����_���7�Z�I�4Hk1˧���#�X�0��P�݉�w������d.��Bч{,�y�YJȥh�'����0V����W2�_�)/�,�F��R
�"g������� �����V�^�����|�D
C��oPDO\'��Cʰ�z>�,w�Q�Ҩ�����v�zC䦭��}�����}� }bO��8�?s,���|(���X����%/��&����lg����QW3��[VJUBD#؞K^�2�`KV�KB�Ű����(I�-d/_���;��κ�����l�k����C;}S�{�V��.���YA��l�J�W8����,ݭU���>�`��`��
-�������3w���	Ԧ��jK�HB}u��_�2�3L#��f�a?�g;fP�<0+�P
�_��B��MZ�
�[*U�Y�O�.� !y�n��T�`m��C��n�Z䦱�_�VuyHs�M�<���Ϛ�� �5����sӟ�~}�
���kw�z�Ü�0^��GK��s��x���_���g*�;�C 	���̾0(����up���[�"MB�*����(umd�h��}�5`(#��յrn)U�n�@�S��C�A�[:�i����Kg�6�����\����W����� ����d `��فu%O�rC)��{5N��%��r����S��M��N4�}3��s�`j\֓��=�A��!��R脪��W������0��r�1=�-j+aJN�Lt�j�lP�W	�C�w���D���w�d�9���u<��;����P���le���ﳄ��3�6�k=T��w�����N���Gd�ɽ��5�'b���("-,�A�pʡMz��|�B㍒�Z���F��)iv�7�CMּ���t
�Վ��y�v	��zf@����M�X{���q�^i_�����^_�����:c��ߎg���T��"���p9����'�����~ =Ν|%�W�+�\�hh)Ѡ��*��䶓�gb��vgi%�11�	��s��a�s��(���7�����	���	5�Ӡ�WM�x"�/�0f�x`��' �+_����U>l�SՃ$������)�b�	lE6Tp��[�V!�U=�e��Խ�N�[��$�|"%�3u�"i�~٦2a������%e���=���U�x��Na�F�/+�����\SŒ���0nՊi��*?r�MoRjO�0���ȣ�Z���c�\�i%�ѝ33��qos8
݂�Wm�����j�D����a�G?����(|�9�r�8_�f
9�������9��a'n�Wt7K�u�no2�#�Hi���Z�W�\8�8��?���E�����3;�ӄyJ��L�k�WPxݦֿ�;�"=�TJ[~���1I��H�����4[��{�U�S}� b�ؽ͹�s��j�%�A��FȪ�d8������X~2�1Vi��p'V�H��x5#[*B��.g��Ap���V��6��씰1&.۾�jA�;���7d/Ub����fkT���΅xw?:����5�l���~_��J�+��D
���/|�ڮqQ�a�ҧH���bS�Lhґ��iӖ��Is"w-26=�����h�@@��5�2��������`�֙���Ё+��E�����h�N�={m{��3	M�j�$)"�1� �5;qڈ�^���ЫN�O��D����9������]�9$�:�&�羢�x�R�ERb�U��)�Et��h��"ܳ��ʹ�Ÿ��(m̷c���;G
�-Ǥ�h��$b͢qbû�F�k���[��0QG���&�'��E]�OS�?���q>-wd�:����g�QWo�a�MA&7ի��9���l�&?��gK�H�!g���/����F"֋L�^��@:��4���OJ�D�G��"���f��[H�ALk"W�:Ʉ&�@[��F�ʤ�r�T�U��_��[�\�{}ï�Y���:l�0x�*��U�=Z�sVm���[�ZM��
��(U¿�w�K����πJ��K+����m=Wj����乃A暡�jq�r6$��tk,�Y��Į���ִUr�|�=�q��'��N�I6A���Y�8���b<�q��4����R��de�F����l��v6v������=�����ӊ�:2*9��nТ ��裺���>6��|�3!/9�m7����f9�v�C��ߛ��t`������j�'����e�����8`5��I�ܱ�8��s�i�SdU���CBT{���$�S���a�L{�9m8�w�3��<tK����eH��ma���J���|���U�b��h�������Tj�����3��'�3-	x�Q�~QB���������7S2φw�+O�����l=
��<�I?�c��Q4��a���Fڊ�{�<2��g�7���⊻�C� �4x$Z}��qj�ȥ;���{�����S�8:�N�xG�W�	i�Ƶ�Y��������^�-kj>�U�^�T�tR�h�̈́Ȏ��im�)�����ee�:��ͫJ��uI��8�����Nc������3����l�}���[�mP?��ȃu�\�Hw��j�bh͞X����t�a�$A�J�~��Y�o. :Mi��e�]���>.)�C��D��E����3-�����|ڶ�k�M8�~��:�I's�aô��t���Ģ%���!J���	�T� (*^"Q{�&gjr>>�5�
R��S�w�
{&���w/0U)/Ujꉈ��p�(2�#6���.N�*�n�⩪kW^��ۼ����q�b���;�8
�#��:[2��
k�;�ME�����琤��׌[		��]����zz�6fMHy��
����Σ@�Ǜ�5����7��'rt��z9E�<i��������Jh�Gj1����z�O�E���?�W�K�,\��y���c8��O�5ܟ�fm���ڶ�����n`Ȼ#��������fQ���=� gBӷ��È%i�9Z�ˣ�K�����ȝM�]XA�	-����<�Ӥ������l��V�f@b�{%�00Ҟ=��8$}}�T%�M��N�z���&j�Y褿rA�Y#}�L�sK���3޸�|&��.S��%����������x"�U��n�����N�j����t���D3/ݱ-�iQ٩\�h��	�]۶>bY:F.�� �F�DY�s�����������[�~�A��i��F!��QtK?7"ns�~R�bl�=+����,*�\촤Cy��p�x���p(g�8>x�-�@�<�s�w��T����W��%:%��/7��f�V�=�W8WN���fL�3�Om[@_�w�����ETW�k��xli�i�8�n\���cŇ �n��t�޸A��9"����^ ">H�Ja�(U*��	/#�FKR]\ n��\ͩ���k����1��~)1��FF$���l�Rǡ�N8zʴe�;!-�>����C�#��.�C��H��XqĶ=e�wK��;Fzg���� ���O#�@v�k��� M�,i�I�K�����+��w� 8���ء�h��Rg����yͶ�����&�}��mJ$O�"pכ2�1�*V�
ĵ�[��<C�NysG�d� @�� ��k� E+��ͫ9ڃ�7/W�X�m��V����xN�IB~�,0�����qO�Cl8���w��d�QC�8^��U�˔FQ�r�׾�7��2�5�)��"��`9�M��|���ڎS���+�rJ�K�[K-CBȋ�2�w)�{6Å��,�_ډ�R���ɶ�D����[!�����_�"R𲦢I�U�"�T�����x�0��E�UP���^B�ݸ�9dM� ���|��!ZA��N���;O�.��.O�L���d,�u6�r7���������oR�}� �l�%`J� ��3܏�˴#�80Q�zSWHt�9L"���C �;�!h?��3�9IWW�.>^�
%�F��7�(�R�����^�#f:n��afX<�<���y|/^�T��9��0�m�R�^2�!��v���1��� aV�F@ɬ����nR�1��)� �g�4�U1 �X[֭�Z����⦱H�9L�Vn���8<3��ݬ�}���Hs���4���&H��i\�
{��d��oۂ���r���Xo4 �O$��Q��[��.�j�3���,�2�V[��Oʧ6X}�LN�jK���΋XZ��*�R�@��\r��Dl��Y���2�J�J1ف�ss3\�b�w=	
#�8Mp�F��$��{-�މ�k�^���4&������ibb�гss��1�<݃�&�@	��W7����/Q;Qbq��$v�X�C�����i���A�mpL�ڤ�'�/n������O��;;�A�uA�T�̈�H��̲>���.���*�´���J���v��-���ժ�����Z�_(���[�/|�E	��D��P�}��9	�7ۡ�{",F��̙]\͎n-�%,�V6�S�[�\��Wi��w9��T��̹�q<t�+{� �-���fd�Q���x��x0(ύ {?f�'1ᴙ���{L��f�d�q#_ㄣ�D ſ�cXYf;^�T�g�,.�F�IMR��7kk�dX����W���B�!ԧ�{�DoD��C?	��+�ڠΰds�a��L��3aѠ"�h��	D�B������e"%�����,`_�Ӆ��~V��a�Z[7�3�l8%�ܺ��w��#B=ς<,z�b��-{���cL�n?�.(F��1���#�?�����O7�"�d���]`9^wA���4�����yR��Zs��z�s�<b�k�YN# C���O[�:���G�=~�"�Hs�w��N���>,Fn�c������jc ���\ܗ�˧�	؂���m&;˜��X�\)t�\;��`���W�0� ��0�)|RR�����M�cwߔJ�sB߰ �XC����3@Ę~]��CH�'�� w��V~[H˃�$���¹��֐�,=l�C��P�Ք���b�^���p�)Ms5�F�(�u;��|��d�c�s�����H�e៞���}�g��c��h�b�\��rб8R����h{Yan�nN�:P�\�ζAn�"G3�O�ۙD��31c�g-�~��[d�@�m���]+X&0�s~)����!�O%.ъ���'msf������荻����Sh{2�����H��PDփ�	�����(���9,>�ţ_ Bv��"�.�p�8����Z�������r_�����vCZd���V��*<š�H���X%H�]�ʹ�-A��{H)�����B(Ev����U�
���n�iO�9�nk�,�ӛb����^�7���� ��e��D����	}Jj�,a2�u�^:�^�%��f?���Q��2֩ڞ��~b�	VBY��MS�z�`u&�nN�~�Qr `�.?�v�<��`�E^o�Jaz�D����*��޽�Nb��My�������m:.R<k�k�,w��h}����s�`$N�{�r����cfT�˻�Z#��C��Nk-Y�+Aԫ��o��B�F,F�C��G��t?b-�t���iT�����U�DO�:���X�6�o����_�Y&�L4����nܼ�`��.���~���V&�'��>�����k6��T��\��g�#������㓞F��)u�)=�X����z�3�`��Vm���1O)��N�n�2	�톭���-�݄B��4�Z��B�$����1 �H�3�lv�ɑ"@��8<�{��x
�麆�ḓ�َ��Y�([��Ysj�Ld}Np`ȅ>@z>�.�x����S��E��?q�K<�P�N�k�8)ESR�JIt4��~��G��#B݁������A�yP�,�-�i���g�Y�B9@�]0%ظ7� �	\�6�|C*����.�g���d&����74�_�y� )��� 1�'5�[���un�)����w��z	[!}���Gudl�JiF7v �,ڵE�����V@��B`����P����Ve��H��Aq��ބ��?xUҍxf�գ�k��m��X��Z0�pv�\�-�Dö��}W*p�n}ľǘ.&�|�<��#�d�R�s����ty#�՟��@�!L5������)y��.L���zr�ZPׯW��O%�xE�e�E���6�r���N��*9_=���!O>��/��eZKPQt���d�#�ܡ�>kܩ�+�P0�A�Z���l���	*We�DC���S��������\|�r2�Ϝ*i��9��p_��B�l�?����i�㪲
�i0���`*Qw���{��J���1����<��=�w}�����������e�1�s��Jqw۔�y�7�� �m�=��:�vu�褹�|Qc��#p�U޹.�Dq.�3�}4�rF�]���7�[�a��Ӧ��E_�˙��D�I����v��kfM��Yv�����ظ��-*v�+��c{TI�*�=|m��̮E�Kf�a��go.��(Wa�����J^o�����(6���l>.z�ڼō�����`������,J�<;�+f��q��Y��-�P�W�����(S��������a#�J��]Е4w���e���5<�9՜!Q�x�"
��C�=�@mJt~�	�Jg$���檒i��M�v��qD>T����܊D����0�n�l'��ZlY��5�&uv�)�Ż�0��H��=%fT�a�ܺ<�[�I�^g���%�����9����N{w����z��/A'��![O��U� m�۬�fFn��a�b����i�������-b� ;H9o�Z�ӌ��0�%݃/�� 	fA.a��
��nv�K#�<o�v����&�s)^\�j�G�`�z9̹��T;u�|��Q�qs�b�:��!����*,f�՜C�X�EBc�0�n@��@#��6ٽ�9��DJ����W��jO!.P̃��ZOsJ��-h��z�[�MT��t����Q�-���pK��B�ڳ�!7͉U��+gp��c+�	�@wi]��o��l���)�O����� �}C\NE�Na�a��!c��o�2���*���a��5!�!����a<r�#ך�$��Z�YFcA���IL���A�{��[_���1��6���'�+�)�Y�5;WQr׹X���n��v��h�n��Ō��'��^N�U�G�. !����R��ܡ�-J�Qt��U��-�@�����`����4�Q��o��uϱ��g~�m˯��$|���g$���8��ͽ�l�����c0Z��E�I�WLa|�j�>�7��܉u�\�$���|]F�}���}�=�m��w�l�:���]�� )�;�U���#!m�(���1$K-��^�H���n�zg�bE�h��:2��2nP���1[����onpkҚ�&�;��/'��NB6���>�G`�A�ң�gF�d��<��`0]uN������v�x�
F)�q^�S�@!�9b�s}P�-�o�aU��"����KdE���7Rm"+ )�g�Q4�%��6�Q\R-�w������}'
�`c[{�l��S|���AVL{�I#��X��1�7+ߒ�%e1���y�dOաx}z�<��F_VO����m��H؊X�9��=Jt+o���}Lb<?�����+w�]��
�*��iS)�ڪ��Kx�T6費&�t٦���"\>���P%��v@E~G��S�Its˷S*4�'���p�x0� �+_�>��fXs�w; C7ն��-���#���ay~m�V���K������(d�����!�ʱA�-L����1vR$-�Y���"���m��VFx�	��{�["y�'��r��0�mO��8�=/�����:>��� A&G@��i�A"�R��K�b�@U|��fO�Hsu#����9�AcG�#i�{�<��mU�تQP���-�(�J~���½�9�5�@i��d�MB�Ǟ�-Ӹ���x_��+P�j=i�5�݊fbA:R�a�����5�rK�iw@���2Ά�5��H6-���u5hhu/���l(3��#<��Yw��W�����q�5��0j��$S�h�{k;2��9��"����Vd[(��C��4u�{�v�L�"��:h�a�	uD\�~	7C�Z�]v��)͙˭H?>ĿAX�,^�����ɺ�@���J%B�z�g3�^�"�-�rW$����*N�o�,T��T⓼�*u�eT5Apb��aMSK�jV���?�X������bjP�+�B��e-�
��æH�[O�\�|��Pٷj��zz.H��ݸ��9�
����R��E�L@pC�#%��@P��> �b^�-��׎ߛ4>2�����\����^iVL�Ü�J
|Kd/9>�"�aI�Cy D0W�M���w�w	�3���s����I��t; �5!g ��J}3-�\��cՙ�1%_T̉D?\%0q����7h�����^�	�!I�0��B�.���a$8޷m��\�ͦ��P��Bj�}Ɵ���)�_���͗�D�y�DR^'�!nId̳��Q�L߿�<�? �}!4P*��D�	����eW�ø� ���L��,*�ͮ tZ]�Z;\M�e�f5S���8�����gg�/��e�[�~�/���$z�Y��_���G~�qq��\W�d��d�M�w�)k����˹診>x�g!�ɪ5)�ۯ�����~���y:�Z�DqaT��x���dS�w��R�u�k���J/���b��Wd����^��/���W�����i�w�qg�rJ6��5i�!z]6.ٿ���F~l�����{l�yA�0�G���XX���|%��t�Wn�#�n.�<�^��yJw��70P�7��`�44m�<Q����Sґ��Z�aT�k"{�p;%�~S�,'�*ULv8����bo���0LJ4%����Y[��v��G�7��2b zA��eh�J&܌��	t�z�x��v9�y��1*�2�,OĄ��z��cU"�]	Y����GQ,L�AB���<��͂��S��l���9���MW�a�8Kj"�Ŧ=.�o���/J4�"G�9�6׊�d��Zt\`�7��S �̋H�g���uH+�8�Fmj}ǹ�1O����6a�L�����S�׉��䮤�^s3����&��#I �-Ė;.Q(��[Zokk�$���D�v�{:���5�RBz��2�Кu�ؓ'�B�7��� �+�L�qvt�|�Gt5�~��Jw���9������2�D�`��)� ۭK��H)ƫ�w�!�l��iG�������W�d�Gь{���sֲe����B�l^���6�-�F�U��uy�A�5Ae?�9⡳�ze�F^����|��3c�c�;���h��4��֖A��B(D���
]H�+L�	�F�̜X�!<�RW�� �ȡ~��.Uֲ�o��c�@bo�~M���  ��	=�:�vFHQ:���Y
���7%Z�@��L{���z�wT�6[\o��l���\�����k�дٕ��A3'Vz=��l�Z��h7"���~hi\5]Nw��릖�3E�%���ѭ��f�W��s���N�����mY6<l�P�����]�(T���ϜX�Ǆ���Cvz7�J�X��n����o�P�b�S�t�y���	�*�	�I��eG�u�bi��G8��ޓ���>O ��L?��?�����]9A�W��0���ro��l���5֘IM�|���~�V7R:ɰwx|��,[}΃yj�!�*�`�_���\;�[m�ئ�"�ɫ�:3:��is!��Q� Ex�L�X�a^��5ဇ�H+�χ�1���0��Cy]Ӥݥ�N�TT��
=�`n�B|YM;��~���b���$�ЃʴU"�����
V�#J*"�x~UE�3���{����T������8�����V��c�
��q�Z����]�-�%;�5�X�e�#�%�)�K/��K�+��م)!������}Ϻ���ݩ����#��n��\��[�b�BK��<J����}A��t�w�I#��"�\#���-ht�8�V�g�w��"vŻ�
|�A���t�۩����8��@�) ޶l��.NƉ���f��@���H-�|B��U��I-3�H�^���߃�F���G�S}?x-�g8���F�d��l���9�x��܇s��
[8��H~�i+��^�4m�5F$��{�6q��׵��~�[�߆3Fۊ��p$���������i��^�$��pEo��f=p�AU�峝�X��sc��$[QF�[�
����4��r>A�2:��X�~�a#}��p�ɱ�z���*0Nl�q��c��
����s0m�b����c _��U���
�G�E�dh��������u܋<�׭d[��$ߺ��~jRG��WCޝ]`a�C�D�>N(h!��v��*��Z��Hr׹q	�Q���g�\���S�u�¸)���Çq���̔��z���tql9��W�\ ��Uy��_��}&u;G��}S�6�n�~2�(��WVI1Z
6�A�-�����Fi�c��L�����(�"�:R�Ĭ�0��ڃ�X��Cם�)��B�,�]�nt��z�Si'=��&�E*����������S����?�&_�u%l��`(�j�;���f6k��� b�\&��Pl"6+)CID���|���i�g����<Ρ?���U�Af�R�K!�W��	���J4NY��/�8�bĩ�����"�	.�ގ���!�]���́�?�y#�#����S��#���.Ou�(�D�����1$�r��:�n�C��E�b�CK���t��Q�4�����<U S�d��S��"`�'������S��gZ�0�n�a	o���;3#�V��
7pi���9��ʏ ���ۛ� �G�;Ú�\n�n�h|Vj:�]�R���H�E�)<L���\�	����"n:&Tl�F��?娺6a)1_�s��,��QĠp�� ���}{�q��~
��������s��UR�D����u^
m �8Զs�+'3��{X�J��>5wu�->�k^�f�q�`H	LX�T�� z}� �D XU%V
?�!�K��b=BAa.�(,�Y"5�½|�^��z�9��L��=��.��`]v{V�$���cK �}#S�}Z;���Y@Y^6�.3>�c�n�q��͙��>�A��LB0�Lo�"oK�gG9�OܮG�69���n���&#+����ER~_��ob�I��JEբ�}ifqRI���AXrT= �x��h�P�S!�y���?���aT_%^zZ}'�F��E}�p�d �fpQL(k��Vy�S�H.�Ґ�η��C������a��1pl��Qm��.��'q�n<���W:��_��`���6$�88���&T�����o}��пS�(EO��>��� �^�+��:��2</Q����`��&��#U#��>VO��L�[��C���[�c������=V5�U7�`�璉㚺+T� �_՗��k�o�hU4[�H�����6H�{�E��_g��1B_z�,�>篪g,y�:��3\�0�K�i4�i� � �]54e8���J�~L��Y��![/��,B���ʈA*����婝�R��W��>U>9�k6�M�ˣ<�\�:�~I|��{M��k�i}tmS�@.v�܂FG0�C����J�f���"���֮�0@�py&�ljmnūK-�^�x/�<g��eF쳮j!����N�I�Tê�ew8��.OD��6�B�ͮS���	ayő`�o������5
";�b�!q��q��)پ�Z���۽���"�V5Qk�4l�7��W�I���F��T�\��Ϝ+@W���!d�@��@
y�0��������?s~�Xqpא�P?���<����0b�՟�z����Վ�/v�Y�vF�;��I�����|mO�o�+vZ��t���:G[Frq�^$�R�V�j�m����
[#`Lz�ܦ6��攵bM��`�&gp��@�.)�Fڝ��ɫH$���(E���L�:�<��җ��ɘSU(N�{<���{)%2���_;���4K,d P-(1�����Qw�nh�r�JJ�$K��YRUP��aK:~�!���n�I^���ڧ��i��u�)��Sa��N����W�� 7p�9�'G���F@�l�0e�4,_��Bf�J���K�bk�=�"	����Pg�}�ٌy��V�j�#)t
^-#������:N��z��[q{���'�����
sýY�$V�����ב*�&���m0ZA�"������9���hTM]��3�+ɝ�8����tAM?�xk�Q����s+�Vhz�h��Y�	�U*?mMH��6/}��z�4&}TZ�!�,�Y��}{�g�7dѾTq
����6�ǥ[Ajr�5�����Esǩ�M˺��~i�����y��QZj4��B��BY��hY8�ػNQ��,�����O�ڹ�4�� <�
��`b �^�|�{'���UЎS�Z;�d�"��a���B}.��t �<̓��5�/%å��)]�]�sl��.��|�}/�O��N�W����I\r������� ��UnZ��]fr�Ӎ�F��J��b	m=�*�(6�����*]����u� �L��Qf�]'	���}�����y�ӏ�=���gW�,�/<��|n����Rޓ��E ��換��T��5�	$�Z��tv��3G�'Yi�Rs��S�yпL��\��p�r�ȣ6���ŌBE�����|925H�2���;'~�]����? �q4�f��h�����ވ'`�BW�R�L�=]0 vV�Z��ԿkФ��2o���I�Mi ��iZZ����&�O;����ƒ_<�(R�:W�z�}9�,l|A���S|*ؤ���MtxF(>�rE؊]r���������n��o�D���Z��Ɛǌ��2�n��*�'s���$?���<��U#�)�S&�I�������1 ^H�T�]8�!Y�y��'Un�x�0D(���D�[��d!q�Q,u0�(����Q�%�pwix�l8��Ǭ���?��]*|��4aR��/��T�/	A%A_�L����z/���g�IB�-�}�m���e�֚q�[�)00k�CcLj��x� O�J�sͦN+�9"�O5 ��YmN �Nn��瑮+��2�=��r�?�.)���-	�P����a��(Q���Z��?lCc�p�%s���oe�j`A�����
�=+�v�԰O�{�>���|��O����AP��D��S6�	��Z��t�Y� �F6#'d%��uX��ݽ���PݢHr�JHt� ҘXrkӂr�� �MU���r�Vk��J.�j>>E��S�FɛjQr� @Oi:?Y�q�؟"��O�wW��/���|�ª.a�d*��CgHs�[0�����)�s]w�*��^O���G��y�|k:�2FO�����D��Ћ��v�zʡ��u��kL&����|U���%/Ƭ$�yS>���w�-L��ߤz��l^%��4� ��Z������yZÄQ��'T���իν��~�������
��Jg��(�ܻ��|g���_T��v��E�]e4���������`�-a�'n%l[fe>���z�ߧ ����!4􏯕Ɏ
�j�]��Z�JZp���2_�_���1faK�u���]��խ�O���;�q�'����k���9�Թ��lrdO�{��(�=��#�щ֋�Ũ����]�>)K���W�����Y�)��l�{�N=ǳ�u7۾o�υ���r�R9ܢ?��
��cK4
~	�q��6R�)ӎ@�#
�K����� ���P�|�D �z�ƈ�P�H�]��N"��E<�m�,�Y}��+��T�"����p�xU �$��좾w��U�hz�(U#Jn�0�L�K�V4�mz���3��&��>1�}^�5펶�,��D�ᝌ��z;��8"�S�~s�}� ��*���k]\�.��7q��;m>sm�ol��a�T�K1p�������ڇ���a����*4��kF0�ap6wmEt(F�����;19���?C����<��\�k�&Rp&2`���.� jUV�-����ӰY��ZRZ��|�<�u,��SΫW��Qˑ�ȵd�������+��N�[���<���-C������D\�%i�Y�E�r�Y��������X�F���;�_��?A+lk�3Vt��Cė��?f�[������'$s��!@)���.;��؞*�3/�wFF���]{DU�o������
yp���#��a7ݘ~�'��B=Y�O��N&���TRe��͆�x�{��JG'� �b8��/��u�P�Q�D橋_��BUj�\����u����i�w���/��},U&���c�F�������Q���T�s1*�g��|���iV�CV�:+��,����o�u�_(�Yt�2Nm�<�0,��7��ge�,4`:=U������|z��7��~B���M`u`����`�s�.RyD���5�N���Wt!"QI�W�i��❘1��Az���f�g�����,8v{ӕ��w�4.�`��^N&S����.�+�����0�ï���Y���}!��>S3^�'�>��yߟ{\6����pJV.�������Q��+�zd3�`zw��ǃ�z6+�[�'o0 tϑ�b��.��Lp{�0��jG�|t�n��:9B�@�u�8��k��#�n�2t�,��@,f�D����cun"��QV$4�{M�c�$N��^��&|�z�4�P�ĺǽލ�q)ѱnm��h��Pi��_<C&AT� T
����q��D�)]�$@=
H����~�йZ����ZJ�g���uXv��>��lr-��/����bUID�8h�Z�� !���L��>YX����{}Ck8��iȪ���:�x�rBƳ�)����z����;���}��xu$���Æz����5����w�j��O���`��WV+d^�J�*��5��b���)��0PD�1��l��������!�)n����&���j�%�q3wV�v|�#��s�[z�l��X39WX8O�K�w�����j����,9;�[sV�
p"��Cg}����]�ܓ��Y��ry�!2��Xa$)��+wfKG���.r�l!x�G,��!����O5�W� HX�Y Ȼ4�H��QK%����㞈Ʒ&�aEa���&���s�ڻQ���,e!z>O��F��>��7U@��%�����;�Lt�9�dI�+��:�����Z����M�GfY��;��Wk�^m��ժ�t�yM�;�&F����~��2�
�}����Eů��y��v�rN]��ڴFʌ
�wSD%�i��=�Y&�[g������V],���(�O�q���(�����!2!$�>C�T��L�~�)}:J���]�k��7Z>5!���e�̜��Bwd�JPe�9Eѩ}mZ�.��*n�Jx�f�����v�����?O��c�/�OKsd���i,~1� 뺨>i�l��j7�K5Q�]�70H]_�Y�� ���X�x�u�x�1Q�`��;�i(��XmWYz���[��aÊ>#I_3���A�
���<T��Mĩo��|�w�aco<R���)���Fs���<���b��**'�ء1���o>�����H�k�!ߘ�u�n:���� G�ǞN��Ѥ����[4����a���+�G@���^��F�#����Y�
%���S�L��*�>�sj@P-W�H8��0�?��C6�BO���˃8h�y�ol���3]N����E�u�2.��"-�i^�2s�A�.5����$v���I4fT�yό��n`�6M6�> ����~J�Ĺv�G~I�؜�p�SeB	G����U(��D�M;z Ir����3�ϸs��+��?!^�H�����c�\���.T��u�x������o}��J���� B�f{X��b2�c9[f�X���e��ر#{����",>��g	]D�&�>.���EM�}-Jp�U�
oA5w;`Mֲ ��4����e��L�ߪ"���%Q��C�Q;�ɍ�t���M�U�0K�TZ�L�D���Lv[����r�b�>��|�9J�c8,QO�£���Vc��M������|a�vPZ0j�q,&�,�e.�R�w���V�+��氢p�n��޼2�]b�&���
�Fg�`{0>������1u���YcW?嬒�a�,9����/�YhS����rv�t��������ya�ʀX
)n�,!-�:��X�R]��^���>���Ju��<1���ג���H���P=�4�x�ВH��3�]=������S���R����)�Qӭ>X�
���J]�C�@
�k�G�{DY"���/����I�����֎�7����C���RY�-�^8~*�OEX�U�KՃIt[O]$�7<����X�uq�-��Mc�������<�S�y<X�بp���gp&`3%��
�e�zr���Ƒ�i���s)�П��f�%5�x�u���]�K �aI���Y [h
�Js�+sL���Ś<�E�8`�lw���C����h$�n�⢀e�¼3�3����/�2�`C�NL7� �^L�]��\��/�
��J#d�H�u���2+�z��{B�-�-���H֏V���.30�s���֔	��G�8*`���I?���vu\ �2N�c�:b��wEU��rJ-��v��0]�F8g�G35_�����"����8��)T0<"{���G���ũ���q@�� ���`:��a.�{��E6���ok��(��7��Rqn�&��OZ��.��lY\8m��9p3i�Ҋj���~�2Ϯ^���!t������G!�gŎ�*�Q��ʽs: �7h�O���Y��Hy:I� �}Ϥf��U��b�^z��R_��H�U��ϑ��Y��$��T�$��X}VB�d@}ǩ9�|RO��6�#��������y�2%!�E����~�Q���l�9�]u��V~�Ǫ|��JA���6f&���j�{s
�>!�lx��BB]3l5Q�� 7Vx|��k �+����;B� �ӛZt�N~�C�	1��"�5غw
�����gu��]����x�
:?g}(��{n @r|PJ�M��X�A�Nx�n�8�?�}t�,���x��>#����Z��qd�dֈ	����0I�%��&vʞ��4^�c��5h����1��Z8�e�zH3Afn㬾&x�`�p�,�Iq�6N�y�}Cc[�1��d����F����SMm�Q�����^(� ���=��
�Tw��M��(u+��p��U�UȌ:����͊��F	��wF��{��i~�8�~�F��M:��|Z�2z�N�S��z�I~17���d� �|�ʣ<֡�@�u���
�[R!�q_{����j�3���6�?"c�(g�!"Ǖ�[!�-jv2��؞	����/�9�%ྪ�`ӂ7m����R�ApraS�2Q������!����_��i:D����}�Nꠢ�&�6�N?�=}mM��T�x��RDpX{ ��k򺡚9��Y��WE~h��/�TgNW�3٪�gZ�Ąc�=�W��]��8���qL�����Mp�~[�=`��l+����O�ل�򈸛=�IZR��T�|t�:ˋo�p�x=0'���P�E���2��u�"�S�گP4�i:��@�H�SQz��%�_<ΡYiS^d�	��c�)ڮ�$���V�p�]�@���