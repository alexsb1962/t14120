��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?���e�F��M#�=
i��
�l��~,�!`t[Ҁ%()�֪�Ч'����gF�ڨ��̌Xs[��'	K쏏�͑��ðƕD����FG�y���]�i~�t�W{�1,���^x�шP�L�X��ka�Lg#i�]'��r�/�rt$��)�}<���a�g��2;Ʊ���傚��<����z,⸍Ӷ4ኗG�ƀ����8�������԰�s��2Y	h;�:����'_�*��>	J����)�E5�t���xY����-c�f���R��N�ƥ}��QM�52��/籼��|�$p`�9�8�3�`��c��IW��լG���@�֎�g�Ee�(p/�o�<�1�M&l9(�Nm7�A�##yC��n1�?�q���z,C�Kq�5�'Z�ӓzn��{��kM�� �O���ձ��~�H��N�Nˣ��ܹ\[�:*9s�sQ�A:��BFI�1]Y�6(��pj�� bbr��Z �����>�gc"��UM��g���m�˽,�T�,�K��KR���>���M�*�KW"r>*���I@"��u�D_A{{n*�ti��đ�\����q�,}�c��s�dX%l��N�-�K�AK�:��<Y����X��t_��C8�lȭHI��^�k�ܖGCcZ.$�$n��p�_s�'����]���81H�k�@Ƀ�H�sѢW-׸�x�-/ a�"���%�
�n����b;Z�R�����}�l��~��)�>�X;�<5%�Q׎����oa�S�?�R$��a]	�Y �H��[Q�qp����U�7gD�=ߖ
,}��;�ҵ�G�Vh�g>!0����kå�p�iP�&����W7�5}vC!o�ġ�^}M�>���n_�n�bYZ���_��\�u��7�˥fKU�m�Qp���F%;:�E'4*á����e����W�軣K�쩹�sDI>�T������!'���u��(6��{��3T(n�Y]\6a����s�s	G�޼�Ͷr�z$��wP���I|~�HrfFtF|툿�y��
����1�i�`<���Z���ň:��jqv�DS^�3-�Ĺ֕�F�K�#�N�2�B{��-j�H�7�&�)������ɯ}�\=a�ϋYw�`�`n>�xۋ���hԽ!���eL-�:�M�j��"�kɪ���B�+3��2�t�{��@rG.�{��Ͻc�/V��7��A@� �y'��Ӟ�
iΙX�[lR`�%������rK�:�+A��^�mOl��)7
Ԫ�!�5v���{���S�w]w�{yȟäL�S����tU"��U�3���%-���fd�V�y�5��΢a �Jk���I�=|�����+
�N�e>���Y�%��\��p#~��ys6�;��ҝD�e\ �'l���0��ano$��9��.�!.�xʘ�=�Z��a�߆*�Z��_��?9��g*��c���a���z�ET5�*���c���ڴ�G�*b�<!#�-���sԯ�; � )���0�PA�놣�F��J ��O �1�H���D.1uO޲�������v(V�E��g���0,���E����}1����n�@���n�i v�L�$�Q�Q-����݅�D��<K�������gX� ���N� ϗǌY1ܾ�n�b�v�].s3��Yu��y�}�������7r�����L|�����0C��,�oiuL�͗��.��gx���滲n�bf���ߥg�l3�g24�ٹךB4K��>��>�p��"�u| Ŝ����Ik3�L;�St���o8G6p��ȋ�n^k��E�y��#�u�<5����U�
߷(Jmt�m�s�������6��ڃ�LH�zrK%���>���T�����U#Ji�@e��' ��*��,��U�ȹms]:�@"M[���6���K*�!s9Kz��)����4�m)4.�!2E�a�'��喬;7���-*.�de{�i��~�\����X��~i�SP�hfo:�����BnT���9�X	x�FN�v��k�V/X
�	{�#�f^|'˚}����;��.=Jo�,N~Ql��3S=�Ԍ�C�M�������c��-?���,�&o�*(ɸj���wu!�s�]c,�z ����<��]�[x�;�t�˫�K@��_T}R]�ιKdר/
�9%���~�"�^��*u�דK�1���]��x�2�P&�/]�W	��8�����L�ͩk�yT2���=ľ�gҾ_�)Ǧ�Ύ#1���_����R+E�"��v����d�5JW�?^@A�܍D��<��k��$�m�?&�E���-w��b��s��E��񝷑��0���R��#��s�hDA�v��|�蒬V����)��^�˓��=�EƉ3;z�A���!Hm\[p�r'�H2$bїc{H�����nR�T��RC`�7���q�l�d���N�s���NI��sy�?	���y���)vG�)G��%ka�yw�m�l|��U*����l�?�ۢ���m=��Ҝq�Q��Ü�@]��Qw�n�_�x�� G���ٖ�	�|�I����"�/�R�Y �n�xXtΉ{
r��~�rc�����v&T���g$|5N!ƅ������ǒC���<�g��5��*Uٛ�H-[�]�"��S�%��O��E��kY�����sh��_��u��]��խ�n1��8h*�1�&B�.�7���Y;Ա}�z=����a�l��cM��'^�o��6�ߙ!TYp%������[��lւˡ��gA~x��*�:����S�;�/�
�c�M !J)�_����.�@��_U+t�H�n��#�j�s7�'�S�D�k-���D'�_��YM�l��������äfE�"�c|F>��/D[�E����4���H ��	��'�%/��;n/\�[�ou����;�%�2��"!�G�3�_aUx ��j�[b�q�B�D�����/s�H�m�Z��6mA�R+�W��4����6I_�!��k1��eU
?��p+��RV��P+�a������"ao~rq"�"�-�&f�ч�Jy�7�>�u����,�V�����-��l���h��eDV�{�����Y�(:��%6	H>�
[pV�ߣN�`���Oy5;R�)ڤ�=:J��Y�HR�_,Ls�('3�a7�+Km�����
u`(�6�}�as�&Q`]M2S����{VD����5�5H��y����o^G̢'��"t��Pܸ� ������^���법�џN�za�t�"��~`l6b>��X�.��I��J�X�
�j#9��X!���Z>+Z�а���� ��o��D��q�+J��&v�Je�tt�nl�i��p����+�G�m.��SM����z�:c� k��� �S��ћ;�;J2�~z_Z�:'p̔��@�%)��l�zȆ�w�4}	��ҿ1�V�+�7aT�����w�H�uqЫ����N�>��bM����,��<AUS��㆛���on8a��]y֨�-��G���ۆ>!��c���i0!u>�+������.�o�ӡ�FD�?��U�_���]}�E�Q=�ѭ;+��Rs>Fv(�D�י.��"��*-�$�Zz��@\���r���J������ڝ�2y�?�ׁr� p{�S6��޽��f�>^��V��M{����k��;�pi3	�=����dP�s����`�mQq6("D&58�����.���FdC@�����|U|i�ByG�m٨j�$������2>9��h�f��q\�*T�az1b�A�y�s��E���+'�G��DBz1g��K4Ӈ��C[�2,H�	lAu��h|�wùK�����C�n�/z���-Űg�~:�=�E�;d�ۇ�Tx:a��f�dq(�chV(� }�C�[�ȅ,�V'�(~4ۺ/���4�d�|���O:�HI?Qe�+;��7�-d:v�k�A����y����*�f���%���cO��-�އ���{��:J�S$):���3 ��[Ķ���7��V�ļ��fi�Xr�]�C��v�a�����ݝX���wg��xI�z!���U�-�ae8� �%���M�t�#T�mO���X`J�pi�M�\�?�b5�?hI����Qz�J]�Q�X�%􎚦�RPw>��<�o=8���賘�O���d���xig�%.�qe|�V��RM+�lU�m�0sa���G�k
��E�}G#�[��?��m��KJ�ӱiH�n6��Z��#�%=ڌGt<�Q}Ҳ��)��!�a�y�lf�{��m��}&�N;��\Qc֝^�}���y�'��\#��+-{sڼm|��`3���H��쒼���X#I�r�b#sbL��I�-�^��?�X(���!;�Tǜt�Ư��F!�@�%��:����Ƹ��� �����Mnv�dZ�F��-���`v�_
c=ў�B#U��óː���%��E�ORNb���qz!uͺ��ŀ���֙��OX�j��v!���͠�>Vu��"+����x#����p� ڹ�M�.wv?�F�F!c$�>sN�=!��}n-k��=0_p�i��J�0��:BQ�d���CH��}o���eYֺ�l�%�
7�Qo��c��q;��E�R��e
�U�b���
B���	�=a�2�>����� !�I�P~YLn$��faS3+;��Y5&$��I�X�l���茱3t�c]ֻ��2�f�&2��� ����r�~�f]ʝ$�}̈́V�{tBI�0�ET:ڇ ~)5������7p)���2�;U\�rC_N����3����~�*ܟx� �8����B����L�X��9��
!I�R�_�� �v���e�c�*��W/��P/~���,[�Kې��v+��3h�c������n�G��&������Z�j7�"M��1���iR��rI�p����2��S`���Z��l�D#H��� ��T�5��
{"ΏP�o�W?��/�[z�?�@vM*�.��tJ/��U��`F����G����h����,�U�"��u����v?�������}��A��$����n;ԼW���~8�Zn2wG��`bL��Ę�G��䘻f]���K��|ﾚ��^���4��֥��e�a��4`}��]�[���cFg���dɅ޲�zXj�t8��%;[����Qʅ��￬Zn����\d����u�nUc���3{�����g/������\�c���|�����A9>}l+�C�u5E#�0Z�P�=3�g���e�X�]����E���kYi�n�5E�F����jn��cBr�'��l㣛U/��7��_ҏ�j�5g�ʎc�K9��Q������,�=���}]��!�\�$><�}yg�<�%�3�Y[[�o�1=��6�
l��1�}ϴ��k����	�*�%�`J�C��`��%r�J�*ZU���(S��yԾ/�i��	';Q�0G{��R1��<&��X�t�in���3�hO�53a [�խ�!:��"��DN9I�J{ŧk�����r_�5�비����ψ6�?��S��u�I�\�4,��p�v���7+������]F(��K��r7i5����!�E����eDG�R�U�J}P.,��Oڒ�-��$��1l%J}�l��Sn#�>�,|�f��F%�»e8l^0\��h$�^�WN��ڃ6�������)Ode�(����������.�=!���͖�[
�/%d�����H�)7��]��FV8��7��s)�b�vѫ�����'�����e����h���TƈiD��c��MHʅ�{���W�NN�u�u-TC��>����{$1
;�z�jaE�P��x7Ҍ L̂���j��ȴA�B����|3�L��p�=����Z3��, [��x��w���7�N�N�n��p@�J�5�;j��j��*L����x`��lG���$�Y�6T	jw�py�_竹y��Y�%� �v�p*9�Z]��b��u\F`xƐ�e��=��b���	~k9�8\W5�� ���1~d�쩟�±�nƖ�v��Qt�(��%�6�c�X�i�������,�Y3(х�Q���p���b���X��+0���߱�6G@\,��D�����J��ʮxC�U�O9�k�L1��`�1��ڲ�}��ۣE6������S�>*G��
ܕD������M��5������W�ly!���������>Ko6^2ny�,�܎�����ɐ����D��FR���Ci� K���D��S��뇈�c�QS��K4������LǒƐ�&��{{_�L
]�I�R�?1B�bQ-�������a_���֪�﫽�u.�p��rN}й���i{���I��^�{�D��<�F�,\�T:E���״n@ߴ�S�!-o�g/�Q��U:0�+&8P��=:��Cl(g�X�j~U�����i(?smV���mF�VG�
��<�V�:jS���1&i��=�o@~��<iO������G���-VVe�ZS����*!u�v��
g�D�=��Ҳr�	s��c�9^��\�G{a��GV�cfJ���t�P���| ��u�����Ixc���J/��t��+Ƕ�S�k'
��n�j�s�*¢�\:V2��L6�[fzL��3*�z�%*�m7��2��e:� Xp�w$���x����x6�p1c�4�V���.��"Ly�) �^���J�N�"��-*1=W䧓tk�Qq&*�B[И�����uhV���#��ÿ�5줉=�%���Tj���� h��\����*�-L�fБ#���lD�*�z���z�U� q����} VK
�P{9����0Q���J���S53��w� q��/^G¯m���CT�{D	��r�6:&�?�pF �H�ݠ����V�_�'~D��G��%r��$���8#�;����#���zF±�][z�)�~(�Ð��Ԧޮ���`���61D����(ԩ��-�b��o��_/�?'/�r��.��.�ɠ�#;(�1i���"
|TP�i)N�脿SX����V�*���-������$M�x?P��/~C�3rC"맙Lj�¼�-�R��ў���\��!��{&���ʉL�X���>��Nx�\��X}ߍ��A�R4{�h��d�*��dG �}4���`^Fz�M��;jnp�BqcyҊkE x6��w��V��S���x�O!�C����hd��}��ǵQV���� ���{\y�@w8�?���y�G6����TS�þ���.��=�.C~`ઉ��V4F��mT��\u�!y�̙o� 6���>��|II���	?�Ps�C<�IQ�A{j��_{8 V�������.��{�� S�J�VD�@�����8����u�e��TY�C]@�K����.�w'�>���!{]·�H�J�'i(�c���h��&݈�<��}�H����g�e;)k��&bnaЛ�R5��$�����M�n5�7MaL��5�K픙f�b��G�b�F�©2$]҆P�5�B�ݗ(&���̵��&�N�չ�0xk��+��58�o�B�C,G����$�4��K�L(�E�S43�E9��_�VD��	��Y� 8
l=���XON�D����c�t�[��b~o�b���ߚ ��Z������|*��l�lQ�a�D�+��bQ�gGY��H]ȍ�rf�%:������q�}AwA4����;�c����RvU��z?E�7�����i�€y7��l>��mlx�+��Q�bKj��d��k/�d�fƤ�9C1�d:��Xk���XO��J� ��*�u ����6X�A�U쭘Xa�%��=��MUq����a�U#Yj2���ѭcik��baa�F���.up7Y	�i���1��m	�A�r�r�j�|��2d�і�"H�WU�[$2��Sk�wCl=l��V�}{��I�n,�c�����*\����%�X���+�F�h/�т/�!A��7�~y��n��ZXr��ʠ����$ydMpM�P�H��-�-��ܠ��N��k�a���	)��A+Ʃ�p��槾#�a���Ex8��#��B6�������c�v��'���S԰�ԯC0���P?�CbH�����^��F�L���"�\e�$�5"�/�Yd��a�,�P�z��Ҡ�1�#-�"�!P�"��f�f�k��B����$�Ae/�o0PO�6��E���%�<�#f��pD��@�����
�+S�����M+9&�ww��˟��ow�`^=�	�0�'��Q�!h�b���4a�qR+cH�(�F��.��P� �@i|�
��^?	m��ʥ:��ce<������n?�����U���,�-N����hat��҈��&�g�j������^�ƴꥆ(�\�5�17��y$�>����0�ʝֽ,�b���`��|<��|�O���(���v�B�5ߟG�ޔr�d���P����ȧA��9j2S��-h@��Dc~٬B(�-m���&_9=Ȩ(�!����tG�䄈s"u�����=[��R\U<�I��P��)2�\Ex���k�p2�O�{�����+"��d�z�k��9?�sa��0�\��kA����n���?N?#U�c�wJɽP�Ahnb�	�~�P��J�o��mu������z;Jɟm?V�x��c�<0vB��fx�T"|DK��|�P����/p&���#���}��(�(h�c{FxP�Cg8�˸75Bq�����ҦcԠ[�\d��<�q�h�ԥ��E�����A��#�o��5���ſk�^�H��3Ux���zEɋ��K�R6���XR�әR�����|��U����^~�vͱ1�����,��T��Z���@?��ec�͘�7���9�S2�633og�GLG^3��.o�FN�@W�����;��ϒTm�q=�:�3x�/�b�<k�	�q!z�&LdɔɯPW��TЗK᭦ԏ�mz}r�W�j�/7ڊ5f%����݋�e�ı�ŧ�����t�|����_�;�}ёy��Vu�]����Q �W��aC�yX��*�'T)�qC����p Z&�^DxsFMh0��hԬ��g1�Ǻ}��{�lK����r7T6)�l�	�s���-(��"��LU�	Q�..!�d�_߮��Z9'���a�`��Y���N��Qw�J���0�Nd�/Z��ᾡ�c����Bd?Br�|�pq�".�soTU7�ڢ�ظ5Y�֧�RjT����*�G��3��R�V/C8%7d&}B����3�����W��b\�E4�}��4���/��#W�NC��E40���H��uf� �R4����!��s��`������\�q].�~A\�����v��s`=ntz���c�Y�:|��	}#|��JL9U��Α	v��rt����nR������͟LBecL883�Y�(q�{��[Š��{�BT�]Ⱥp�C�����y�9<=�Fc�y-��h�����̸:�@?�v�10��4�!��wp�9�Gw�M|��[<�2�8�(��TP��E�=T=!J��=Ҫ[�����d��ҫB;qfZm�}�d;�}n��Ҍ,{ɣ�2ߧ�� dL�џ�S;E5yB�uzQ������?���b'z��=�d�z���`<��.`46��n�=���q�偧�an�9e���nv�x6�JR�[���2���x��} �{A��A+��7���L��E+����}��9��CM�;_: ea�Hm{a7e��8s���$�ZX�p�_�u��Eh�K%��׽�M!'���EG�gO�l�.a�rf5'��&(�A(�}�S&���xW8�;>�*���&{�X�eMT�'��P�O�PMLFi'�z[�A�M���cu�VĢ������y<�2%a���i6�!'��&Q����L��s��s2 ���-�+X�pp��C&�K�3;��m^�*=�8R��t4P��gQ���� 2Z1C𷿣[cln�-�k:>�,Ϙ2�X??ϡ�i��Ң֮L�F7/�C_D���5���~a�R����%�5��s�ߙ���9�X�4/��������y���#A�i�uG�j�~��Y2d� &�z�vu�A���N�F�����_�u��H��F��k��Y4U[;m��H�>��K�q~ߛ 'Fz��Z����0CJ�=<Tc�&޴p�N��/ť0���/�҇M�w۵����:��7��%���i�'1EUA���9lI��w1<�k��*͗h���l�i�Sw����:=޴�'�݊��`�.�=��g;����S�r��Q𨹮���a���?AG�#�sP[%͛H�RK�EI͜ZB��A1�3����oH@�/� �f��	S�B_d?]'�����M�9�0��Z��@�22�#�����mÒ+�L��A�ub��?	��I֥<B��z3�S;����q�B/J�'�=f��wBkL���؃�{&c
8,�Ё��MR�k����#1d4����Y4.�8��Cf��Ө�J9ʭϸa��S�4��S�|��q�q(���?��;��$ĩ����]k���y�#h�n�4�R�D��)qw�I��>�M��f�K	Y�}C�\�^FPc��O��~��������c��L���e;#|*Ȱ��^��킔s03�k���YZ|@��c�g��@��]�B|b}¥p�����!n7�_�9Ҟ��: )�r"���l����P%/A�.
�Q�4��sQ����'DL�,D<ruh���k�� e<�=_���AO���͠����M���e��g<����E���v��c�WI��{i_�lhS�������Dq7͊��`cm�n��*6-B�,4���.��M4�s��z�t���z��kpxȵ����j�OR��[2Ѹ�iG ��76v�N��3��N�/x�$gyj������"|�*���zR��*�,àOL�m^G)c	4�6���d�/� ���$&u��sz	��''�ZS	�yYo�+pƪ�\�����H�M�Gv�<~�y�ż��S�����0C�-��~���}q�a�#�k\�Q�������K��,�\`��񍖓yr�gr��b�E�)�.��k�wC�4T��M��M�R��]7Zy�l�����hu�Ж�oP>�Ҏ�6���� (�&��<
7���G=���3��������k���3	�b�nFE��ޣ^�F�������S�&�l����@r��z�'���ҋh!���~�Fb��#I0�x����1�)qb�D�����)^��Z�>?|���-R7MQT�Sf;�8��д��M3Λ��7Z������S��+3��>���d����:�{�__z	��d� �^M}Ay�Xz�K
�|�
�=o�b��䋇��5�h�ژ����2Q�]��Z9Љ��/����T��A��	�m�ǧ��}���6,�1r��1$���hvq�ַz�p�#�7[�&,����7�>2�d u�Z�����UgR
�YW�ҥ�N�#�t�N������&K�k�W��o�*�����B�=���#0�%8kV�J�%�8�i H�6*GZ^��c�O��|����0� ���x�Fa����(/��c���V���i%�\`���tE�,
t� ��j6h�|.%Z�B�L@��7�[�/���J�DᚲN��g�b�!��mw���q��9���e��#�
P�:�\�-f'���C���"��ln��*kd.g�|��2����#��ؠ��n�)XLU�� ~��e�3��N$��د̅8�or��m���2�c�*	H.�s>�ܦ���ńͽ^UV���-�L/T��|�h΂C6Àg;8�����`�Z��-���u�{�5��R�'Ҭ��2������to�`��7Q�I9;ʄ�%��o��!���RU�z�C;bW��[��ص�k�>mܕX[��P��o,�
�����[��b8� �R0"ݾbN�CU���,��|no�5n��C�W�f�]8�PȜT%��D!q�C�_��$�(�S@f���]�THW�����͹�ג�B To�_��i�pYd�Ƞ�"�箐�B�7}�!g����|�oe6�IW)r`�V,�Xz%�p���ZއMh����F��=���`#����G�j��"�Z�����e������*w���a�ׇ�7�jBm[ZUWb�Ka�c������<��.���
K�e
E���X�
��u��6��y㧃5�-�����D�_{Z���_`ko);�]hxV�ijY���N�� n���.(��9i���;jp�c��Y�����ꆹ�a盖F�۵������k+�4)�GR{v�y-���u����eFg[|����5C�,�~[@��T�����^3���X@�3y��`��=����y��{p�=�J1N�����A���`�|��iPN�}!Xn�b�VG]y{�6��V�����O�SJ~ҟ��B��Ĝ��T�V�1iR��@��ړj���3��ZAwf��F�Ǣ��Q����5���$o -;�&�C�k|���\n�҃F.���Mz
@���l�8��/�J.V�3�;��Ǉ��B�b+��Y��yv�8��, �.\a��#f��z����,x�FE�!x��5}�yHљ]���E�����N�'f=Xİ���XR ���˜���r<+��A�0wR��5��Fe��q>��,�
�"����������1��T΋�5�~�พz�c�ɻ����8�ZZDOkOw��-"����N���L�d�F�_��Ki8��"��5�}z�!KǄ��y#�禓%��Y�����;|���,�Mb�4�7��g�*ŲeG�o3��SC� ��v�U>�F_��� ����,5�����!X�E�ju̎��E��������h���݌�ܪ�6�7�����1e˒��N=B��b�8O�����&��=Ӈd�:B���EKz�_�ye@:�
�� �M�U9�;��Y�\��/�_K^h�K
�$������{���k"|v6g�0�\1~��}"{�2�����p�?k�H8����z߲�="(�
���/S��ad��>�\,cP���`r[^����oNK�f�]��5Ŋ�7�w�<�m�K��9�詷�~':;��Y��v��'͂dmr��A����D50�V)��G�-پg)J�׷(�ۆn�����i"�h��ܠ�ԇ��I��JX�`k�z���N��+�l�ڰM���)w�=�_�n�|�嬫�6]���M���	�ߣˑ��D뽨Z�$��_� X�P����s@�Y�Ԋ��އ9Nx� ˍ��aӧE].b��>��7�l�,��1s}
綬�
S�)�ܨ�}��dA�=���m�噢I�
ܡ�r&Hf�TI{���� q�U��ز��|�a�rtT}�[م�(h*�����B���`��t��~\���.R�WA�x���O�J�.B��	�U��<y_#���C�?8IA�\�E�K��v2Hg�*��ֲ����-i枣�κ�I޼P����TG��:̥��2�����ϗ�sP7�9k#��8M�����'�� 5���ћ�� �t6b��8ψ9�OL!�Su�E�����O��?��D3-U�7U}���睌�@��ɥoid�����M5�?p:��x,�XjR�	Q�M��Ϸ	�a���D#��(�l�gY��>��YF�� \
�p��I�gR�Pf%ʥ�ԗ�.����#���}$�iY:c��S>��L,��l���^œ����+Z�GG�Ga��=�����xǸ��ˇ��Ҍ� �Q�2V����4|k��TS�����X�4���I�����n����	�]� P6��.�P��G{}ٟ���&�;>�q�Rc�)_��rfM4�c�b^z^<g(㙗��ɞ��4��tHA��Xʒ����.��qT?�� ����j΃�Y���<4Z��65iSEȰ�]Th<G:fH(3���N�x5��[���E)ý�{)�C�,j�=7��h�
�C&-���О�\;�w �� "�C��.ƚ�#��˲S�!{��8:/�`ѡ>���S�o#>�E���m��a�*�yS�z��z8��Ç�p��iIuS���0�d��ɝ%Z�j��z�|5�+*VSd��#&��Dȋc�4�������A��סz��C@&�	-գ~�߸��
"f%�gMq��1S���!_��"/5��_�!��)��g�oܯ͘�~^�}p�QL��N�I�1<�o�a�ج������J3��|����@uX;���}y�͏M_� �(��}��D"������L��J͑��mǘB%��7=���=�1t�0#e�K��?��jjA�X�'���1��h�S6�+�o#c�XB*;���b���4�.K���G�8�!��ׁ�Y� G.'�9C�9Nx�w5mGR��@��.Y!�
KD�D4��L(F�� R(���(�tQ��n�T#�{�f�J��t���-������Y !D�n0��:PӲ]6�`L�Z6������jm�¼M��(.��Cܮ]�sxv���Ԕi���٠��2�T�����+`��㈐Je����y�{����f_�d�U=�Ơ��#{z�^.ĻC�4ē�W��	��ã����������Pd���f(|mm��db8��HD������"{�e5&s�0���M��E�,�e'(��F�6��(N�,���%)�������Og��!��复*)��N*WnrO��v��
+a^��*<jq���G���S|/h���%'p�Ѯ߱���*m��/�P����W��fȶ��E�ªu�_H�*
���<��v�g�H��p9� ��9���i�=�,I�O`G^��PU�k��3����u����D?_�����<<�zZ�RK�j�Jcܻ[*����Py�wB�Y�J��G����� Dre�]@���t��{�7��]\�q�8S���#덄'� ����F��W��[߁�o\󱋗����zC�����1$z�������������ʋ��W���`��b��Ϸ5��`H���Щ�zR<��*f���=؈:����3�|#Q��4~��
x�#a�bv�ʜ�� �o�1;�54C�\��]�q�1HJ͟�;|���3z��&$ޡ�� �S���2��L�]يQ���ś��h����8�U+�¾c˪2o�pc]���-�"/ɱU+ޢ����qȶ#�Y�&�HAY�ܣ��W����{W�� f��X����V�"�S�������;� <�e[�� �<���s(��<��G%��TU'�O���b�p�} ��x�^P�WLU��.(c��(��C�¾T����g�-�-�K�CX��%��ˤ��Ԧ�]��$+���{#�O�>w�����59��Q1wou�(�?'c� �B
Hn.j��$MQ�&��"H�24�x3�V��Z\�Ni����{z�u�킊]7��/��r�Z��S���I��d��;���Y��V��G��ԟn~E��0d(h�w&Rג��쳩�۠A3kD���a�0���A
x��A��1w����yq���� ��"�A���,��Gi����wJ,_kg�v֥��[�ܐ���|��5tM����1Eu`G�Ŵ���{�rj����h_�iVz@��LC8a�2uQ�gy��+6Tۧ���^�ݢ;�׶D��5sRVs��xO��W!BgS�c�uγ�_�ew�N�]��5���I��ԥa���E�Ӻ��NO����>��f�H!�P(��#9O��%�pC�e�\�iʎ�Ƹf�,�qkǊ�S %�{�i��`+����۔��$�X�"��#�:�^�B�����ßt���;S�`���7'�H��/MDwD��.���/�J�9���t�Yۺ-�P+���v���\����+j9���L�K)���a=�!�MB��f�D(郻1!�̝������O���hz��z���-1�"	�/̀�Β��5)��l�"{��f l�	��;j���q�'TK�� �ʛ2�M�b֘�<��{;�2�����%��'I�=L �!�%c��N��_���
�(�p�FD�nU�V���[�,��1&�ӓ���-�d���Agl!�Y`�w#@���Q?��G����I�CpW��7��!Rɀv�-�y&dc�$Tg��*p<~{�|�I�L��	�}���I$��/c՞���r%�H�"���ɤ�C��q�D�ܠ��In�!�wY�(�S�{cX�$�b�^�l���Ok~�5�Z A��
g�3�S���}�x�lVZK�ظs)���"����$�a�������\���[�$�o��in�S9����ji���g�>�T������:��{�a�b�̓�Pݚ`�/�Du�
�w����Z8N��aP&i�V�2�"�s�#!��%�:�x��t[��+b��W16�K$����,l���y�v�b���c�:L�Dʴ���ȅ����+���I���L݆�p������CLm���OOO=ۋh�>DIN2Y�~����6�<�',��`-L�t��к�B��OC׀)�we�+�CH q[��l����f/��i�e�Хqi�F��}J*&cb����}���Mk\�����ag�g�g�ȕ,�(�����+~���N�g��(��i��I�`�bQ\��G���}��ܵ�=s���pO���S ���ָv�=�8i!��R�>X��-�d~��;Op���>���2 �J��l�M�����*)'N�ڱ���Z0�}A��R\衴�2�WR� Y��ބ?�^�+qY� O����]�F!q(�l�4�??�����K�Nݫ�$���Ⱦқs�gܕ�zk�� �gϯ�9���Y4�X=���`.�+��F��\Ty�61Z��v e��5�"�^v�|�i�������3��´w�?�G�#�؀d]���d�
�=!?q�4s���^.'�Κ�R�¨k�3gx�W>���IA�1�I}-ǄW[�b�=]�����b�[
����Q3~��v�2qm��@��@1~��Ibg^f��OS㈏LH��u톟�q�W���d,VZ:�c��j��Nq,@������`a�)Ţ���^�z�M�0�Ll��3zT$��q>���`1���#@����sֽ��iM�c�ۡ6����[aWY����s�d�z�6������"�)�¤Rk�cn�;�9��.R�����+�A�Q������ȼ54������4��3q�xE�m�3�>F�4�b��)௫:�F��D&P�!&mi�:-t8�A���p��� ���1us3�17S�D$�q��*9��j�H�c�3��6�e�(�CgH@���|	~��
���_?���{c�à����TjY�wI\T�4�p_�7�	��f�O���)���|�8����u��SG��4���0Mܶ1�#�B���F�d��4��.Bo�l P��/A�8�J��q�S9W�$r��/��2������u[�v��zNZ���p��a��Uv>�fO$|4f�u}k+GQ-��6b�Uڔ-����9�E�-^���0�h�p�����(ٚ� V�ڔ�)W&�d��zd�J�S��Vo+u@DiAXEr�A���r���������
����h�?v�^���� J��c10m��W�{S�/���'[q	j�x����:�B�Gƥ���`��M���D�0iA3����Q��H�4$��1�Rqt�\���b�C�V��C���$'�D��0��9��`���4;�E���� 9_3\1\�3]�2c�_"�4Ɯ3�9*DR���o�������Ά�o4�tܣ^aW�|�V���}�͑y�Y∻xVnPN�\vb�Br�!�	�.�m���y�����;��,�BY�܇Aa�+��$q�$���9DW�]�RF�Ͷ��{Wm���6Os��O.0���)!��7I�����0]<���ʋ�\����AU{�鄬���R��x���+�bvR��o�zٌV oZ��p��ڞ�
���]?�;��鶣�a�+,#�B؀�sV�:(N7Հ��e0��*$S}I�w��3�5s���7���̄ύ(�g�4Φ���J���!?�S}d͇���(� Iٞ�`��b�k~�D�;:��Տ�:�6��O��������H{�-��p���y�f�	m�`�Sĭ�:A.���X�A�E'��њ���#��Cޱݩ5�����PEC��&���2VX'\@�W�40wm��e5E��y���h�*[&%D�)k�p��O��;�z0ĥw���	������UN���!���
?3����=ִ��<C��N�o>P)g[:,ERΫD]���/�-*�"�l>���7����*X��dM�R��{�R�n�~��y\��>w��]���	zr�Fd���P��r_Y�
���4�O�;����*wI�T�W^����0{�[Az���V	%AJӃ��i�ֵ~��L�$��TM	��(�O-	��������5�iu
f{������AZ!����4V�G�-��݆eZ�B���d7���������kpb�h[��S�w1�����a��V�
�X.�M6���p�S'})��w�V8�s�&��i~|(��jM�g�ǔ�R�#o1��Xy�-��@G�Sq���HƵ�{O��;uج-��̠��8cnT��𱭫.�FdD��A�Tjt���"4�/����?x�JTF&gء]a��L"=���͹pV��[ioYv$R%O�`U���0��nUy�~q�q2J�6������>(t!���W�oB|�ǉ��~��+TZ��aa0H���q�]l��������&�"fj�;>��G/a��j�(�}��vZ	sק���܌c]���}��?�D�b,�M�OZ��
.&�;�����G�)����1Jnv3�4"��N8�A����K�eZ�xT�X�7���HT���(�-E���*���Ư��H6�A�˃��3@V,{ؓ]݇K��d�(�?ft�٨���
��z8�m�]��_M�_?=K�rѱW�����5{�� q�.�@��;�ı�l#���-��V�*���5�} K��\�����u���gu��s%Ʀ>"�[AI�=�b@��`����V�T��Y����_-���9��#?G��o�g!��J�){��þ�&ܶ�<�����N#^�����;� *ڕ�b��
�.�[�f��61L��-�%���M7@�S.[k�+�_>Be ���"�ڼ�9�l-���t��E�x���V�R�LN�m��e��� �HS��9�J�,������o���4ݾ����"�5I���@�o��Y�+���j̺�p�8�4!�_8t˷��]�7��.���/Ⱥ�����xF���w�C|�UM��`�0MB�N`i��@8�KB�Y$ N5�c}0���2@�i�e�Z����زz!J���(�I�s%tOUU(���y���`l�R��{N�E���d@��e�~*+?��8y� X�n4^���7(�5ov�>���j�:�ls{��2޺�0�`6��f�҆��I#Ʒ��73҃O�4p����6�ew�ײ}7xz�.�Q:��3M&�����<[�[��5yo��33���P��ӍF$��E>�����#����������@�K3:���S����u�����S����uU�hc	��#k���}I�"k���[�|��u�2@��e�
j�}�ƱE��Ih���0�X�/�f fb��+���E
)�H]�.@9|���L�f�yƈcV�x�.�� -�l�eGA�o+WV�����D4b��#��7C�h8�XԬj�\n/c�����w7�S8}wQ&K�#A���ኄW�6W�Bj!q��Z�fX{?x^aB�>,�s��@)��'�I���x�z�k�&MPs�?��h,�?�GҲ
f�1��n�K9�cC�v�'f�^nX*�4b��K����Z%ha����^�0e;��6���sb�Ϫ$����2E6	�A8��l���f ��<e�2����H�e������,Q3C�KEɱ(
~��J�8�2�.s�������x�u�p����f��=TFh�p�M�������Z6Z�o�~���2ḏ��n5Rx�m��\�����?sj��A�h:s,�<��]7��2󸃙��L���s��<��2��Vn��N6���N�{vkrd̠g�,ݘ��Mz:��D�=tGުS�Q���>c6�{�w�tw�DtMeً�3︫�&��$Wن�h.2��*����Ն����Y��l-8�����J]AgM��%��֩1.��:���ˆ'I-��餔 �o�������!����$cA� ���!�{�atG����u�Kǈ���m�e��c����`����Qw+ˢf���+g˄�[!"�V-������*Ӫ:��^"_���`��!D�dX+��T��D�F$�a��:>ui�sP�k��w�AJن#�s�/����b�O7����`Y+N��~��0����d*���+OM��X�����m]#�M���h�ö#��9�4��L�A𔭋�9߹(�����@R���*?�Z�w�W�Hk�хD�Z� �����"-�2³ќ��_��<�N�[�C�4;B�P�NF�]�:�V��iw���r���������%w�A��W֓Å���-�3��	���;0Op��v�����9����ʓ�^9v΍u\� _�咂��v�[Ǎ��ݓ�h?���R�!:|�Z&>�#���������3��FSy_oJ!�o����gy2{��P-l���Z��zC��썠�����I�c��:v�4W�z�~c��w1�?�o Y#�?�~'p=��ט�����Vk��K<(0���C��e~����2=`�+0m���[A�ET��ޠ�"�2�#I���(Gɸ�;�c��-d��IN����)#�Y�n�g����E"nN/G2\P�]�]4am��� _c`�~\b��%��ȔTjo2O�Xs��KJiB�v�X$fgk�CS�FR
���oi,�����R�N����B#�ip����--��n��	��FA��TVv��1W�� ACل�],���/Y��rn�aX�[�0��R?��i̸��fj�|���\1���1���5�fRS��F�hq��w�w��b�ŗ��i��
(#=�Z5S8�1!�:�m�L�z-�@�f�o��-�
G��|����нC�k��KM���Ib(�NL]�[4���;�3h*�� u
��/�� L.��U]V���<�AN"��uL���ʸH�m���	T�T�%�1q�>���\Da��A��i�e��٢?� ��+t�������=еx�3��!�i��%���RP���~OlR�� =8b$ra�D�-$��x�#�E�<]���ӹ�n��M��EN��3r>�/���ZưI���:UNf��vКmb��}S�f$RCу=	�+����M��M;NK\e��Ԇp��L�
����{W dnP�����k���т�S�+bJ������KOM�<f���W-���"�dN�X�)S
��m�U�"����g����p�p�k�N�˭��2!(�KNC�Q0Y�Ug�R�tj>���{���/���y�)����$�Њ����tn**�Xf�ǽ}���7�����m�<�e�u��T!����T�jFB��Y�QD?�m��D��8�1�Ҵ�g��ċ��+=?��3y��c�na �	T�Z�_!3��`�"F$}�ߕaM��2�A���}�z�PU{���!�-�r9��k���6;y���zB�'��İL��m�=���=Őb`�1u����!�Am��C.6�M9:B����Ԃ����KM�e�'�bO���U����E�I�Ӌ�ɥc�^*M�@��v(�\2�%��g���#)��	@��,5>��4ߢ{W6��PLX����G�vjm'�����'��&q���,°�(3#vn��(��У��n��]n�sUm�ц%Ug�;��U���ʔ�rBz�h�!�X�1 �Y=���lg�ߐe���Z=>}n��\e�Y�M4�q���ו����D�T��1i�Ni1Ϧ<�״2�������ѹں�z�c�B�0Ϗa��l�b���J��Z�΄0���C��Ah�+.���p3!�=�H�_{l�+�IWd{�pF�� �iR���-*��Oq�<*8W���bLXd�l�Q�3kb�.T��T�TSp��H�O?�x����H�j���7�A�u�u�����5�<�g:�}���6� /��@��]����bH�	g{*��Ňa� ��#�b��I-p��
E��Cpl[im��#�3�+~�c�5ӏ�%��|^+�<��+��W��Z�F�T�)��x� *��Q(��
�o<�H��"atD\���9���#�������`"�׃�N��|+~�����n�S��
d�d�Z\��KY�(��雤�g�Xp��mL�L�	^���}ݹr�F���"�`���������X_��%�K4B`R����"��K�6����&f�g\jDdyn�K�'��ت�����bA�/��6i�&$3��]
r(L��A�X��#X�\�`��6UB�<B��z'��|���F�z#�~0�34�A{�
���g	^���
P�e%z�1��l �k��Z���u	�c�BH���8����$$Iώ.M�P���[��'J,L�$��b�?��8���_fuPU��1�ܨ�% ���ut!�i����AX����+�^����b���6��U�W�a�<��W����Sox�0!�=���C2���������ӕ�Z��a_���+��u��FՒ��8�qT&�.��p2�5���0��Vמ�?L#'�A�$���v��Ą�y��+�3"�դ�a��pԦ ߥ@����g֔�;ԕ�wM�M�Nvl��*�v �Uy�#�L�gm��3����u�~｣v��K�~-�h��n�^��f�{~���� ^}��e�p���'"R��U�?�=�yG����[���q���2m�w�'.8p[O��[z�m�$�]�rB��vX��[�	Vɓ��u�Y!��'�s\U�\U�ź6H��Ss\[�-ʣԇ��/�L�r����WE�b�[�Ib���Y�hN3<%���X���E;㴥>�<������>%�N�!Kz�Kt6H}�#���ծ$n��:籺��/n�%���(�7��MgE���J�;T;��uEOUN��PL��DV���oΥ�� �"��}��K�#f���d���� �:��~����YI�od��lQ��>�F���v��������֓�n��'f���7�r��=����FX��35�p�h��3�