��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O��^x%���c_��$i��b�q-����O�-~\�MRTHx��Z�\0M?)���w�`+���AXS'��28c�
A���j!�ng1�-⦜������Y*�5��F���c�ۚ㏏��� <6`� �\�N~ɄC��+���>S}}�1���>Ac�@]en��}a�˨�ګu\��ʌ(jx��sR������/8Ew�t��s���<.oi����Ѿ��jZ��E�<��B�^ ���%8HY蝈�%���gK<�����_�	_)q!��w.ml*�DT&^~~EvT`�3|Im�+�z����'������G:���S��ye�K�X�M��hr֤�Ƚ�F�^ xC=^g�|�6@
8FH�~���o���p�\�u�o�euuM���Y��3w�=x,Y���q�Ia�7=��UBQ}�dܭ��r��Y���"�W�m9�z�<�ۯQF�9�4�*Klܫ���A�:��ѹ,���vD�G����U�楇���<4ݎVP��rs٢z{�����|D�ا�|Ƀ<�Z &R�Wqh������6�3Jh�5��F�{ �^�n[��bA+�V(-9��'ڞ� Jj[����Γ��o�S?���(v�LZg�)t�� ,8r:L���6�W�ܣDm��	�v3r����w7ɍZ歊�'@=�K�LZ��0��4b$�������.�7���Ā�2��CV���snJ�-75���Y�^c{$��'��?j��:�N	˵y+�a��At���$�rgc*I3����>�AxTᵏ������\�Q�G��T� ��H&�� N���*�,2��8YW~4��hH�Ja���N��ZԦ;	��Y��S�{�4�A��O�� ²�x}�bX5Z?��e�������2��
��)�
A#S-����A)�u��ά#�?.S�,�%�(r�&s��q����	V�P��YWp�a��:ꎱ)����(�?�-z�AMz5� ʘA3X m����������*�z�sN�Zi�%��i橆"���n���O8�G/60$���t���tS�9s�	���nM���M%G��R�_g8���-B���'0�_%Ģgh�UDa-a2fƀ��U��F`k�򦨉���w�u��Y��5����o�֙a�Cy��	xcE���խC��aD��>���fl�6$s��[	>��f�m��:����1��[~��m����к���J�E���A}���:G�8~2�6%ԨR_����(�/J#4MWm��F�b���׃�&���ì� '�����s;�i&�*pF!�\���X	V��ul`,�@�8�4D�ML�|T�x���#�@'-���{�ϬX6-1���/|��T���]�g���GB��GN���#%���dk k��&XN$|�I	���5Ȅ��-��0L͒�TIfc��J�A��$��cLN��\Z]��R�7�r5V����!��-��[8!+�9ݗX��V�'&1�լ�&�:0��v�2Kёwy�E9�����w-$��+����\)��j����h�k
��[&/���{ȣƸb4�p�F�����^<W����6h2k��IF������8�X�z�g�sRYtF���]pL�Ǥ����q�V950Σ������a��X��;�����BR�,�W���e�Jٻ��������8�{�Ru��i�"*�6����(Wn��m�	�/�����h(+�:��۟
_�1���ti���R��v�}%$mֽQ����;��gH���|��/�+��r���p��d@J��
��b�to���J�J�FT�5sy�f�*�W/Ŝ}є��*�#�1Wl�$��V{��]=�P�;T���5�~� �T��\Bq�֒�J;;��7U����Q��O�����㒬!��c�u��S��4�q�u��
3��S��:_�9۝�Eu���v��'MӅo��C�*F��fv1��JTe��
;��rg���p�pӂI*
������.�����D���b2Y�pv���Q�Ԯ��5s���A����z���]Ok�JDp[�^5�z�HY�&q�X����b�X�x/
��'G�FV{��&���Z�`i��p��ng�P�Q�J�<���y\~�L槰���ZF�V7;y�jH/	D��Υ�*��~����$�Kt�L���0S䳌?!>��G'4eS*�˧%(��Fj	Q������I����4����J����&�+����=�q�~j^1�%$͘@�j��G��$��|wl
���[_��rIǫC�"3��Kb�mp�kiX�'R~\Ն�{6(��$�!��1��'9���-'̳}~+A�/1ҟ42V�#�)A�T�0a�=��d2���3}��:(O��釠!Vh�5)~G��N����*s]S��9Ԑ����M���3����qxGDt�su�!�����L�_u8��)�j�V����!�����j�,ݕh9(f��,^:@��^�aH�w�.&Ϣ�.�Шd8�2�gi�*}^?��Q�@J�^O��&�h�	�׋���.�h�%S�[��a0b�1@h�d9�
a � �&�?7SF��)�ؠ�Ϥ��햣7N�D^3�T��"K#L�&e�Ss�"���7�Ꮼ��E>�   �5��w:�� g�!�Q��M���K�Z���X�� ����w��`a�-��� 8#� ]-��tN�RpWDf� mVN�_�.�Id�f�T�
9�PwD�*��zas�O��al� O��B .ףL�|�\fc}C�7�+:�]
��Rh5~h]d!i&�+�{�n �e����G��v%�ؼ�N{=�!AD�CQ�e�>�?Ȅz��O,���l�h)8X8���I��d�Κ���KY�y<��ᠴn��'���l)�7�B્�ӱ�nka���]�{����,���m�?��Z�> ����/Kb|y	JOuݾݣ�~��>m�@���Y���lp��k��t+���X~���"��dJI:kCJ�^J~��No��8>��B�,Y6hg�HO\�3tO�y���`��(���}�W�$I���Rc���Ȓ���j��k�)�k���u9Yg�},h�1��P ��E�#}��{� ��97�Wι�y��Mޅ`�5��kɝ���?����|?�H�6b�D^e�:�l��}�t?dMN%Wr(^R��j�;�o����-{�dL\�u��F�3�D�d]�EE{{U<��	`�!%@K�͑�s���tN�K]Y>aV#�Hx���U\�yS�%�AB�E琑Gg��&])A���5���W���Y���Wz��c�9=�$�y��ŋ��1y;g��k`�v!�8�Č��Ĥ+I$4_����Ԕ�C�+|�8��2`w=��Ȑo,k�(S 3�z~�G���9�Ɲ|�k	���q�&;��/�uͭ9^
��B�̃����y�������v�7�B[ ϐ�ɥ��y�������"�V+�%���_1�&���J2���Y������%�}:�"i��i!	Tcw���wI���mV���g�\>��r������+�����d��E����4rD�7�1�S�	����U�tŨ�Z����Ӗl/�q�Ƥ?�j�T�b#�}���c�rJ�M�t�w��#��m����&�g�� l���J�}:���-��������s��$�;�vd���|E\;p�g�+��x ���;T)��T��v�Z�>���tdq۝����v��١��n�h�k\AKX��) ����c��a��xh�΀��|U�r��l�=۷C�<��Diw�������J�m:~����2�9YM��j6�<8����ъ*��d �
��[8>Jp��Ξ�EZlG��;>�h�D�zPB�7%��`���f���.��I���[��m��� ���Q��F�4h��;3hk�ѓM�_�.��񷶦b~�N4@��ᗃ�J^���П?bF*n�E{
b���b�6do����c�M�"E���ٟ��.G�7lr�oV����$T���$�;˔�.piM��&fC\FlЖӭ����C��߯6�p�A��ѡū�8LV����;dۺ%Ì~����v��۹�ks� )�%�����:�a��ݕ��#�j�e��a��	;b�g'���=Y���b��!��#���c�yqw+,4�7��;C-���@�M���t�r�T�1�O�* ���&�k�/���7g������*!������I$�*y�� �ڗ���i��ԏ?x�ư�׍�Gە)J��t�V?�a�7�Lر:2EO3�_
"�ɸ�B�v���eB��R7��E��B8�_q�|##��T����H8�r���gKPL�Q�گ��m���@��m����u��0�����sفz�2���,;�~��9����%7��;6=�*�?���M��ߑʉ�
����vA_F,B1���C^Jv	���rԙ���$V�E#=���o����\[x#0��- 9�}ʝ���@���nCU$��{&�Dԃ�Wm�8����<�Y��>�PaW�
ȼtPY�)�5��9;�Q�[.KBeU�z�ziM���2S��ڸ� �Q��C��e�_ nz98b]���k��NG_h�Z�S�˃\�͌�c ���ʎ/
ٴVGľ��/�1�Бq�P({R�J?��8�މ���~M//����l�dm1������'�����"�����W%�����	9s�2�v�AT��?B<��d����t��5?�a� �m/{S��K��*¯i��¶Ғ��v�+O4��B���5H��C���])>R�G��9��JL��+ɂ;� �.����'��S)�hK��^d��y
V�k"Iu��=���%��V���6Sb%����^��b)�_�j���L�	U�,����h���c�z�Y�| 1U�_�̟�:��m����1��`SJA��1n�w�*���&xW�u�jΉh�x��@�	������Kv��N��[у�*B�>`�{v��]��{��|Z����䯚q�+ʔ$M��J�2��n��ٛ��}b-P}�IfF�0_5��4Z���G�]�6u�x���4��T~��|Z����Z&I��3��
0�����REM6�K�2]�Ur[���ă�'%$��|�>A�(���_Y����i�E]�=Uwmя풏\H?�����δ�*���j�ƺJ��A���M��1,xԝ6�����^��,$�<�F&N�Hfm����Oc ��e���I$dj�MX7z&��w�W�i��e�ZR4�N�z%�r�<
]�������)s�/���pk5u��!�.e��E����VŚ��b*H�#}�R���ލa�W������Y/� }����zr�P�M���l}����E��q.�m�ԅ����Nh�a��QrD��kk���|�O@S+86B>���hm�q�ޠ�����Ā�:<w�I=o81��H�O/zY�?Ѣ��ԷK�+p�ՊRU����"�䓃4b"��:S�j��e��p�P�tۂÐf/��~����b�i��s�~���t"��ǂO͛�s�@�~��������.Y��Z���5b`�\��y<�3�Qn&pz�p®H�t�%�G�����6�1L������Lfs�.���o�>s���l�_Q��f-[ S#J�c�j�ȯ7��Ͻk�����ݜ	Z�'A#؀	�wN@�;�t4�E����<�AMa�%�y�+���F�)��k�W+���O�#:eg|�ǎ�'��e���d���jؼO���!(���R8���7;�2��K��}�l8s;x?a�T�g�(ʫ=#���V��N=<:�L��IRo�Y���&�����1��nm�T���?��3BM��d�E-�gqR!�a���r+:�*��t?�<�9ẍ́�Rf�*��Û5z���M�v��_ ߹���*����Թ���w$~�}��c�����0X_� I��n�T�ib��j-��2|+��+�?�*��X	/�5�d^>�Vd�+��R�[re�����z)ޜ��P¡�$� �/�m\�����lE?���+���B���<S���+��c������O���$&��e�1�\)��	!��d��N@nZ�=ZfL� /!�	����l���k8D�İU��}M��e� g�#Y��I؊���y]Y�|�3\Yo��-�
�٭f:�W�.+�s�jT,�>�j���3�2�Ԓ��Q�wu����I�%�[~�x�}�)OR݆�gU�������P�Q����י@nolݫ�0�=WtRJ;�_v�4��8Z&�hRe�g?z�5`��iv�K����-��؊js������(�w�,(�CB���������7>�`�I�P��E�yY����NAf�0 `���1�����G�U�#
��P����Q����3\�9�֑��Z��9��`�gߤQ�m��ĺ1ik=�\��%5�x��տ%DL�Ӧh<��ʭ�ӯ�m��S*C:�H��p���m�!t����D�U��/��l���+�)��v�m�^�3���Aw<mw��.��"���ztw%�-�kQ�%w�69G�գ���e?5�T�a#�9��[��j�%T����sT�ŉ�3��~���;���P�ҭ��&��$t�=_��K�7���e�ū�#���+�Y+ns�Pdz��*p�~$޺��½��4z¾��|j=|$t����Az�K���^r��]e %���K���Bqtϔ�
:b.H������hȎ��`ǅƞ��4 [fk��r*o������b�%�1⡾�s�l	��rß��2�p*��!��a�Q�L*���Z���S|p�Wi�2�&�nF�J۩����&%�]̈��|-3�~=��D���GB�'�)u��5���i^	�� �+�3��_p�N}�J5Gl@G���AV'~kX#p"��]3�$/,+�4ؙN�_�_���'Y�W�\iF������$��`U�t��l|b��t ��,8�E��9��qA?�w�wʊ�A%f������=�
���=�ٟl���N�h]QOԵ�`v�&�(����݂���?���Q��*�i��0�F��q�h��)�\�,�P����<M5v�;��-��e>�Tb�'�.� /P���-�H+��(��o@��$�vB?b-�Y҄�N!e	j�ldh��EP��!R��˶:�)����5��X|��O+��r+O.�k����Z�)�dY\��(�%�$B*'e���X7y q\pJs��?ûw-�