��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~��_&kQs�\�K�v-���M��3�:��!Rm�-hH�rL�.Ĝ'�i��u$'c���T�Xڣq
�W���Oh�
*`}`�n����� m��؀����)r0V ���Y�D.W�������q���~_<�0F8�?fq��Y�����l��jYw	v��q���1�L�1�>�%��^V�aϙCۉ��Ю�e��c��t����ی����O��K:F�ޕt�%�R�`�ɒM�1Kӑ�n�̗�����MZ<�P	_��Q�3}�g����&<�>1KAɵ��/
��VH�.R��J*�F+I�Fx�|Ե�j��{��Q�e��j���
��ƚ�k��`{&�6�8�{�3�ϣl�'�Z5�7��b��B���W�
k��5�H�/�~������B��֙��I�w>�oP����W58c�xsXOQ�7�R��(�|	�M��IG5p��t2d�=���t��^��k�`��M"73�S<�W�(Z;�"K%����Z��� Og{�	X�'�k��w����?`@���-~����TRt::�)�[����
j������B�'�g~�B坬K/����t�e��Vﯼ����&���7;?�ܶ'� �����#z>ͼ᧥%�ڡ�\�ޔ��7�����I�Z�X���yY0n.�ȸ���lY��G�ur��G����A�m���pV?� 2��sh6�&� v��Ca�(����y�ԩ�՘Բ��	(���q4-C$� ?>����+lz!��t!N��?m�HS��Nia�ⷸ�l����	IHzU��|��2�&���4vн	U�嘓Q�3�["Ψm��_u@�rQL��M��� A�3��S �]�?�j.�|�wt�C~ˋ={���"�pn$S����g�����։��(�b���� ��߷�M����<��X��?d��78�Mߠ[�?*)E�#��VV�Omu����4A���6�:���GI�ω�!`�2�X��T��������`��ͪH���cX�\6G�)�ؑĶ(ɦ=����G?�о�����g�m|v�S�=O�T@�w� ?]	�~�N��.#��ۄ�Om�GG�-~rX�2�8���g �!�*?𞮷��5ϸ��`��&s�������By���Y C[�CgQ�tՉސ��]>���)��/��M8:���ft'6q�g#�R}��>�;�)7t�ca4����1�^�=�A�rP�� nC zîg�N�W쵡Bk(�|.��6��A��$!�ٻ�*���լEU�gM��K�Y�H-��FU&��4����U})�VHBg�ά�����r�^��E�d�*EӰ�p�S�'������I˚0�<q�9�d.���x����p��H����Hxt
��S�[>���#8`ˠ��@���r�����.�ADzS8.5��w�2�t��s��/\ȝJ#g�Vw�ڭhT��~B��.0K���3Q�p���mc�۔X�S6�ދ>g�Z�>&�"�fٽECf�"Ȁ: �чE�g����z�_W�t&�/{���z��5��;~�v*����J���{W���zP�j�hQ�P�#���
r!+��A�(2�J�&"�ɸ"�q�-���v�&T�\��8���8������2/o8���j�WA�1����CV�mv51��HJv6�¡R�o�����������2�@�&Q��O�lC�g�T��ٓŧqc��:��xQ{k��,�׏�(��<ʛG�h'j�WeU�-��*։���Z��k���a���E����X=�f��,�T�1AybӶ_��ٺ�SS���)�oϊ�Ȃ}9cf[]�yTׇ� p�7�!͛���	B������'@�r�y6Z�#��pVJ4N&e��&=��z	pb��:���B�1�D
P-�l���*Bg0��i��n�/�A���Pn�a`B. ��8�����G��JB�,�p
+�V���F]�EG(U��Źp�+u`�u"B!U�g:r��D
��,�N:�`�.��>[�o�97�nY~|4���}.r�3}@`~�ܕߏ��BJzi�!mQsI_T�Hp��-��X�QW���i|��}����Q��g (F��_ �fƺ��j���INm������%-��m���w5�6���E�Lc�4:"��,�X��B��QȬe��J	_ʦ��<���5Q
C��},�
L��690	J��K�<����?!����V��2K(���5��2yhc�|�,�b�MN?�MX_ey��>\=�3,��vC�<��L)��fPM�C9�sF~^�Okq�R�����en!@?�JÃ����bV�x\��k��<~�J�����ذ����y�WZ�@>�L�M�Pu5b��>�A�1�Y�I�Sd
B�*O6��jD �1P�6n����T8�X��??�������<ԟͪ�P�sV�`�G��Ai��Y�h����0�ĭ��`� ������3�М@���}�0� r,C�j������C�Đ��a��Z����vqM&�V�Ȱ	ld��GDL��@�?0�20�Cl@��f�l�jw"N�C�hn.,i�%#��còFc?�f�� ۀ�B┈�($�D�N���{�p�`HI_�x�I�Ҩz�)i(�����PZ�ӌ,�
�s������� (/��SQ�7���q`(�cp�W&�~��>��:+	�T���s@��~��z�A{y�X�p�H�'�,O��9��%����pR�җP��7�
�R5�Ǳu��0?��T&��!���H�x"]�l#�����9��Q��YId1�L�{��i��Ɖ@Gn�^_�I:q��UۜI�ΧX�ҬF�)§̳ ��W[���;Õ�8��IN@�}@y�i�P�{������|����+sb��"��7�=�G�:�� E��n'6��-��L�6���I�d�plD(|k��7_�l|`<�z��4 Ԝֈ'GZ!�ܰ �U�h��iHA�����镥' 
] 
��fl�a�#B٠����e$��$�4�a���MG[ SO.fS����c"��ֈ�%)�Ta�&�%�5)|�G��#��H�Pju's/�H�y��4y�����۔��� �X�j��zo!��^RC]����\7�H���vk#���v��C�#���ª#��e3Iu�����c��v�������0�^\eG_�j�	QlFdxa�t��m����;x7�1�0�w�fa	l"r2���nǉ��J�T��W�������+8����V�4�Na�8a	��r�SR�1����,i݈��?[�CF������)~�˹�x��6����ȡ����`��v�4�n��ǈ*�5�y��ӫ����Ё�҆�5�T�����r�ʫ����CL��`��������b���^�t�o�y�A�,��~쫖(��T�7�~��P�!*/��Ӯ����2�9���&P�́��j���ݺL��P�LZ��<y>�D���'���k:�ۇ�z��C�$-�~!O����L-i��.� �YFU�>-o�`\ �e��,����I���t"qbaؙ x�	�_�,�<U��X�HR�9N��d0|�Kq�|�_�0)�tLm7C9]����W�8����լ����r�J\hK�	j��Տ�gYJQ/���?Ӵ��Z�Zi&)V�V�,�H������m�K�J������<�:�_�,H�3���*#O�'ވy�!zwǓ��oCrP9	AL���=Ο�;_6H+����0k���4�\eNG��d,Tx�4�0�!�d)�|cX�Ca��L1|� ��RZ��q���j�~����ۻ��9i���|��1ϖ"~%�Wn�HN3@R1�5�W��� �=Y��ˮ�y�X��AشC��g��Et!��1�sjdiP���ȁ�q2.3:��5W���ӜF���@y�R�J��koV�Z�ޠΝ�l�M�/�+����uS�6��LRN�/��q��F�x�Q�Aeq��}�$[�)y1���.B��k�]��=��ֻ��5��	��rN�_����:}�.\�C�k�BN�����=�<� \���l�㽋���g5��N/U��G�fE�<� o!
��T �)mj��"j��IZ����=��
�+�ϛ+�p�?��5���I�RҊ�����Q�-x)}�Xv�Xj�iB_��?���\�)2�����※�t3
���gWπ��B�@4��j��(���~�d��<��9�QD�1����zNe,�9*�\Ь��-zƳG�	�~�K/[�Im4�� GU��O����m^��tp��S@�'a�=�>��sGx����^�xp�M�9wh�) �S��z�M���l;�!C��[�7~��H�)<��W�e,���iٕ�M��YȻ��R� ;��$ς�0#u(���IA~�)]c�lČWy��c��;=�k����WKz�ծw=^��J��]�{C��P�"�P&z��e�0�UzY���\'<�*��0t�\��tu���&�_x�Ű��5@���lFw���aq�v�wE_6X�p{��Ɓ��EOb
[ε�	�R��u��T�O��v�8f�ޢ,4ƪP�Y.��y6��V�-Ʌ���v��[��m<.��
�s��$b�.ݱ��i.��y�;m��ֱ��de�`�	x�a�����Mۄ@h���nŜ�1��"j3��Xhwf���ş���^���d�_����'�L7�����K)���+�-9����o��v�֧�EI�	�d��,��d�9re"Ѫ�����&�/�i $��'��/��_ �N�=#z֞Q�8cuK[1 3V�����`W'Ƴe����ќ�n�\7l�:�b�aK���LU�T�3�^�5u�u�����m�D~�<���3������K�i6�l�w�����d�VAI����[?��T��X~���\��� 
o��*��$W�r-<Ȳ̄gB�1Jj��Z�v�U#m�,4k`�,^c�Ӳ5)�|�����!<y��@J#�'U-�t��/��F�bL�Ϸ�\]#p��b����	��	NwH[�ud��/�_|��q��� �m[���Y���G���ރ��0F���X��X��v�����W2��
��� ,�TJ��eB�V���R�"�d5�Ю�ۿ��+����b�$D�3�����Q�&���Nk��l��]j�D]p���O	�N
A�_�P/��u�oV��#�#�	5vZS$��bby�ic/��	�;t1��*��2�P��i��G�o����տF��U����AH3�X�8"*{q�T���pJ<���%G��c�X!����U(	q��@DbY;���jia�2�>:Ln��>i���3�
3�o�[��]�2>��	E1�5V�.�C ۸O,��Q��#�I��L�N� ��c� ^���o�g+��IF��%
Qt��x�*S�k\��ڰ���&Uhnb�c}K(?��,��ȗ��*b�HF�7��i�H%`�RW K�܃�P(����i���i�G=�f{���#ߋ���>�y.�">z�H�S�,:])�G�Y?,Zg�6r�^�}Wu�/]�K�>y��ȇ�N�`��0G}�P�z�>�sZ�e�`��1�:\`��v�K��J�M��
�O4���~z,�G����_�2�6���RX|��ơzt(+�za�F9���M~8釢ɭ �^i��}T-T�dw`J�i�6���:�T<x��V�T�s<��l���P#H��2֐5�J۝��1�Ug�;�e߯nՊ�{�[�79N,���D�;��ߟ=�;���������R�N����OO9�Ŧ�&\��-�:TcŘ$�\�C��]j��V欹�?��ӽ�b� i�m��ed%��iSfp�aM�G,G��K9�[x����N�b7����w��в�V&
�{,t�V����S���y���[�G�4�$vc�2]ax����(��{���9���}6ih���/Iy&J�UۛC�i �Ս9�A�ؒ��Ď���Ê�>Y�\�\�E��KU��*�ء~H�U?
z�,��8$�I1V<K�m�'�>G<�K��2Y��K�U��<:�z�=��(�����@�v��l�m�0�Fn�T<�~��wϠ������^���tal�!$@k��^Љ��^����4wO�ǣJ��%�;�<�!�O�ڗ��S��o�~�ʛs�@r}�c�s�[	|���l+�v�"����=q��C�w��i���C�q8{�~����B������eE~0��4\�'
�͊�!ʹ�?U	��	OL��9l�+�K�F��]�-}���!%�1�s�%�uz�i���Z�k~��blUyx-?6�0L��7�=kP�3H�qI�gh�NL�P�L!a+�T`����!ǿڶ&%I����^�!�W���R�q��Ɲ�;��U�c�8��z�[RB{�9��R��d�7\����A�������j�w��>v" J]��2�n�B"T�]�!Q��U���ʛ�Zl>�s�W���x�	�y?�u�؃���C�gw���
{����G��Xi��]k�7{��h�x5a��ً!��&r�Ϲ�G)��BQ<&o ��!|h6���>zA[��,����iy �km����������V�J����z&�� �`�S6�r<�[���g^�y箸+�EJ�	��}ɱ,G-J�+��7ɡ��ح�Ⱦr&���_�m��c! ���2@�����r([b��([TX�� Y�yy�Ɵ.@�z�����]�W����Ѽ/90,�u�����~���<��iw;ɒ�60����y��v{-�~���6<�i˘�T�5�F�%}q6#�]�#�	��J�VF�ǃ����=[:e�;r82?��K5DHRm��q�	�3J�Ce:�o��%k>á� �-�S
{� $b��AU؜O��]uJ/�-`Dv���<؇�G\Ԧ�<C6��u�5b,���~^�|E�=��Nt
Ξ��D��Rt����I��D�m`��U�ֳ���q�`��Ӊ?��O":�w�ƥ$#���@4vWk5G)����j�z�\ ~�	;�Ty�}�nj���tz�D��z;���5|�_[IqT�CO����3���	���O-C(8�E�<"�l�$�H\�db�S̮ܯ�*�g�Pe>:�����]���3+\�'�a�:����*�b��/�j�;iVS`�/�v���t��C�M�ґ��Ҡ��P��w�#E_*��� "����k�]�6�"�����R��m���֌j�x?�����1��K��X�i�S;c ����4��XG9�6S��ÿY�cZ�`_�sH�J+��p����dA� x�f���4(șH�K��y�a�Х���h#�m�EI5�o:�,�ɍ�bN�2>��P
�i������=
}m�Q��m�?��8��0�l��E� �.O!�֥.
�՛*���������R!<�/�e7<4�1���ֽ��h.�Ͱ�Eo�ٔ�ڬG����ؘpݥ+A�c|�8o+�ͫ��9��w�u�>�iP>�B����Ѐ�6�Io��|4��X[bC_�Nn�x	ql�}:�^�rE}��
�>&��[-̓|��R�BH�1�I����C�?�̮g�7#���0F���k��$jMp��%�:�=�[q���&�;��� ;31A!��=�pMUc�;z�jk��@TFl�ΚD�D���T����EZ��G���X�}W����T�3�sJ��>�P�8#�H=�����9�*�H�i3J>9y| $<�vd����}j¼�y|��HR�XU�}��؃j��^�R���������������:XOr���!1ؾ���4��O`I���1?���7ӷwl�C!�_�w�J�"mr?V���i.T'BB�`�xY�tF����u����M�c)�Wm��=����`0�1|�P>ߪ�������Lc@Θ�!�D�������oYf�*�Y�Y$!�;Ź��#o`|���S9����\CO���ZhK�X�1�"Lg��;�mL�Z�m���
�Yl���4�s�궑L_J���@�H����wU�!2�́���@�v��i��"P��4�G�P��^��kE-�/8��Z�6�3v;T�γ��)Y�'�E�S�A���Iu���Yn��\N����+//�%������d�;Y[��33fr���a������V��R�����i��H��bӳ'�b� ��T������k�[�u�Ľ>�h�Hq�Y��/���w`[(ލ�?/�/FfJo�$E��$ܛ�nfh��������ژ�z�C�n�'"����Ж���]	�jQ��ŋ�+�l���3�^U9:�_����梒t��!"GD�EU����hC_�L}n\�FGq�G��Q7>��Ƴ�
�K�8��/�q�i�xUxM���7���p
�{e�9�	��5�qE�c�l��S������t��_t}W�cX�L7Ź�?���2�$!�(#��֫.�S�U�%�N�J�O�C�����崉�NE!��� ���G�|!%a�_�l�<n(�w�6��S�i�J@�5^9X,�	�c�J"�C���IN�E(v��ځCHȫ\����_�����	���%����د��Ƶ��l?d�4D�,�g��Q�F�2V�Ü.��_`�$�����cF~Ʒ���hŧj�,$�F��Ue¿���T%��'�}�G��鍸���.H��4>�m}�V�� �.�n��a�������5q>*[��^�:�qX���d)k2�(��/��m���� �Z��ѕK_���(�7��3�W���z(j�K�����G/�sP�	r�$��0)�E|������(�zcvkO�Tq.�9�G&���' ����Q
Ms@{Q�1�2%rk�����"G�x�u:��\W�8>��*ܮГ�R��m��O�]Ę8��CMџk��6�Ӄ�rA���pa{��r�ҙ��1�~7��W�"iM�@&��-��Xb�����2_�Y�4Ҕ2��R�eJ���vk��/;�0�咞�7#��	e�e�����!Ƃ����B�B������B�Iؚd��ԇ;6~�wh�����55�֧�墊���i>Z�jwׂ����9���hp�=!Oۅ�H������A(�Iy����IUi$@~��!K���m�p�@��|<���[�\�[�쐨�|kȜp2E��ev������e_( ��8O�݄ҩ�o�M1�fK��y��̙6�i��k����LP��ab��+���s6v��%� �)��q�L�u6��ef�ﲁ�J!@�5$h��ΈwK~��2��]wM�ݨ){����P�$�ʏP��oat"B��`1��9a �.Ҹ�ilw����������<a�%������6y��h�L
;�j�9�茠����ӳ2Mܶ��0u����-	�^�o��J�$�o�}�D�AIz<+�(\��6Ys*�f���4�������6m*�H�LGY_��F�k�5�3EӔu�m�t����{K���P�K�N�4���1�-M<;�jߡ1��`�p��ڶ"�����0�7]ᤝ!�҂���	G/Gt����$��Ɗ����n� �#�ү�҄N�ᱟ] $�{waS��ˍ#R`��͢�	)L�p~[ ���4cx�R�Z��1ax���xV��4��V��q�Z,�̸0�͒A�\��X�i��:<���b*Srܖ�~^[6]q��O�U���K�� 9�9��g:��v+~J��m�r��Xj�g��%=�\�䄩9v80�^T��:_]Kb�)=t�O'󦹺�x%M�A�R��l��!A�e�]�n<�+�S����]b@?w���:�e�����d�|��x�����޽��/껯��a�P|P1�D[$��HU�[.t��*j=�`p�v@>Wd�[��3��2�@���s�p7K:��A��x�f�������$�@��>E¬�#y�I�V#��������޼n�>v�åh���g�]��o�k�9�����V�_d,���e{|Q�*$�m�J����_#��G@d��I���L3x/��c�ʴ��b�Yg�Hn^��t���e���������� �Nq���\G��?��UAk�鯧C��qW�}���d"���"�CW�	1i[�2Q_�)c���#�uap�1x&
(o�\!�CF���pGT���6TԱi
�=�ಠt"��Th��mx�S0�"���v(�V��f�n-%h��d�3%��u0pkC�$�Я�O���[2� �aAG��~A^4U�u$������V�Xհ��T�����cc�����"5o�,�3�X97k�%���`�[j�����1��Y)�����"������3*ex�Y�
�dϱAI���G�;(����1�&�.k-^-�"���	PF�'��B�X���%�:��ԠX)�)�k�#'g^��ȣo�㠷»��u[l�ɨ?�����gx����Е
���K|���u�n|y����A����u����H����C��?$1��z�����-U7;��0bV�#j3Ksԓ�kq��ᬷ���?�����8����z�_-�o���#��ۙ�}87�&y�6��<_��7�>p:s�t���v��a�WL�t�C��9�w�H�E_h~}Ϟ��`�,��Zґ%�Qk'�����9�ÜbP�:��u+�^1<b����ʂ[�)�[�9!�dvӱ�Y:.�P:��}�%�4d@Z���&���>����
K����*��KHؒЦ���x�o����yޒ��L�k�I�ۣ��a�5� g�����W��U��V�1*����6���wu:�E����se�1�r>��GL��/���+�/���S���y�-�3����kJ���3n�B}`Vo�r��R�X䎯�9g��3�b�8RH���W�Y�v��}��c]ߵ-�gD�y����%A���^%��^�GGy��Fd����+9$q9�`�Q�,_:[Pr<X�.�|.a"���޻p^�w�����7����&��V�j՟�-��C�3'�6��AF���g��h���?wm`��"��\ӢQ�YK˰�χ�L7W��_���![ut�o��n!�}4w�ǇY΋`�+ur��U�gu>e�o�t�@��f�K'0^,'5��+Q7�K�͋�� �|�S�$��d�?l��{x|r�0P*%�H�P���T��Bt��6x���D��iakK�Ln1�����L�B�vu���h�z(Y�zE�I��$�}o��,��8��\��#M�!xDeBA�����s�@���9�U3Z*@p4�O���:�=uќ�� ��%v�����J��j�z��4e�\Rv���	7��|���R�l�xy�D5����["�:mk�ؗ�4�F���OO�hB������\�/o�OWr�K�朩T�P��j����h����&2���_�z����[��.�@�-��;o�`��P�sz��TD[��.7�����k��85m7�-Mp���r� �7ӻ�⅋�kӏ��� 8њ�u�� W?���/���ރ�߭.{KS>/@����F����eG�}����8��zE��A��!ϲ��ȿ��+�˛]��Q�!C�����X<Vg���𽰍�zh2t�e;8h;g~}�Bۊ���&Š�O`p��xvdk]�37>o�* �����Oi��M{�aQ��ݶ�fnҳ�X��=OCGk��5�R��"����,�@�du��/ ��U����Vj?�)��|�TȖ��2�E���:x�8��Q�꣥�eJ~.~����S�����vՑ���3u�R�V*���[��r�1��Žd��
���)z�Q�y*$Ḩ��A1�.�9:(��3�m��f���$L#u@��YYr�xۗ3Lc�����Z���)��DP�it>�ZQ�ç�-�0��jQ
K�n|��֫�jT2c0J
Т!IЪ90Xu%)l���qZG�ȿB��O��:O��g��i8M� }�BþpM���p�j� lD�~t�=&��]+��୭ ��V�s@y1����ęKB[�-��b)��鰦Dw��reђ-a�O���"KI�� ��D�v�q6�7�q���� g͹f�e(����4�� �zURQ3�ZM?�����nF}��G���~S�*�hy(ӋzR�;H�ك�W��F�p�dh5(c�9Ϸ��뾈�"�?�P�L���L�D��(��5�lP$v�r�k���9����U
�2Y�#�p�c�xek�l? R�'��� �fP��)oj_�q�AyOK�Y�?>�����
K[L�e�����]��+�+�Xq�Φ��$�ɢk7��M�i��h(:>���HE�	�	;�u�<=]!i��*���\����LX�ޘ�;@�^�0�SZ�I]ԧO,�A�,���&��5�����jB�;�7�9R^M����J`��<i��By��G�lP+E��4��$� ��kR��
~���Ҵy���|��ÔO�~����_e�sGb8�L�D����m�g�ԓ𛇶�i�-ڸ��
�0�^������~l ���^\�W]�E=�d��(4t���8ؖ(��I޸���h���������!;�0������_M9ȿ��@�$[�[;R�W^2�m��� 1�	(�,0�.%h�l�kt�1XRr��iw���x9�m��:���K��"�R��q�E��q(�˹�pu[�G�B�"������t�r�><�v~���!BO,	g��o>9?X�L�57ĸ���sF!&�t��{?$�O؎��Bl�F�O�nf0 4��qP���´��c�Z4̏2�I-;[v���1"È�͗��lL5K��n�}1\5*l��R��T���s���4�I��o��w�2���Gp��d�?�'�@���EF,�6�=��FpU��U}"��P���`ڡ��-ɐ<�����#I����6����&��;a}�3s��W3��T���kr�G �W��'�MZwY��?6)0P�	�n� 2/&���@L)Q؝�g� ٞ܂�N}\��m ���{�-�:�������K�Y�&� �C��I���#���P��;g��O�L���n�VJ����TsQXk@*D�Y���^��/}����r�aYi;��}6�Ueqjks�^����;��,����B��E�S�����%'��5�~���t��$�Y=W���Dj��KRT���C�gQ���W%@o�hߚ�B�K�-4G,��P'	'a�f�-��n�`#F��)D�&�|���ɥ)OuA�Gf[X�
Me@�:ӫմ��T�EQ)�jg����P��>�<WՓ�ŀ����D��@�
B���D�����+P�.�ѭ�{�_
_~,б�+��4�>�v��U�����l�ub[̱��J��+�s�hcm�ldMSJtK �Q9G�Oi�F_
�
T���1�J��;�P�w�����1�k�C|�$����~����0����kL�x���ʦ���%,��,U:iH?q7��$	��t�w�Q�q�1E:���j"�kZ1h7��F�~-
����0,
p�vԣ�2�� 7璃�I�T�X5yK��I����lo;����Ԧ�+��8��|MG��78�-L�RTQ����5}�b�x@Ф��|�[e��
��B�-����4�&[5�f�ư�qj��+�+��Y B�/yZ�_��. Bp�\6�.�.8��s�M�AA0)ZZ��I1��J;l���3�n2���!�v���V_?�Q�Z�GͮX�
q&�~�����7
�h���5�~w��`������Pb%�R�Rzz�Ui����y�L湳��l���{�/�-OD�_y�/j-��'�/�-)��2?ٳ9j>;?��;�z�x�q&v�(��E8a3m*�E�v��i-��W��P� ����H����Տo
�ܐx�b�����i���m�����<W����O���w=��6�o�����|A(��5��p��E�9�d�,0��}��x�݆��k�N��`(_ʲ�/Y�'}�Kd�J�D�o,�'�F�xm$,�)������'p�lHV�U!2ڧ��f�&:���Uߓ�)�5�A�E�����"�"q���,F��9:=�z�\��`�A�A�xNf%7c�QN]r�0���q��6����o3V��diym܈P�īӢ��a�������:%�`t���E��ů����ڽ��i �Cړ*I$��Uon6�K���a�Y#��;Wf�P����/s��#���	�}�4���S/{:WDWhTdךK���k��=�UC��r�Ԇg�RُHiV����"�22�ai��k�Q'�30mJ��G���A�]���AX9�L;������*!��U�	�'�kU�f/���v��&��tl4Z��e۽3���s�K�\�^x9d��SF�� KTb���_�WG(::��<ґj�(t��j��
$a�4'�A BƂ,U�F�o��e���������q����23ƫN�/ ���z/���c�ix���-u����Z/Ę�F�n�_�d[r���:�e)yD�8��=d�8V��[�/��_LkV�}�db���2���[<���,�u�"cD&��i�Zv20HZY��ܶ(��Gk��I�SK�u��oM�K׹W9~��呼��{��,ㅓL�W��7>f���p��eJٜ�
���[UE��� (�g~o��>"Z���ϑʷ�� M^%�m
�r�zW���_+���cE��<�+	�'Kh^�%}���Ñ�������t,�w퇂J�n��{�rTw��Y���}�<4$}�=��?�u�Nǽ�.��
!�ܴeWD&��qҬx�x&pꆜ�y�7���o�����mBm_N�뉈�����1Y]8�O��=�X@�Jj"��j@öo�^N��M�F�$q�Aތ+33�+���mBQ;�RA%&?4+��b�,�v0�$1���C��у�)b]��G��.��,ux�j3W�F����b}��q�9��~�)��.ݘ?���c!t;J/�wc����p�]5���P���)���1�y��b���{a���XHlh��h>XX�=C��}�Uw)0�Qץ횚-/�-�D��S1r�B��֚0lt�:�bd���5..��j�sHSV��Aa���܁V��6 ]<��CkJ�.����34(��y�
��hr���n�
${.}Њ�y�`��7[*F�����I�y�KU��`�������n��d&�=�S׀��ω�{�s7[w�E��ݴY�Y��u^^AhR4�l�����qgSN�#w�x�U�%t`X?�1�t@�/$G,���n{u�g����S\��霻��NȊx��ōU[�����j*�ҏ_��D7F���끎��0��ڼ�{��`T�� {�����y���ds�����D@����_��/V���6'�����cK�虞��ÿ�s���?b��-�W��v:�p�qv�u����n��i�n�֏�	H��Ql�d��5�l�ې��:H&�m�n/��U��Iy�̸p�@����_DSG�|��<
l,��PA,8�LȝK��L��d���UG��#���w�_ڲ�ϯ���C��Pqa±(��y����Z���tRU�q����C<��S�.R�+��'�1\��(�#lΆF6�	x�{T�B�'j��쾾sSG����	��x-Rt�F c���H�2d��@B����oY�e�n3{?pzM.%�v��=�A'�.�A�@�� ᲀ8n�s�JηCsHS�Ȯ� 7���G�DM-��a�,{��)�v�t|��H5iҽ�R7^�E0=��4&�������Lt��Y�N��g�M���'`��X����k2����� ���b=�)=�4�ӋBOdb�Ý͉�M|W�u�_pf���@� �"��ə9P�,�)_)O#68#I+�oq���?܁i8:��E��6m:���n�X��F=h���� ^���s���?�����'#�;��3ĝ���{�Il����j�&q=��� ��ή��<I�G׮��G��VRv8)���(ft����� 8��S-��h�8��O%�E�ڌBign�+iR����r���d�=�z��Xw'�ÁX�:g5�^���U�	�/�2mB�}���z�x�:m��1�T�h��j�Y'!](�FL\j*h3���| ��}Z���W�	<'�J�Z+&{���"�m�0<Te|�O���걚"�� ��`�.�:���r�aٌۤB�p�^aZa�� �C��7�9��9�i�#5R��3W��ó��B� ����

���ĵ����e<��湴��V�'�i8o���%���T�\�=�|�����k6��3��Ĳ�v���Ʀ(�3n�giLzdJ�S�0G�Y��S���a{�+R�Ը ��f��8�?�����%Ȳ������$�K�\������~����\�	XP�����{��{�ैq�!�z�8�H���7��G�:r�4t��yu/�R�Θ}M|�H�U�]�9�9�
c��*����l̑��N�E(�t�ju(%�@����c�D�G1���/=��0������]�H�1(�2����Dm4��a�hx�L�`>g�i�XxBbɂGШ��_���	�����C���en��g:ę���;�0�Xs`u���"���5�1V`��I��_��kb-��4�-#�JQ�Q<�/}E��N��h�ޱ���Ҟ��`֎JG��x'�r�*�oS��RtHc��U�m�xK({�7^S�-��:{�����i�x^~74����	^a1�iSd�¬�P"D�w�՚~�V�}T]�/-X�z���Dd	���Jx�2͏gs��Zu�=R�% vlw�E����=C]e0�����)ql	��9�}�Z�ˋO�]�D���./ă�j!Ɔ� BGKe<婣#��h}��Tb����N����927 x�.Iz�����u�I��d�C�y��]�	�mV�g�ɺ������@�[q�أ_Ӽ��Q�V��Z�6�w���řy' z��m��
كP�<���Ĩ�d �$[/6�NB?v�Nz�Ef�bx�(�*����V�ǩ$����G
�֠�+?m ��oSr��7,d�?�@��u�:��G ]e��m1��6q�"����/�e��ϰ�J0��Q4�>������4����ٖFY�r��p��~���ڙ�]t�L�
r�Ֆ��S�T!<�o�;�=s<��"6k���|��?z�X��[�^ȧB�6��-���<��ҟ׌2���`K	rM�3ס\
'�MQ^��z�(�nQ�S9�~��L4G��	�o�_�4�)&��&�u�2����Z'O.�#����
"�J����O�/��?�ٍp
\M�Eꂍ2Ii-0]���q���
-���$+-�p\�=����"�ҭ�+0@b��$j��ʿ%'%|5��%k��9!�k?6<XO��+���(�G龨iU4O�Aژ�q����v�;)���(a.���5i�O���$	Lu��.}	�M��������p�5G�{��E�y�?��5�O�`�kTmŬ4i�D�F�A�Y��qo�:#�淟�ܚlG�)#׊q��rɤ�Q{c�3�ѵ�ǌ��l�2�����985s�	;�~B�������w�l����|�6,�e[�E!&�]L��kM�'j>���*r���U�1*��C�Xe�m�K�+J��l��J��$�<|vxJ�F�
� ��,U}#��#I2�����!݁�ز7H�j'N\�!�e���-M=wϷ�|5��A)��{���&�˝;';�ǁGu��5T7í�5�(���������X�0���K��pˠ�xq+�Z�n�e��"�PJ��u�ѩ
̥�����J�}� �$J@�P��a��|dZ�y�C�fĘRf�g3�KU��u�P�_F�Xt�.f�5�I��3�����s���NA�_'��J$��u��t��C6~hB�2��cӃv�>H�;�A�u3qH�U"D��m[n���Ӏu��ƌ���Q��D<q���������r4�	(k���#qE	��d��b��:����}Ja�.(���b�[:�k��l��[˪)`�^a�g�⁇R�����)�m��B��r+��
�
O��]՛�7hZ�/��Q���S�DTN;�Q�M|N�ĕ�G�� ��Mc�d���"���l�/^�
�">����(s�{_����6���ģ��cT��(+��ך/������ɝ�
��w�}���D�n$�g��mi5���9�z7�hٱ� 4 w� ����Y+p!��Հ{^J�x/`�y)�N����ΰ9b�>���=86��i�NuTƞ/]ZD�_a�o�<x�;�C�p���>ԫ��K�N1��9U���T�A����k5���R��'Y�;�Q�n��*l�p_D9X<$�R��B3�� �4>;��Fz��&'�h�
K���,җ�]�*�@F���=��Z��K���Y#�@�X��-�H��1)y�b��0�%�!�1U!���(�T�h
N���Z'��2�J_��bpr�k���0^�`ՔН�U���Ǹ,�1c�]ݑ�
i#/ C��<z! HK��&��\�-k.31�{�R{.�/t�`�f�EgjaI"�����g7�m~��D�Si��:�y~'���rP�8��+I:�m�~1��fJ�ك�擷�5*�K������P�H�+�r,������NC�#%��PA��?�������'�+��/�A�
���g�)��Y�g��W>�5�EX@��E�٫B8���a��3�uz�l�x{�lq�a��dn(�m��#i����s��Y9䪗�������&�hM�"6kS�����*���,�v��`z/��5B ���d���Ua6�(�e�Ѣ`����4Y��hY��4���ПJ25�&�m�hUPDڝZ�/H�&w|�u��=���i9�Nt�.��na���jQ}��z��A�VyZ� %T�SoF�C��v=H},�T#�x��ƹy9֬������ ���P~j�9�,}r�,���7�FK&��b^�n0waй�Qn�