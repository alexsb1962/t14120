��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����@H
v��T��bg�KT0=��?�G��X������8�,&Y���a�g,{~��ۤ��C�'�%��`K��6ӽi��z�V��&	0?��vq;�����YO�;�x��������Q~�yۮ����؏O��x�����Ŕ�[�b�{<��B���̽�ue����<2��p�R����[7�w+�#/ ęK��(��{$)"y�}o�P|\J`V5.|e�v�v���
�=���\8��>#Ps�9'QQA?����#�:NP�{(溴�����=�;;�%�qT9e�℄^��S��g����1�Ȑ��;�$2t��gnr$K�@B�ަ'����zTJq�K�7{r��PBˠY�T������v�Y�4��w�yV���Uy]�D\�b���l�y�j�68�׼��1z�;�*�x��'T4�ݑl@�Wh�#I�C�,��N)ZA�C��
"��;j��eR?����������;�;]~�{�'���j��O�߼�?? ǫ~�v�i���T֎Z�}#9���i.�0�8��ٟ��\�@{�v����,i�xi�h��R��;9s3��;dH�	�j��_��M�$S�u���>AL��{U��^���i�z�I�wZ����"�L���|aR��S,��J���A6�i9�@�	�;�W��j�Ȕ	���?BXfU)�C}-�)(��־W�y
��H�n^���t�k��%��u�}!&��%��c��5L#t}^���y��.�~�G�W��� ��ʴ��z������H�I),1˓m�dC9B�Y��D�d�ܐckZ�����ow����A���7d$LexT=����G�3L^��(�^2�;r�g]�`ر�ȬS�.#�4=�Α����u<J��7�)�ot|��(#�g���h*1�_z��P�����K�
�ݞ�
/sx�*�b��O[�/�6	8F��)!�Κ�ħDH��-ԫ�;qS�������4Q��k�Ԧ7L�P��Jq)���d�G]`o*S��j�<�)�l�E����� �a��9�
���͍	��K�6�_Hkʇ���W��A�F���7�,�ٌ�����+�dI��W&��3Xz;Յ�$�1��m9I�������2����|��&q�#�`�0�sD�r�-~\�B�0�֐CY2���N]��ԏ�o�ѻ�dHQ3��w%(���К���XI\���3����9 ��H��qF��������h��%�~ke��N�D����=,� �G��c|-�_�	>�/����<����(�'Aiq��!̂�%�rhJ�-�	�3E�0�rB�DZڈ�/��sqa�r� hӇrfͭ�����A�|��G%j*�F˛!U��hk^�Aa¸��MM�6Y*��ԏ�D=�Y��6S�Ru�=y9�Lo��R�o�"ٞx�Y��A�2�@����y%��f�Xo.2���S������r�Xz�v7���?w7�rށ��7I�k	ĕ^� ~�`�Qr��x��e|����I����4x�m��G���*ꑾ�/ i�,���kV9'd��f��Ѩ��n��ΰ��V�F�*A9��ˮ����[�K����_��)@���i��l��+�s�1�>K�n�ܬ��$F4+� '�֭v�k�{=�/1Tj������|�z�*�(cICe^-ĎI��o���4P�E�r��r�Q�͝�1@�@^���R�+��p�r�Vs*�W�f��PQ~��OBmQ��|������E*]�lPޭ)�,vQFD��@�,�*J(}Y ݉8�z�*'; DTwAOz:nxn�"�W4������4���:�~�ڌ��d�PA� �WDkd�憈�[�{����u��>�msWbO��Uǉ�b���iĶ��نTC�ih�oU��\z ��ch[��L��]2%�9Hꔅ��uUr�ϭ+���	��������@�Z`��rs=�=�~fU��I(|���+�V��������L5�%r~{��P��.���`4�D�!���a��{֑
Y����+���mQ�����[6Řx0� �qe|���}0 ��Jb	���{S$8sgq�
���g�*W7�#"�|�z�Apΐ�� ��t��bH�/���v�O�2F��ߓ���8�_i�8�}�s}E53���PK{�=#"��6!�MI�7�Hq ���Ʈ�IB���6Mp>��i��@=���y��n����j\/&��>-}5���N��c(�;��{��v/E)��6j�D{W4
?���5 0׈\����Ҩ# ��\bBP��s�O�H�J��:�G�$��3�??tQ���=_7�|����#J��A0��݊u���~8�/cU��Z�Ba@�^2�Y�S,nN�T�%Z��|j`L�|A�܃kM󅨪��*���й�3�Y@2Ze!�L��s��r�
}��~ـ�G���T���Fn�Q�WZ7�^̹}C`�E\䂌�)����a����h�[gK3>��J�mnl�q�3ǽ��Zi����l�܅-��:w�l�ke�۠YEi#rٔMhY-ω�J >0��M��(�峾���~w�]m�n��g�I�Ġ��̝��Ã��׍��w8�o~�o����Nһ~~ү� �2�#�D:ղ���v�wz���v�e"���ĵ*J��Pe���X� �S%:\cUOϊ#U��o(�&�Eq5���t�fM����ƣe�o;��U����N�zgkDF�I�Ǹޏ5z�/.�%M�1r�\�@H/ҝ4ri�y�=5>ӒH�Y3�bl���嘯)�xxc���Ptxoۧ����A�Y��N���orG�IkT����2-g.'��H��ˮ��/m��Û�Y�U;6X��BT�9���4������/��M%(�+���`|8� o.Ɯ��&���zŷ��Ê��Dp)�����0+}WzP>}za�uc�:��5��>oEnj��+@ЬoĆP�C1W:Uu�3�#�]���S�C�Sf3��r��m�%�&�AP������P�*KȷCZ����#
���ޡ���C�Ǟ�+��b���zE�K�~�E�>���M��̣:Dw+�������XPd7�u}�=|�s�d42��2o;��^�:ކ��L@�^46�FR��U�1k��e\�r�D��%.Qn0������%Q�j����!��<ȳ���-{z�x���{�
��|��:�Q}�󿊡+�jk�Ͽ�tq����N�jq ���u�V5D�R���ޥ$;��4�.���ҴhY�������^75\R�`����ewf�U��{���hx���0���1�rNeUVV�7��@x�j~ʌ�T�|�w] �K)�^A�h�=�Ƨ�t��cL��H#v�迼p"��ɦ�	�������M�b^�2���V�}+	�8���cy�� ��u1����`����e�"�ǫ0x�MJ���}ObH����q�E/�r�������j#�Y��y+�>��ÇN�\��32C~�@s���J�*�T�J*�m��=cݏ� YB�y��	h���slX�|���� ��4�`���2�b���f��I�(�2�d,�$x,��y~�p6�rFߧ�� 	�"xF��x&��`��L�bVz5�l���cnR���`�]@Z�b�>G����"��~���iw�X(�<��t%9ݐ���L�(�E�����#��4׆�+��n!M+�fja�ݠ�ф��ߜ�.�V�r���n���b���QQ�2��-1	�:���*�+R`���lݥ'6��fl;��@	�zx��4B��'���.��6,��������W���^���UI]�ާ!����G-�k�2U{W�P*�ba�^5��}`Q-6�wt���w+ @�j��ac���+ Z�u1W �����e˙N���b�iV�]����ѷ�w�^������o���~�X�H&1��	9QZ&����H���	��;mg��ʊ-��x�ߣk�t��N�A �Q�\�p�h$�]9t��NZ��"hvJ@Ц�����u�4���j�6Ms�����?mF�[��6��R�t�&���n[KnG���[����"�G�q��&z���A�2�$�&��(���8丰�K�%��)y�pp�t4�V�;+�5_m���k����i�3���-D*��;��)lͷ恟�Ck!~#R�4�V ��6gkJ�B� ���Ѫ:9��^����/�P!,��&'��Vo��IS���'X�B�Z�&n��ˮ6!��4�^\G�J�����G{l=��=q�J��<2G�d�d�^y�E��B�Q���d.�h�4c5y�"�?��5�h&�����o��~}?�f"4��L�C���ԉJ�Z���$/�Iy�����i�[����b~�J�p���?-����ԙ��M������	�WG�V��{���e�y�K�'?�Y��	��F*d���`T}�J��]}J�t���?x�I�u���?n�%���;�~����]л	�	u�'z��^����j|)���������6(J�]�}ӯ�qȸW�P0Ԓ%Vɾ����{�k�i�7ι�m�g2��+��^h�$"����d�|TX��:�QgjW���v��ŗ�Qac��۬(1�]f ǀ��/�{5'@JCq)%Qsg�w-.�;(�_�Ƒ;�H��z����\�D U���g*�M��sT�(��I͙�F�aM��w��k.}a���% �$����1�^iiu�����x$��6�Snd-�y@��iB�m�G~N�<iT��č,7�J�0��9�D����TN�����#*�s���;�oݠ�}�Bq����)�ݧ���\�?����߯6#�1E��!�_eTH�,�Bx��Æ�z�"������gBz�n̮�������IƯ ����1`k#��ݓK����(��T�F��'��qRmd�ŽAw��s���b����͉w	h����KO��Z�4X����䴌>��-�Xn�R)_3�-`P�Y9���������k����_T�-�g{HϞ�I�p���d�f]��+-��q���6�D�4u�Ə�qo��A�����y&v��۫�o�]���edL��i��̚*[Y48�H&J;��`�t��:�j�J=0���2y��Rſ��v!���!N���3�<�ڜ�[��S0G~_Ё�Z2{���@n�C�x����Q8��e���-���BG<�=Ψ!��C��hB�����N�rs�H妫3{qY�ǩ�H�Ro5߬�G��,�����@�J��I#�u/i��~.�u�Pش��v��oa��1�' =�M0q�d�>�h�z�?d	� ��S:.��lZ��<�0��G�)��}�;�u�/]b��ӆL4ߖ`/:��xc(��nX=!�֞� �#��q���epԢ�M�J�Gc�?0�2�M^(�w-.SFΡx4/�"�fƢ�[iS�BpZ�R���}�"�,%�c����ݛ���K[&�<�8��䀍�1
��R�j��H%;�׺�'��D�j����V����4�����iM�z��?� �Iom��{�;�톺tb��ê0\3�ԴX&�}���F���'�~�yO������J�D�a��iqj7�{��359�U�p�G�_y����e�~�U��'2���3Bga���w��DB���#��e���� 5.�Q�pF�Pہ��^�$2�=�a���$x=�K�Js;�Kꇅ�F�%�m��>&�m���H��P�fK$�5x���^\P+�oQ�(N ��B�˅�U� �s@����:ID��j*�'!	��2��$�T��_h����k� �R.����Rz�M����)�p�J�Բm?\�Xu�c���Xr6�X8�C-e�@]'����l����=�܏9?8��Nڑ(��[�A2Mv��N�ȣ`T��o<�\崘�%R���?u�q���P��ڜ��ܟ����u���5�y����1Դ3�>)���l��r��A���@-�Kj��)�u֫���3T%��|7�U�a��`���5��'8wq=�/��"�s{�(���zZu,��;�4a��;.k1@4k(����!�����%i�Wh-�{��'���z	8j$��I�$-���D//�`��g@��+��'ȅ4�5?J���Z8I}g�KL��-�U�eS���f�eY<�v1�Te,x�������-Z���\�=�'.v��
&�l%���U��6+���E��i��SP�eY"�k9;�O^}������k*|#���|̩���4�r"f+�}����6X"�x���"2Ղ2�����(h�KS���k�4ZR^RM�R��:��+`�}�p2L�
�Jה��7N��b Ws�:��P�5���q��Uttj6���G��>��6t��Q�����DF/�+e0@_����z�e�ϳj��;j�+4��s�׼t�����B^7}�.s���>��G��K̥AE=�f��F��e��
eSӫ�[���>�t�Y[��`H6u��.�Eh?�>�gHp��Ț틗��>�'�yݸi@6X���+]�֊}�S3)�A�Ȃ��I�v/�b) ���=���,��5�	Pg� )L�Lɵ�=��X�R����H+@v,�?;�ԃ?�\�T�.���C�������'ڇф���U_I�Z�9R��6�m�L�;�w�nMӛբ���:���c�P�[�^l\~�5��� `���W�{I9ݛ��yS�#�fbҏ�؋`��N��%A�4���Q�B�x%� @@�(�/2'�Ak�f�9��%K]5��W�CĔ�,�aCn����a��	�p�u
�ЯRVm�S2a��b9���f�ԭE���1�c���t5�+���#�Β"��Rh��YL^n�ɶ	�l�ٱ5N��3���X4������a�ɸ� u"�Z��$[��dv0� T