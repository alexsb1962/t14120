��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\���=��sl�^��V����Y�D�?oqbN�H��/�u��;�oqS�\9����)j�Y��RZ�x�h����*Z�Ű4�_�E^�&�<fN���:j���p�"n3����V�P�T[A��'��*i��~LYWϚ1��ͅ��j�B1����/�~D�]o�$z�$i_�p-��Q��MMf�Vr�TC-������S�;��G$� �Y���I������jX�F"HmH�B�q�.� B�F�ģ��;S��dcq�VN&$����;J��m��
�Ϸ����*�O�y,�����I�%f�O# �}�m����?�p<�)� ����7�7nd^��H���fVN�;c��/���k| \�_V6@�b�$���gg�ʱ(��F0������&�9&dk)�,-��?Uc�={?��ݵ�%G�o�Y��3{��4��d�m�Uοp#�/YJ���4"�?F�\?|-�G ��X
�`4�#qH��Pu!���NW1�#���1�*�$�	�,�[���P�so.|2;�ө�{�i�4fk���;�L��=�~���,ح ��T��!��=
:Y\��^����L�M�|�9���ť2��Z�[��T���8��F@���e�r����I m�2�2���`7�e�$�v���/�,J�V��Ӗ#�6�A*O,Љ���ψ���N��x�w�"B�~Σ�6�H����� #EҦ�����j^'���0���Y��j��u�����*>n�/�ਐ�ÜJZ�����z(���ot����ȥ�\Ƚ"��u��VC��zJ�@&"�b��)(]���Bu6�<඀�A�����\HX�tE��K-�������F=��e��kn��^�A��H��4��/��ݷ;M�8�L5wFUv���4��
ް2����6C9�V�F�r}�7�pݥ�?1�>N�^E���{����u��F`K��z��mWq
�����~�Ġuޔ!���~ֆ�6ӿ(W��� :�}�X1�5(���Xi�X���1����3�������vMN%�1t� &w�Z����4���f���K%����Kc{����A���n=�?m�3[�L�����_�ה��e5q�6p�#%�KgTk�f�?0x׵���*)�[vR#-=��>���E�?��=�3
��S�;���
A吼��V�ʖ��ۖ	��͞\�o�	ɵ�RАWظ4t!�'�I�����jd����Hד��
B��d��멥�����6䗆�j抝zL/;/�?�d�����˿�)���3��'!��r��ֲ�Mc�v ��X�&�˽a��҂��j��h��G�_���xG�r]--| >���c��v6�����L��J�S�t�,�C4x�n
��8G�C�����D���g����O���6}���4���ҋ3��?(�J�O��"��
呷 ���E� ;U(.�=�!���|m��Y+,� �y!3z����H;s� {�]y�gk�F���d��72)����Z� �>���3��:.4.�qo9l�%��B�; ʃ���+�\bu.���t ������Ĳ)	e��$BGX$G#�J�w��[^�)�.IoC�!��<��g�}W�@��y����NW{���OC��7�GOx�Ѓ}��1�9�"x�r��[YŇ�0��0���OU�]�QV�?
�$���T�ZI�.�"��9&��?y,�K�6/�ǘ����.��'.��d�N���W�A��9�����#��t�J�P��~K|0��L�"R����Ó1�"N��7i��*t�o���!�PS�b�TO���-%���y���H�޼�q�T!���E#b�Ui6&��������#A	 ��[�t餚=unL�R�.O�~'��^TX>���v���W���?k~��%E�5��Rƶ�C��7���ۆ����@Wp>�R��G�F���=��Iw+����4f��e�#�s�!}� �49�w���}&��Og��Y�8]������7�z8�I^�~3�� �h�e�sW��������(�U�-��Nw���E(�.Mq�'��y�I�a,�m�L�7���Kވ�Yi�J̒�nx���}Gt���Z�zz��m�n�$���4�]���O.�W��>O`�w-���D��QNt��V�	u�'�&��T��� �n)�p�p�=�h�R-�������}�1[|J�S[�8��hk,#'"��&����D�"u/*q�����c �!WA�'�SU���G��o8��\^=�~j��̜�3Juk��Vci*)X�#�2�H���@/VV���[ŕY1����\I+��F�%�ua4�vo3�\x��+�P����Ӑ�b�7��-�_���S�'z��қb�rh��{g�W�i��a��U��M�<��T��6�*�բ���[v��R8[r�[�*�U�n��n����ӭ����,+x6�e��f��z���E��h�	)�2ʶ�~l/�,���^zh�_�KE!}��γH���0,5��"�,40�f���fN�$�zI쑪�da�7�k�+�Z"_?�$�F�|�w7�(��MxP<1�ji�B�43c#������M	����� %Lg�FL*�(Ǖ�+���lH���l)���ǧ���ZQg�p�h����7A��x���x9#a*ûoCf`��wo?�!��]�\׮��b��#��/[��f�� ǹ�n̤�FR bA��Xl���{����bR�l�@��/����BA:��vkl�&u'����g��|��"w��y���e��%�@O��p�����H�+)RƋ� �H3��2������}P��b���sʒZ�`�;%f�I ���.�׿
	�p(����w����cc���. ]��K�^����S/�r��6z��/�/7t��j�k���(�������*9'��L��j��K>��"O�=�D�Q��s��l��䏜�S	�bN@���;�(��/G�K��
ܚIMXl�e��*�߅��ÁƏ���l�J�m�ɏe�\��<��0匓��6C�;^�p�z0�x(��.�p�%"]�q�;^W���>�s�
��~_�7�&���%L$��G��'��%�ȘP˕��#R��%,�Ǉ0��KC� �8� O��J�V�(W��_L��7�	���/Q�S�lF<�\�4�$�3����#筧\�e3�\GkA�E̫�Qgn+�6`)LCʀ��$�Q�J0��*oUl"89���:�ǺS�y~O�4Fm�4:�xp!1͸.��Z͒�r���Y ?��_��^8��K�r#UH�1J���tR!�
z
�[R$6ӄs�'M�ֱ2s��DC̯j�ő#[!3�I�V �=���)�
g0 ��A�*�r[z⚚h,z0'/\$]�pz�!@bٌ��hm%I������U���钊S4���h�#A]�^�+���ߟ����Z�y�i#(k��r�����@W"�Q�A��;�a���/�)<�%I���BvTC%�����Q1_B���R�~�\��}�g��<�r:� ���}`G�
�X�ҭ	c������j?��Q���_a���+m�J�5n�&�.9^��>������'�[�U�}�.M�!�ʖG��b�{p�s�<�3�P��d�|6�j��왜:]�3�&[BbܠI�U��'Zfe��W%�P����G4z��e����r��(l��/?�d^^�%MĬ /Ɏ�K��@-Uv~ק��W�EX��]A$|�i7��M������6&�fQT����$��͞����Yq�ٝ�P��c/16(�:L�`S�s�D�4�Ҟ&��.�cW��֏���!i�X��Kc<7����}���`C\�>�c��*�n�k�cz��I��)��'���%�Ճ��#xv[)�&E�ZBc�36е��>�\�Ǖ'~l�e˰N8׏��K"��.���X:�{_j>�n�ݑ�3�<Ȩ��H�'Y33�?�?;����Ԗ�?É���I�q
��:l.���.�s"��
"�ة)%��[k������[�E��(C�/�]!5�y�5� c�?S�ԙ�,���G������3���^nxj*JSP�{`�0�q�@)'}ӭ	!��t�27v�����1���#rJo��)BDp��B�UZcK[�ɢ�@}i�x��]�	M]�����!�����H��<��Y���I��Q�S#�t@�m�m"C����Uw���2�ʦ��$�D��X.�\���n��%����@[���G2�aE~1Ɩ�nX�2Py�7,��I>��X>
�`�/A��޲|_�7h.6����l������j]=��H�{&&f�a����i
'�w���*u�B[7���o�b#p�� �x��d��C[l�҈��Y]�}6�����ݭ��|����З��z6�L2�*,�p��C���@��UBT����`#u�'��	hK�ȵ�������#F�~c��|��?����	%�LxXċCUգh��d��
�.��"5c�ԫB�fy�=�9Zu��P��5a6�3�YD9��8����j.�U��}4���b�&��J�^7�$Ȥ��hP�o��Lq�OÌPP��!2"���/�t�Kk;G-=`�?*�\6a���G�<T��D1��=gޕ}��@*�Ar6��.Ո�y)����p�ZP_D~K*2�1�'#{P��AG�n	�;������C(!��p����;!��q{_|�0�N�
4ܙ_jO�###��h[XN������^1Q�2�����ܨKۓ��S�R oJ�ұ�oK0�E9v��g�*KG����ܙ���2���É�f90AQ����$wǒ�v��� �\\�@J�3�?:v ��D>h�}i�rf�����?ʥ�{*��Ř87��I�£.�95n���$"K�ݥK�&Xrv��5�f� �C8�Dt��
뽿�b�bG4L��2<2���Ry,�Fo-��9��,~�I��;�/m�0�c�@g���K��2����_ӨۄC�/��,ȕ�y;ہsf�8x�}[�4���K\���+� ��?�Ȟm�XU�F�]d�|[�w4����z�-��M�W���!I���vf9�iI]�H�W�d�� ���u+�!���3�9�-��Ap��wmo�hr�2��I4��u,�0�p��>Կ�/Wo��7[���� X�I�lf����Cf�r=�X4籦~��n��bşW�
<7��EB�C���ߌ`'x<@ڱ�[M `�-�A����\]4~��u� ���=�����gE�1�[SBq�}�q
0�cV܃���71�T�CZl8�ݫ�?Z��SL�>��l+6�9������!w��1:ck�HP�����Ծg��/~��{(��</H�3 XJ5������	ʲ<w`Jr���e�'�C��kb���"�W��R���#[$�r�(�nYY�\ٙ�P�6�"-��Ua=��
����3k�❾��� ;��8EI1j�,l��=��3�9B��g8�c��B�B�ؒ��	�S�Z�r��/���j�Xx������A�����ɩD�5=C��^4I�L
���}"�F��o��?�Ț2D��Ҧ�r3�kK'Md���W�>�0ɜ���bo�����V���6��CwD;pO�U�����.rYJz����D4�����"=-���w0"=i?���[!���~��o�V,87�I8Ng�5 ����,���D,�j�-�W��_2Y]��`\g'�P�4}��=���T ���s�D��b��RĢ�����2W�E�_�E�8!gXJj�j|��`��� W�@gu��y�r���l؀{U�6[��� �l��!X�?��?P��vZ�����Ô��L�ƙ{���l��M��2���UX3�)�zȰ$y�� �n_K������.*���#�zȔौhަ�J�n��W0o&�H��V���H��P���h��+��LL��k�;�m+B]z}���?7�v&G~X,��]	��a{�e^Ӻf{�,ՙ�˸�vW��W�B�����h	&�u�P�<xiC5?���b�c��.>`�g�{��#�5�*�L'y�rfN�d[���T@�:'�^X#����zIY4�P�\�n;���iil���>m4^`
h&��d���B���9�bD.�j�ٲ)7���s�%�Q��d#��d�'�Sԇ�ݚ<��qD�Bm��t�(��qc6Ƥ�H=++fq���ԠVvP(,�&���s�}0A��)0� �,����JB(�R�^�t����Vߗ�8�,D�x�m�����&�dU�&̝nߊ1����7�z�g�;/�rI�_pQ�cX�-�z;BA��5��S{sF}@I$e����� H�����c�ʦ���#c2��,p^X��Z��#�+ԧŉ?�kN>rd����R+{r6���O�U[���?�N�'�� -�{A�XL-ln�%�2�K~j9��}�π�%�2�ʫI"���[�\g��A�1��iOj%_�j.�];���l�o?�Ɛ*f"CM��t����_uw@%B����f�A��z빐G��*� I,���-:6�Ş��L��v "y�!�� ��!��<���l�"A�.#�a�h���j�r�^�~�{�"[�#]ZZsD ����ow�O"J�WҼ�_.�pc�*>/�aؖ点�׹3��TNe�í���.x�pa��w��x
�Yz��V���Լ�n�~pI%�N�5H���?���?���T���s���3V�����0��Q(��E�	���O�k���׍eYd��t��`̾)Qb���ߒ���O���
���rHO>-�6�+'�>�g�Rxr
˗+|*I���&��_�E�9�z�UC
�& �b*/18B�)��1����>�A+:@����h�w����9��� ����\��Sb���l����d𽜩,��0FK����(C�QU~e�l��~e��[����mf�O2�d�%Jy{˻�z�C(�K��m��VH��Τ���!�QN��֦a{��ʒ�߯�\eF8��Ĺ�D�wY���L^���� �6h�1�6��(C��r�NJ/6B�W�)�T� ��,�P1t�����FB�mk�fo2���`%g��rV�>׉ૉw(U�����s/�4���=`_ܼ�
�$}?�i[��Ļ�G�ͱ�crup*N�61�+�Lj� � �/�q���Ar��P��(Ao[Bc��ip](�]gλK����S�8���N��[]p��G�TΑ�U�H� ��O=:RG4;5:�M[��Q]�k*9��^���ތ܀����F%�&,ؙ@���E
�����
��������-k0<"�^y��6�sHG�}��L�"�u͎��o��_��+����Ɏ5�*ލ!Èh���괿�M�gNk���f�ϝ;��烐�~R+��m����Z�ܗ�}���ss�~ci ���=}6�x�鉗m����$7 �qF�.NO��R�w��w��
�ˆ�X��e���E�Z�	"�_{R�( ƚq�;eB
�e++�!0=��U3�s�si�yr�0�n�f��'� r�(w@��y@'��c�(((�������~D#✲_�M�Mþ��(�|S��=sA�p�$}�	f*�Y�'1�/`���
5��-�z$����#����� W�>�R�u#��w��0 �bѭ�ƹ<�<a�ɽ|8�m��:��%����BZ�)5�t�`e��qD8�s���4<BȱgPHk^9����z��pѱ	v� ���ү�L\����}�(W2��Vw+���޾�Y�d��1��#y[_�a��455����ް���|��@��Q���g\�/c����ɺN�y* \�\7Nc��(A�\�{��K���#+u���P ����d3�n��I������l�+�$������N-J�\��}�S���+j8���E:$��ٲy�10[�?�f'�]��][��,�����{��'I[�o��ԕ�k(����Qeр{7���x�q���C�pm�찫Fɭ8S��;9ݬp��=>)�?�Y#p6@P&��R��a	��,/���X$V����'[��<�s�o�@�L�̳W���Ȩ�w����,E��i�%�I�(�H��wݚ(҇��U�i�z��{���	���*(���~S��y��̯V��ïX�U�`���p��a�6
<i?㒎�P�>�.x�LK��,�������}��֥�8'_NXy���C��@�Xn�w�#W��)�Kt!���OD���O�gl��HWR^h�5�%V(���u�5��i������S��\����ݞ����?@��I����$����]`�bK|=�T�!@�MB����v��=4�iM�n;�ˆ:�^�ns��0�ɢ�,̀��5iݴ7`�']�r��Z.��"�U��K"��v���r�M6��q���e3�����e{3�mk�!V�C���^�F�<~ԉ٬\ GIsh �B�xARi�=l/)U�9VGP۷���N+�̸}ތ�Y7�7�K��M��`G7�?2�a���}��$81��02�ߐac���4�Pn�jyɷ*S�/�w=�).k���p�_�F	@��_x��S=>x�x�)#�/���\�ɗ���%k.Hd�(���̲�+��rL�d-�9r�=����m�v>��_>�k��,E�tM���T�GΑh=�_K��>��0���uႝ~�:��y'y�I�w�e\�B=�}��w��%Z��hm?W/�>"�2��y�B�t3���<��.��P�d���q��{
�sf��-�Λ�ǙS$N�g%P�$�(<lq�%���}�d~K���p<,�aK����҉7_|đ�9&��E�Z�pX|=��<�#��Zp����6�q����%VN��v�;�a;�/k��̐��|�{�]�e��nԿ�:^�X{�)�}�a¥��㗆���+4�z	�[����;i.cN| �CP�G�������)����P���LZ�����Vw��v��'5�*?���@r�S젚�������>ި�F�L�K
��5OE�Z���Y1�,���Op.R ��`i���c�ؽ��L.K�?���3��E�=c=�`?�Ӓ^c��0A�2�.��9<L62�#���ـ����D��]ѿt���2�0��QS�IM���Sc�0�O�����+~4��jZ�.zIlg�s�u�𽟄�0ΏY6ϕwb�Qܝ������M)H�w�QrI����um�n� ����b;��kH�Ft;[ʘ��������I�,�&;h��dU��q�B$�wbn��Ѣr��h����s#�套,�Mx^6���\��8�)�����0���a�ՌR�S��iLS*����bh̀��x��7%p�?��2=$S��B�Yu�JgWԈkg|8֌548�%�N����ؖ�%g6�!�	�,5�m.�[c�iA�MJ��oF���0�X఩��.vv��Q����]��Tw�%��ܬߗnl[��d��g6��剬+���eQ�uv�t.̩��j�_-D�3�(��L����Cx'�;LպE�j�݉C�j��V 0��7�}	١e���<S$d,��y�m4�s�2�\a�{��0ڬX\�p�$t��-J�Nn�M�aC�NU)�0{E�&Hl�g����"ݣ�#pr��t�*w�]�jqSչr_����}L�J2��֔$���.���ZR��r�vfz%����u��E���<�V@7��v���q>�~l�P$:�!y�2��#q$?�d��kus�]�J�A��V��9�lnv�F�e-����7s�b��j���e���x�7��q$ 9K��1�#[5�b嗍O�R�bF��2���˲b[L��4�ے�A���7d/X�*��)��S�w�a+2<�^���r	��`�βh,�"�XL��o���lp��*�c�[��
�6=���
m��؆QF0��t�
�.ß��L4i��[�nx�����0�������r<����ʥ���bj�	`���֌mGU�x��#d,�+��W��p�e�[��#���!�]Q�!js��[o�5�,�Ǹn�l���Z�r�$/��l�o�c�Q۩F���\�L2$�xH���G�%��բ�)x��;����q�͗j����8JP�g�Z����Ab�􆢌�%\��7�T���lp����Ĺǆ�$�-�o��g�lf����QP�Dd�!�h��H�qt��jj�g;M�6��ʤ�"d���FtV{�a������D.����uu��:ۊ�V�[*c�P������)w�.x(-
��E��$��|�_A>��d �LL�(v�uX��'v���G<��1�VG�Z�4R�ncj�r����p��i��&x����w�Ŋ�K����&m,qE��Z���y�Z�%a:�<R�}	�
�(�����\�@�V�ȍ'H��Ƈ�UǈZƕ� �HV6g��ʞ̲�
P|�l���M�*�F�Ŋ����p_VU�N��4`�W��`����#�	��+Gk���iF��2�!J�7��C�h�wY�/�Z��� gO���Ju�y�z���$��m�۰P�\Y�*����8
"���8N��IE��A4?flIn��{ZѸ]�4��R�ń�[�v\�A�RG+�ԭb���� Gw��,���yS4B)߼>4E��0�#wȧ$�fYl����f���A�2��1�v7�ب$��_'3�*�Kk�W�-"Bd��ʱ '�P�}p%�|A_ P+�P�bӜ�9������EǸy��kdw#��XU�Ws"�-*���!�l/��j����Z��v��3�I�����rz�|�S��z�F�M���L���<��6yUX�wr��!�*a�L1yp�a ���n������S%�5fMh��sQ�_��M�H`������] �=L���A�"�d��+�1�Sa��Q����5Hd��d>Ss�Y�7e-u�?_����n�f�,{Q��&����o^�d�խ�^�aT���&�G�����Y~�/W��7�j��~��L����u�b�č��s�F�"��E�4c����Y��*�.�u훅r��Ѳ 9c�" Ew���:�ʻnYX��`�Y���+ن��u��#G���KP9��������ʟ�L/�w{�:o�-!���! e[�����D�R��Ap����޺�e�/�%���3R�'E��!+K��{�~�L��5R�/�{j�cV�Ehҥhp-�ے(O2��E!M�~!d����[���L0i�#�n���$
+�ܺԀxfX���l�Ĩ��z)!���~	r[J3��?k�Ë&�st$��kv���9Kn�t���;�T���8�憠��8|T�Д��-͏A4|��*�q-V}�(�d<�P��c:B�	���MlL`H�=�ٶ
0��:���Lo^�c�<S��([�_�T�E1��i�C,�� �˂?�VFba���9��_ ��{���E�Y���X3���I]K���n�3]�r��°��=��J!�kПoˑ�[>��S�,��pȀ7SDur�77��)�w�sw�Ehy�p���0��Q�#��34ٌ�Zũ3��}�%��AmDB�	 u��&۱?�W�tx�[���)=˽�o"=�P�f�Y�0AQ�~0�qD�剗�X�����"?��Tt���2�p|��!�ݷ\��Mgi�vt���u����t�u~g��iL���j��z �͔(9�6N��#�Z�h\@�໐(��.\S���~ �1�c����߉�T�dpf���*ı8�c�c��~�����W�Y��$2*<��3k�3�mBq=�vXK
��l��{��J�������Hg������D�o�h|q�rϤ½3�����H�u��zP�e���OeQ�O��8�_�>�iY�ʜ�����������^%�a�h�)��L���ݷ���Ň:�!��g^ �CH�/x�ICS�@� ��DB��:w1�b�Dٞ��-(z�d���N����BE3b��'Oр��߹Nܥ������f����t���[ۄnO\�nK�� {����+B��W�|�]���mo�k���z.P���^)Nu��(,���p�+��EBY\ORfq���yq�F�%~^Jy�����
�5�<�bh��2�օ���`D%�����ӆ�a3@iK(4�%�z�7�S�:��"@�l|��Rz�ݦ��I'3U)�oK�C�^�E?Gr�,����|�Nի���oC�����oԪb�(|�Y�/Fjً�vȾu����N��M@�ܮ@��������T���J����)��s�Haq΂�*�k�c|�f�bYǞ�f�gj5?�s��N�ń�6�0+ +���U:� �/:��ލ�����	��y�=U0��1 �^܀ �!ß@ߐoбZNʲ	�!y"�'.����ˆ9���NcY@�*�E������ U�R$w��Ac���uY-{rbM�-�d��*��ֹ��;��6�{�S+w��Yzo�(�)
�
�k������et6'�����jÃ;�� *�.�B賕/�U��-@_���ھ���n�׻��M6��j�U���A��3�cw�
O.���I�k�ba�k��ZSC#9�B{���;*~�׀ן���	\2a���o��,��9��Y]!ڗ����k%���F��A�s|��/�9�,{����D���^�z����3s�w���ؖ��
�Ҿ{����UTD�*�/$ ���vs+ΗI��[�W��q����h�D*�ɐ/h�#�I�M�?<�v Ζ�v@�����9�(DjϾ51$�8GZW(ivf��Uth�}O����k3��������f�p�_�{���Ih�$��H|���Ѯe�� -���R�.�?:i�����!���5��o��,�y\�Z\;��臨-p���!��˅e�)XL����}��Y��5�lڑ��5��$/�΂_<Oә���+��,[!ˠ��H�J���<��h`@}s���3��(r��n)�r����y���F�-���`G��O/�>0T������N�'�S�4�P`l��[%,d�KH�7�e�%I�æ�OȽ2�NfVlޑ>?Px�A������\�z��5ͺ��f_����V8�h(r 43���0,S~/1�T�&#.�(a���������Y4>y��iIEAf�� W����B�W�9�P�쭿��)�(
|A����IOE�8��BJP����ȃ���=��U\���s=i��1Q��L>����j�d{��Q������&�����Q�h�ʧ� �3Qf�rN��-Z�*��&7Ƅ�m%��,"Ld�n��L��`I��8�|+��WԜ�����O�}CK��g�d�ƞ��`rP�yt��߮�v�A����̕p躞��m���]E�z�� E���,��iբ���gҦ����oS_�MQ9�fy�@����A��$YUTF��Nzh�1�`�ae�VlR��Z���1Ik��`��[�^Tk5`(3�(^7��K�?�rR@P�肿n]a�.�n��V纒�d���Cb ] ��`�A-ʨ�;l �K�A$ܕ'��Av��Z�;���m[�/�}�ʊ����,����ƨ�ń��$���q�vGr7�l���W��ȟ({����Lwx�ڜ�_b�3� I|0�!E�u��a�K����RIL���"o�4&�lkq��	j& �Q���*�
z`!r�%�Z��L=�n���9�L:���џZ�$E$6*=�colP���E^[^HոF1V�(_bJ���H�ZXƷ��`1ޤ9�����u��l�;*���))��U��!X�"�G���,9eM����
�Q��7�muj����֕�'&��x�Od�-��9BF.V��|j��)!���kN��NY��@$�~q�;����`�I�A�X�'~!|��=��O���[
�Z����+|�YO{iB�U�:[�cN���uQ��	�y]�aIozƈ�S�
��:a@�ߛ�k����>SĹ��T��G��9V^�h��jd��N��"4�.��U��!�t����/�')��pR�3��]���G�G��`)dA�?a!}sG�|��a��i�m�n��/ַ�e9ȁ���.�e��E�����7��}�8P��7���/z�t� �U,�H~l����5P%�:������ϸ��T�A�|Ӣ0<�Շ�E��`���������ӫz胱��>���̱B�G�I���f�7���-;R�[��
�")`1ͶT�r��)�́M����vH5�?��\��f��վ��/Ӂ��¼'�x�ΐ��N�x�Zs?_�Ó��L��x��?ڨ	�N��B�^������v~W�H�Kq�م)�䮭�x^G�Ԁ{aD�H\��l,IJ<�i}Ň�<'��)su!��%��k����%�����+��*���5Od|�J��Eh1)����,:���C~�z���������J������Rr�DI8�Y��-��IQ� *Q���W��zv�����Ҏ�w���uC6�Nk�1�Tq��7����gbh��tl���I���x[��1���3���\b����t��,E��wUx��M�U���f�Ba~�G�в1냢/<&o5��s�#�<� �cڥ��
�Y1�k(4��X\J��ͪ�B�/ �`
�B�d��ȭhy���A��u/ݜ�'Q�=�����.ؘ�$����I�qd)�TV�
f��餔<�������=<��hL��H�����	��cB�A��\��-���V�7;�6��N�F�N��fg����D���ҡ�d<cL�`?�{��.5��`&�E-JF��@�s�CQM�N��$�w�X1�s�&�}Ť�خ�Қ�>۟���}m�2�o_�6��O��-w7�BJ̯fA����F��(�S�%9�k��y�$D��߀m*9\wRǊ�z/�-�o@��P�+풕9���P�cG������V=}JήOv�>�G 'y&��B�Cԛ�m@�kg�U��6� 5o!+����+��	վڎE�{���M�Q�·z�xue r�i�b@4k����D�&���V�\`j�`R����5��C3���M�{N��Q��D��A	D�(���<�קȶM�g��"��P᤼��Ny@���T���CΚHI;?��t�I�s�h<z��'4$\��kƩ���*�|Gy���o�W��,��uػco�Y&������(�#ג->0��
�������[K4���ca�`�3o?�*b�T�'?$�G�M���u���k`�'�6Ј�;9j��bKA�RR(�h�l%���#IZlaO�Z$��Հ���	���7���4�8���-����(u�����+���D�x9txM�S>U�m^d_�a������:����V�г݂�d����ތ�#'�E
�>���d��F|����T�xa~5� ��7�nx��u�����y��V��%�%�0�Y��G�C��"����YL�q�č�i����������5"��Y��A5w���|)���Mq�c�g��F�\MJc#�9=3I>�bBIZ	��5o��5��XE�t�=��H�ݩ�H�*Y�dތ$�	&�M�g��W#�cQ#,KI��|Y_�'�6C���b�]U�i�ǯL�g�I/&��h��+�����:XM�B�=�IC�!f	�|	�h�V�$y�Q)?��)��C�a4g�gm˙�g����"�a����LSV�6�#�� ��D����B�8��2h�1&N#�,��X���~�Cb#��G�t�'{AYWW����[�%~����n] �+q����˅�m�H�J�`7��s]M��ߠt�n1���=C���U� �%q����}�A��hH�j����as�Dz���55L�Dˆ�~k���y6J��Ǟ�` �S+����/�σӭ|����SO��+G<,;�m��K�VU&��L��RO����7j��L��ӣ�^/��N�Cn݄��.9��L' �o@�nϞ/�<C�V
h�_c��m�sҒ}�^���3 ���f��뤇\[�,a3�����%j��9V^	ҁ��!��$��2�8	��M�Hw[���
%���;$�JB�_���`b[B睈9��$]�^�s\��<�UP&h���zT���
����9�|�IU>ܒ�02�(p��\7*|7�Z�ݗm�p@��$f��0�\���e�Ȉ)�̜x���?��l*�|;���3٫%'nY���h%ae�>�%��mח����|f����k��Z!31�:��Ƙ���R0��1_��g/rue��h-�祄�$Q�q;A)�
X*�c=嚓����
Z���!�S��� �ʈ�G���q��P�	uE�w�w.Qe+���{D����2�s��$JQ�����.�o z#�~P:H�V}O������^{�V�aT��3xu纆�)���mEJ�o/���d���S�9u�C�����IL���FJ�T�3W��d�̗v|�M?���ް�d<%�o_�o[���Ax@�K��3��[۫��,���t(��{T��QY�1�Z�s�z�g?�S�J-p7��0��Y�hO\�&c��E�:@��*@�2�@h"#�Sư�T�z+��1OU�1R9�k�[\���)�r��C�[��k�L:@��J]tzw�8g8�6�5�@��Q*k�t�$�m���o׭RK�N`�iXe�Q��Ov-�9�o#<5����NS���F�i�cw�+8����LN������G��c	��f2r)N�vI093X�,�s"Q4�n�Kg�M���p&���v���|��J�E��K>$��ɈY�p-i ��3
ʖpD���; tΚK*�{]VOd���܈�=�/�����*m��y?O<�+�e�ꍶ�|��c;N�~������z ���ZG���x`P}֝^T}W-�R�m��1�lHz$;��ɺ?�^���NNf�P쾄w�H��1C��ڟ�{L�&�\a$�pxH@Y��v�VV=���r]m�ؙ���E8�F0��@���hrJ�.f������'�Tf�e��1;]b�م0
2�;s�L���1