��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����Dg��Q�ȫ�K�� ɉ���ޘt�:|�M
ؗXh��Xb�Le��7�-��Q�1���>Z_�5�1���?��hyҔ�o��N�	#�X�x����&h���puV\EԼ��Tg���4�2Xd�?���ck�\��S��nQrY��5����N����)i��{^�`Cn���့nA��ߩ*��~�[/���jV�3��N�WE����7a�R|��t�p�*��͆ԕ=~h.#|�>XZ�|?)\v��Y��*I\H9�<W!�D�ʢ�'�V��F��4J��2�a���ӫ�ā�q��wYx�E�h兑����\�wX6*E(�����i�T��4�o_ �s]��Gx���+�����1{���p�f�Hm������r�kkI?���㈹i�98��$���w<���^���������p��o�@#
Q��~J��<8<�^�m�Щ/���x�ʓBBu�#�e�m#��A����-�8�0HŌ�f:���r�W�#
�!c��Y���LC����E���k�B���I�2Fp�pHjeg ��AQ��X���g���6꺿�~���-�w��W8].��|t#Z�G=I�kv��ڱ��q�w��d��G�6�)[��_ߞ�!2�(�H���ܹ�#:\�C1X-�ا	b�������ui��lT�)w�H��:�G!��� w#�xCH���}���.�E����Wi�{/��b_Փ���8
p;�d�;G�p��_�\� )���a�Y��|�5�!?��'$�´�|V9|Ptm�Fj�B|lEKC.6��QDG���IohE���\�����TFk-I);�Y���LV�?O'4�G`
�3Jه�N�,���at��J�*�|N:P�|�I q9�=�yW����KӪ�/�,�E�|B��e�I,��y#6�9W���N%P��� ����k���(+@��Ҹ!��4RS�^�-
ˈ�
��_���?8�A��\�mv ��$$R���h���H���`H]u��3�P���;�Wk���|,ګ�G�^]{���B�*؟6����x^dD/A�|Cd�g?rՆ����"��?����Q6�,��C�m��j��A(.�E|�Z�Y@��bg��JNhD��e�O,���9 ���.G`HX�e�
����s�ɒ��(?�����(�t�9�	�+����.k�G�'�8oϳ��΂�S����w���qI��`�6�#�@����)��{�)�Pu���yX�	V��x"�Y�d�C}���h������0�sq������S�)B�G]GX6���1���<�ld���W��|q�<$ڎ32�S����x�fDE}����+���P��}t#���cT��+�_��FIw3u�7�G�}��_�����v:C2x������`������h7 �ӚW�2�[�F�8����_p�Z��������B���������.�};Jc�42��Uc�n$�%����Ŀ;ӻ]��󑜚	����Q�X�	XlO#�W:�
�����	n���aY|���`�W�5+�xG7b�&��݃]����6�-�L�6a��7:�P�o)nBn��)�(jlW��D�3e�?�٠����
�,LP��R:$Y�T�|�-�L��l�p��b��F��7S��Fh�����q{��o"�S�w~Y�	"V��o���[6^�_s?�oN��ި��R�e$m��p�R�n!5���Qr�.:�Qt���۠6���X��4�Z�D��<����szi`n���~OϘ�T;W����u�4��_5!g�^�{^���5?��B5�?b��bgG�'���3�JO@�E��*.H6��o���ߵʭMy��,Jk� Dm��A?�H��9�Sۇ(�`���)���-���U���E0����a+G-��ھ���ϳ�a�" )u@���}4|�tUb��Z����
ճ�(V��Nw�Ț��(��Q��m������66@j�(�X�L2K�3��[��]b��B����qbi�-�a�p�ɦ�`ś�X���2}'���e��F�h3(yｯU75G����t���V��x*����ġ^M���a��7��.�]��J�,��� �)�;ʾ�Τq;SE�� f[&�Gr�X�s����"Ag���F�s���U=������h;	~����Cb��N�و�(>i^�A��B~O�K��h�5RM�ΰ{̊:{�R�'!k0�ޣ�U֞p}�\&h�8�]�B�dXyZ�3��9M0m?*�]���RR8roJ��%�2нد�m>Ұ� ����<&	g�N�0���m��W�g/�7�_�f��Mi�9^$�:l:z��w�)�W�q��]����H��<t^"n��|͎y����un׎¬Xs~��[<�Z^�i7�gj>B��zx�Ns�D�K�&���%Nz��:|U�>�v�v��;�[?�_M�_���*��k���{r����u�diVKM��R+��/n��tL��L���Q�I����9(����p�CSW �5L��M��1�Es��r��h�rv9�εc��
 �3�$ŹP��iĊ@����$E?��s`3�`���$]��J��t�1d�v%��R�G#h󳘟9�7$IT�S���%��w!z�A�F��s"�̎��!:/l�����^X��u8��5�ej��+{��0t���;�B�N�s�_H�y����4�K��v�e'��k��5�.���M��؋�fnH�\U��yڮmkQ]����@��"�Cñ"b� Tل�T{���1����杈�M��Y%q�{�?^�xaP�<�YpFu�Bu���rXHJ�����!��y��RTYA��Zz�u� &Mf�cΟ�ǈ}��=)�y!�>���H$)�.2��d㯽�Z
�L��Ѣ )c����*$ǘ^�f3��J����'	Kq�����٩������w1Q���"�|�Ep0�5�7p�,
����8�ѻ//Fd���Dtĸq���Tk`z�����XWm�i"��V\�ˁ�U�~����9F��)�;JgZ�Il���0�3I�g�#�Ə�jO>�r����9}�f����"K�7~�0+Z(���р: �q�ɡO�e��!^^<Kh�_X���op\ek:Ąſ��JӂiIyp'	�8��e;E����A����%Ѹ���I�ߌg����gФs����m������~T�x��}�X�l�y����OԬ����$mD����k�|zjH*��٭��r��K6���Ε�	'�i�*�j�p<��Z~L�������{w�fw\3V42,8�@B0�p��MT��;f��"o���m�Ǖ��FXm���Jp?vi&U���W�gj�������E�Ե�ܑ�Rf��e��2�%nH��Xl��E��}6�=�#�����D���JK���H���~&��v��.�GBu�^u>tL��@B�"?�$�q��س2>6�
��^��ސ.�MU��MR�4v�\_Q!��@p�˷�.h!^�>�Yj�g�Un+��3��,^����UjrLLx�K��?�͑\��gP�gl�?��L��1
���Q/��o [�,��y4�Zl��/�iD-�e��� }�	�4>�+W��jw^����gj<9;������ԩg��߄C�I���[�h8 ��bEXVY$�k��k�5��J�a/z�P�s0��Ol����&������>���v�)L��Zj�q��p�B��QM����nI����F�*��xi\AY��������� �1�x1b5p�<#3��g\b���������q�_��飄lBx���7�1R�SVضS/����j"���<}���%��U/��J�� W��V��ܳޜ,��$(�{�1��w־���pk.����]���I�����ޕyU!�t��qƪU>��(���2~��] r7��n�qUU���K�CxuVcp�%�'�hT�?ѹ^Ǚ�E<3��]ʅ�5$XÃ1Lc��V.��]�^>�[�I��/M��W|�-�o�|د��8s�����MOXM�'�/�r^��� C(��zzL�����&��!����\vƲ%���zvZHH9���	�A"x��U������ <�i�[%N�ߌ�?��<��,N}|���Nұ�?��3�o��g~Pʆu�E��l|L���\u��M��w�8 �Co?�2e~ֹ�3ض�V?�*E�z��&-˰)μ~$e��N��b[XLEZ:�e�ڌ5�7�j��G����&ҙ�������ǧ��_���� ���+�)r*�N�e���`��RS���w{��ryc�=qU'��Ί�����1q�ژS�8�[�ر�g�Y������Y�QQ�˙ض�ٯ7��z����x���m��D�e��\CˣJ�/	�}��7�H;�b�2����n�W�}�l�̱'̩0T-�H�ش�*��a�z���H�6����4��\2���Upsh��>�.�c���c�U&�=�D��!���$M��/�:�!�����
��9Jg�@@��!�;qL��
���9������"�>/5�D��Oqd�ުW�!�y�@3���h'�5�E�Nz��o6��b>q�C�̈�}F�j��
DJ7�F��1
�>�[��7��*�,�)��	�}ͣh��<`<>%y
<���>��P��p'�,e�|v̥��#�UW�޲/��d�A5Ղx-�Ջ��:��2[<�x�����~����i%g�NPo�ءc����z��8aZDQ���C�*��z��P5��h�u�x�?�)k�,	!���}+q�#X`(��f��YEit��ޚc�J�5E�uk�oX�~(�����1��4>�6�g�Pg>.�D�=��l�Z��HA�����V���UiTIU{z����nUKL&F&�'ݹTV٘�m몈����")���E!�@g�#}"!0 6X��1�k���@9�$7�K˜b��5�B*t��8-�{|�U$4�(��c�7ʑ�C�m�pK��ԃ۴bR^��8��J����0��^����\ғ+d5��,&�3r'�)�2']���a�$�!&[��(T��uY5��E��k�G�i4CT�.������[�=��؝D}��D�n�L^ܯ�O��S��)��`r�E�I�M����w!��Ds	F/5o��$�R��uOr�9��[�K���X첄�����-�E|1�S<�E% �.�GR���
W�J��c�_�H,�l��U>f��3L�h��Q�U�u�×�"}�KH�#�Z��ǀ'��Yf�.0��U9���q@�,ɷD�n�h�;k���S��6G�p�cWUְG��Z��ު��;Ä�J���ML:�3���Z!,���K1i�z�-��%g���E�r��j�U�4�{���z6���r��_��Va`sid?T��CD���%�~-,� ԨZ8�t�[�>n�L��^gL�?'tZ�M�AxWu�W�)��/�4�L׺F3#J�<IG�vIY��U[-i����_I�`	lVO�S�G
*w�_y��^)�����D̤|d�/��Q+�e��>7�Sh�|�}f���Z�8���ݡ���2
�=Y]�Ve��~08�0�bW����}nȧe�~8Tl�&�}�.{I��\�V��X�� ��:���öB �?���DǞkE���@�B:�+;q�{��.��+�b���Е�x��0f����*W8����WI��N�{��t�<%F�V[�S�<�����A�S�����ԏ�U�d �1�D���ˌ��焭�2�OhcDBR��4ٳY��IYKBz9��'�8��e�3'��{�={�>m5/�����gZ=/��C�!��f���֖J6����%�9+&�J��Y����*��zgXr%����	/�i�탇�t��X-!�J�eU��+������U�d:�7�sK޶��������g`h���kP>
z���y�~�e�]�47�?�v������2@On5��1�o@WT��1�,�|�uy]����D&�@���~]�*�@~Q�(��������K��o�p1F���3)�.�<��x��ِ�(Q�pG���_&#�g�×�b\�Ao\ϐ�5���ex$��"J�'�~��d.8�;�M��-Q�U!����������m�����ju�uH��3V����з��c��Ӵ�X^��K{�N��?�fB��� v�T���+P{�3G��J�r��E�X0��_J�����|�r��w3����
���z�.�g�����fF�b|��N�H)Z{�yX���Yӌ휬�C|g[�,�y�Jv�^9a���"/"����m�k�1DC����p����(�8V��/Y'�S^e�[�z�%^Qk��\��X��L��_CA8nҤqCm[�����rB�f����nI�w`��A�f2{j�I���7{����� !3����WW谵o�
����.��4�Ib�� 1�fG�w6��I{/Z��,.��8g�<�;Y�]Q��ܒ8�D-V��5����Z>����Җ�M���kW�w�W�K%&'b^�煓Ȫ�$*��1��,�D��r�ֽ3ͨ�CU� �,Q��L�.��.�u�@��6a��;�ha=P]�8Ա`�v�����L�#���2c���UŃ��M��:4�.<֪�ӧs�D�����`��r���&�=��J��5��	�Z' Ư\�@��@�h/�4�gM0��[���i*������$��/�2���5r`��?=�����ީEu	��2��Fޓ'��h"&*����`�0H��p'D9=�/�[�<��ю06�a� �2S�(���T&����N�(O��9?x%)��8|tf�K������WZ�V��Yv	pO����Z�;t�(18gǭ%p�  �x�h�^��L�L͵��N%l̤���l���	y0���ʉϬ��������F���6�vcP���;�1�x�"�G�|�<��.���J����vT���M�~�DqG���2?�Az����#Lb�8Ip���Yô�n�ItU"������`�#fH�9�=��<@T�(��5���I$X앷�H�ԏC���]e�u�cV����颪+��R��A��O*��5>%�XʇYJ�b�|�~���q\��4� �$]����� 8%	*B	�l�7�#��D�bn������t��*?4��ƕ��Uԃ���[��Jx�X�̱����J�EQK�~�#:���w���p6�7�ę1-��l�o�k�,�E�3� �m��^�rDy�k���X�!@��
��y��V҈l�/RP�~�j�;��Ȧ�Ԡ�Qf2�1�$�>^)�ҍ�Ϣ�G�5������t��7i�j�w/:�CX�l ���C��u ��M���C����~��JRF��h���ףu��J�(�n�qD������2M��yP��Mmc�@<#�����Ub}�a(�Zz�[�� ��E��Q�
ݒ"�T��^�[��@���0����<v�te*Z}��}��;&>(��e�_2V,�h�'��~��n ���`~�n+�;펬����{���.m�}^��o�(%+��>�]l��sȼ��ӻW�Z>M]�3c\��U��b��xb�?�:�c��v�rX<� �$�Ń��|pv�FB��/N�m �>�C~�$��qe��9��\�S�F�n�ۦh0�K����0�ĝ���W�/�M�G*?uc��*G��>����Q�����Y�
�W��!���lu��T�tt	u��b��l ���<�A��s�\�P���r��"� _�-ɬ�5���]S����u���$�[�]��L���2�:����K�����Q���qG��N�4��k�f���`�^��f\�1�������y���Ԓ���$sNnA��8}C8�U.@��,�;�#2��ë���N��2?�"迠B��=��s1)�8��L`��<8�x���sF�
�y�E��m�nC �hDQ�E��~[�!��ݤ,�_�)����\��F(�����@�E(�Щ.�n��pp4d&�l,C�?�:��|ŋU����^�\1���K?Jf�����4>�js���Vm*��ŵU��C�ѕ��E7(��S%H�bH��x(T$`�y�]�kLd��@>��]V/`�7��� \D�h3���"����QiP����	>z��8���Z��0��������Iz�=�A҈4�n��<X�28L���?],���K)}o�]�?u�C�ͭh)�����'��Y�DU�F�epF�4E^��;���b�:C�׬=�2��2�B���0��⸩��s��-�����$��g�UƬ�h71��%U�6a(��k������څ�o�����[R;�ЯщViNK�5;M�ޭ�R�F�L�kSZ�R�vMԐl��,��0h�]n�����<�����p�Z��^��
ަ�r��L�&j��3|ӑ�h��΅�UpI�FY�:��M ;�?>q|M9C1�C����'�p�ݚ7�o�X/�C�R+�=�W)	��m�YQ��J.+$1�X����X�+��I�s��̭o�_����ۏf����1g�a�g-�L�N�VǑY�yԹ����B����d����-�YI�}�7�{.��/�sBvw�"+:3���V$1j�|�~e���9qгS\b�F�~zڈg�y�0Fۏ@�7���Ը�����j>��e@%����/HiP����.�w|�DWE�X��ԯ�A"����	�||�\��%�kHI��ߗS��;�'�v���E.Z��H�K���
֬�QW�By���Yo��ǲ@�۔�F��/ٶ����$��C��뺶
c�R<��J��9*��������<$�<��/2iz�7��)SIQ牢_��<a^��M�:��M���
�������B��$"ⰰ-�Ü�ƹT�)^w&��4�'�.��Q܈n�����A�$��A��셾3��h=��(V[�_�S
��/Y����A��-���|�GQ�E�f$�;@m� �}%-� 0�9�J��?���ć���*́Ƒ�fqzE��q%m�ތ!|�>�R�� Z�.��#:4����O(�/���e��o_�Nf�� �]NI1�;;���f7Fj���AБ�;�S�͂'����y
7JbͷCnϻ���CU'Z�����Ղ�<^���'����;;@����"� ����ZiZ]���B��@�!Qw�2�ǣ�	H�u�Θ�H&�l�ؘA�E��?�����t/cH�%1�kf�	�� �kB�FN�H3#�d[C�]?ϓ�&���0��˩�`��i�L�;���>T}z<o*q=��bN,��(�����ϳ��C=o$�]�wN�gL��$8Ղ���|�\U�S$�`���W|9���C3�]B?��K�p�`�TB������S�B��������n������-��gnc>,,�� 4aɿ�`���m=��c�)7Dq���|\�Oh�I�}K�_��.uNe:w���{p�(Ң���K�s�"+&�C!�/��dw�ڮ��DBU��b�ಛ'��?X�9_�<��%���}Lj#�a�Wş�F���W��lf�}O]V0�,���Qj�j:2�#f����I����f�u�m�J����¿������Ă[&fZ4�p��I��F4�_m@yz �Q���Ǆ���2`.'5����r�| ���R��G_�Uc.��8��N^ ��hrT�x	|�� �aR�T��V��%����.�)ȍ� �����kχ��ϼ듦ӥ;K�@'|I���	eY�\Ʀ����Pyy�X��4�P��]�$R5�
��)��(�_�;��n������.�V��1��i������> �����w�B�u[��1\���e�#�@�u����P�	�8s(��yf�����i�eQ�xY(����#>����XK[���%k=rnc)2��g�b.��tC�'w&*���P������am����ln�7�M�JK������L~1ױ�����AVO԰%��'�����(���~���v��4��]A_���h;��Ͻ��;�!
�p:��W���������	q�0[����!���"Kr�c9P��_e�r@���+[�_,���N���f��EF	�r�:���	1ʉ��Β�@����G��$òp��#=o�s �pn�$g�2or���X����M�u�&7�*W?r�T�ˁp@��p�R���Ȯ\^K��2�dr���,%q[j�h���R[%��"$�TR��}�z��ó:�sF����+!򃌖���8��=�����ؐ��:'[�5H�eO~S�m@˟nP�������I��d�B8X�f=�{��@�+Χ�qG_1ڼ�$W9�Q���j4��3u��P|Kݜ�%�V��wy�����2�s�&:��{���+q�$i����
Y:1g��F��H�����?�\�E&�a˯_�R���K�Άv#����d�K�SP%���i�z �����p�w&