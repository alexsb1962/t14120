��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�Lژ�O���3��������F����Q?���b�V����Ţ� K��Q�G�D��i�o�Yʫ�|�F�V{:�� �{��LBB���Z��^sӽy/��[����I����k���'_hx\�Ƥ�?���ƫC8�r��j���?�[�b��Gk����s��$E�C���Iv{��Ϗ.��R+!9u@Gf6�e+~�7k>�_3�T�@�@����58fW�o$�T�h,|���z.yhb+�[��>���W��Oѹ/t7y����8�A?X�Xw��J~���k.W�$�'��(��ꉑ'[J��TF�S���o�z󷬓�I�UW���{�|�M�a���@�F�J�Q�tx�tEV��Z��i��lzt����#��I ������T0�=C��'1#"V,���)�r����4p1����Ɠ��LS�d�,BbD�י��)�@/
X����0�9�C�'�8�5��I��*���ŀ�К�;R�g2�9B}������Qj����F�5#,VF5~z�wY@�g�ږ���jbY'��&W���Q��p�>��@牣@N�#���Up��]���ߏ����\c0�4i���jK�tƩ�H-c�����d�@+�FRxY�,��~F��(��y���^�)P݈�k4<�w���Z���?4���E�}��_�á��š�0ޜz/B��Ѽ��#f�݌$��3��z#G �W�fĨ��H+hnؐ�&�,�Ɍ��9�ċ1�(ֱ�{��v�RF�T5r�����F6�}6��2l����Ɯ-pw@���
�O1���3��~1��І6	��v�A���@�e!����� S-����193��n���2aD��T�=��2���;���(�
�^e'�3���;ó�p}�a���^8H�@�H�=�
�/�����=#��J:)�&Z��x�Z���Q�HD�)bD�kk	Y�Z��`0ꦗ�ɷ��{gr�_s�ԡ���Թ�3�e�����lC�Uw3�D.")[N��=֜r�F^����d���_�Ý/t�G�S�D ��"�U5�΂L�o�A哑ːr	ڭ�#���H>��8��������C���,)�C���g�_�,�:mvi�<��doZ�K'�[M� fJb���Ν���H��B6fOo�'	@��_��&�05�IR�~^f[=�B��5�Z�Bdw���gf����Z�Mdn�A��ͧ_�}���@��(pO�H"Xʟ���2�xw�e&%T
&�5i�	�M�
���6UI���&e^��<:,�h2�5�Q�4����Z�ݖ����`�F;,M#29��p���8�m�j��-�/=)��)��!D��.S-Ms�m�Y��Zm
f�l9����b����V�.�@5���ƨnF�!����/V^
�tn
\�;ک��A��j
\)(֒�V�����S���M�r5�CQ�l<=-4��e�U��\>9��X�Z*�ލ����EW�)D�鉜�3;���&Z/0����6�՝��L= �Gc�EY���{6:q ��?�L��r2�H{�ߜD�z��_�0��ݙ���bE����"������h۬�q�H�	!#S��AyE�}�E^�2>��L*�&�l�\�Ek5{>���Z�@?����)�cuf�evDB�V	9/�ERqw���j�A%Htd=�ę]�N�N�,���>� pDt�4�G�ʛr��aeL`�v�S��
�\��q�0�~�m�E�ծ����B-<G���Y�lԓ��H$�Q*~e�@��E����p�U��
tcn�]9;�SN�_V]eXbIxs�`*֢)������O����U�FY3Ɩ�Q�E�J��3J>�}ޖ������Q�$C�:���m�0��sO	�K���9o���ߌT�4��H�H��K���;��I��@9�h�\>��w5N�����g/>�kIq�n�,
��{@��3~M1�:gF��Fz�D�ʓ�Ν*�SҶ7Pr�W�{dP��G0��R�w|N�r˽T:��1�`����`���Q�N���ub��L���lcׄB��=�Ԓ5,�RC�
aF���~V��{���4ZhW��'��Z��)j�l}�]�y������*P�y�sg��a#�{���`