��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:��������uA��@��y���<����xDET>��W�����C%�=U����3v���hj��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\����J,�'��i߫w�+��J�\�܈W�k��ɹC���"�a�e�7^F�d���m��[2}a�����6&���)��ᢆ`�"
RC�U8��_��0@	�HyR�QgB��-��E����x a��gJ���A�K ����ɉy�Am��X��2��Yr�+pd<��\�݃��H
u!q\��P�]��c�纐��w���7���f�Vm����dg���LF�S'nc�|�t��
�%�Ut� �K�p{�u�����4��`nB�$���^�٤���8��❮f�$(޵�ֽGviϟ�#[ ��/=LJ�U�;6ô�Fbҭ��@A��s��<g�,�:�\ܮ�_��{��#D����c3�`MI\�M(U����<�X��Dj>�(*?+p"�ȉ���=��ɞ7C��q�U.�]y]��_!�ɑ�0��΄���84�Ӄ��1�4���RrC����Vd�/�|+m#�=4�up��G��b��Ԝ����E��߇&B+!@�q�_~�+�EF��t�S��MT\@Yۈc��R��Z[����8CK����	�u2�����]6sR�d��*�-��f_.����X&n�	�`�/��+�R�߷3����>|$�"�� k� �B�X;��-�'�B���\�t���X�u�br�,ߊ�&�e�A�DHk=�U���.�5��Z�}F�"�c���-+�z1]��:(v�X���E�X��q��ך�sHQ�������Y�X=D�s�w#�sbê�A��Scu�c3]�I`�
��(r�W�Xz�#���3�'�U��o���q���9}n� ǗG�"�=,O`����xZ.2!�_�`Y����%'t�&VP�A2Aq��M�iL��ݥ�2Q/4�"
I� ���ڙH�^�K��#B���.�խ���Nl� ]�z��6v��ۉHR��Ňד޳����D�f0���y�9koϙ�>5V_��j���_!�Uٙ��ы��v� �x���^����JX��
�g��	��b��JA8�֣�-`�L��6��d��4��	!�Չ�S����\����?�7�`Ly�#HNu���^�]m+ڈY�N��w	Řk`���H(�E	�K^1D�v��i�(l��#�d�U��I������0�� c��Ri�D{�E����¶a�#��}<�v.�D�ݹC���(�)�)-y�[�_OmQ�S�-A�Q��⟌љ�^a]�ܠ7ҵ�#?=���F�~F�� �q��� �9�C��YP����r�w�k�]��dD����ww�������Xk�qkF������sfp˓��zCT�����ut��N숽�L�����m�a��gI�/6�u �����V�s@T��'���`�s�������H���E��ۭ!?���\/�����׺L��U�5��ЬQwFL��Y��&+��m���ޅ��\h�Hˀw<O8�oD>h<�E�g��¸�ϫB�s���Q��"h<ۂ6tx�����%�(���N�<��A�9��`�r�Zʨ��oy[�'~�idN����P������U���k�4�j��Pa���=��W\�2/$F�5�]_���)��Q��%b���n�]X��\mn��G.�ԩ����3��II���O�͓��b�XIV^�5�>}ڶBAw�'q�C��`&̗�ES�J��I�ʤW�S���ҪV*`JA���3�lO�K�٤�!���Y���p?������߃O�FoQ�~4o�X���%`��2]]VK�E=Kp�X`�)�9�[��fr�ujo_���H����d�?Ĺ��'Q�Nz���~PvPi�+��X�{���[���Ƴ��5Mޏ�c������I
ô����@����k�jP������|1�A���Bp\��zy�����H�L�Ę�1���m�7�4f��W�+��uo��va���௞Ҽ/��$�8p�'b�~��ᩊ ^hv�$���e��( 
��
�0鶨�4�r�f~w�+��*_ǖ���CC6g����d�B���$��Ycװ���"D=��g����cD�=HQ+����T�ٽ��~�-�z�>\.�T�S�.?�='��q��jy����6�4��4�c#���Q��y�x��v�8g�G�t�<�ϟ�����rG�F���?FF�Ȁ8�`l[��>W�+V%���蛍>;R(�5Ղ:����$�,���ڦ�H
��������(`p���i4�W�#�Pϓ{��t�������,
%d��Y�.���})�X��P<�R�<m�Q���O�i/	�����L3�#[��i#��[:ڲ��3S�僩���Q8u� = �S@�=��o�K����!U�R��{�*RD�aގ+�Lq����?�*=�����42@;x]i��_с��3�+xz�`�Ҩ��aH�#�À�R/ ?)d�9fA�]�JJ��v��V�KŁɠ�\IWm����-�3O:�+56����|�`�l�#��D�e��$��(r=@2���q�Ȗ�2�ۄRQ���Єm5"����=�vgC���l�E��s|Ĥ�k�~�X��1a��=o�K��ɦ���]8,	���P�{����a�+ ���;�4�\��M84�t;YU�3��@��tX2��T�\48�#%a�ED*��}Z���B�n̿zG�n���7\@,�G�76��Z�K�.����@�'I"$��P�$�;X��jP�C�oUx���Z̆��gdѴʤ��+q!�&C'!��*09��{��z�'��Nn�~4 �� ����hX�s&�	k�Y��?�ĳ0��1GK�$欩Ml"�l]��g����c����(1*����:������#]�6���$�!�Hz��L�h*�5w�*'a@S`�D�㊎��Juvv�x�� Z�4�+{��6H��]����԰��ę-���/�剤�MB1_֨�F;r����YyU���ͅF��K��-�~6L��gթ=��P�I6~R>����#��<��j�D,�o�r���p��7N���8�����]����2D~
� ���1��s��p��_�g)i�����ު�2��U��������[�0$��9,2�>?�L��']�ǥW��VUv4L����.%�u��;�@c}E���?�i����5~�MB�߁��_< u@���jV2/@US=O�P�;�����7)�B#�x�Ee�`�<���7�F�Qz�yJ��Q�EWٳ��ګv�����A~���u�z��U2��rc�i���%U���?�����,�3,�U+�U5B������C$�����8����S^�7�����&�������G�$V=^�[����b6ti��*�iάL�9�s(����h�H���Ȩ9a���mv�Z��Ury��B�H(����].�ȝ,�4�����ҹ��#yd��Xd�j֚�Su:�8j�F�:�&p�#;RUۻ+]�Ǭ '���K+Д�K�!C��t�ٵ�f7nx|Ŝ���W�u���-�%�+$Vwɲ�"���46���%Ο6�T�˽]n�z�k���"�tW�S9iXճ9[9P���W;)�|D��Flp��鶁�]lv��A���0�_*��Կ����F]�
ܶ'`K$���w�S;Rʸ�Z�����0�-Mj}KL��*��2q^��L>j�(#�]���m`ٛD��v�͵[C-�:����������!t�)���DGE���b�u��Դ�$�+͏/Q���T([X&��G�����%#;U/�K�sɲK���}���IYES�rׅ*�r�7Rj?H�q ϶4B���� ��Y9V@'6����{����W�ꈃ��Wϋ�L ��M1�ڍuA'h&c��g3���t���>�w/z�2#���R!��p�WC��"��?��^n���mo���Ӏ���b��b��'.'�,��x
2�r��.��uǁ����[��\،�A�v�I��?[w���Lb��[.(���Q�s{��=)��{[�l�
>��~YHyG��v�%�,B"F��)n��*�c�e�(�N�r�Hj[�ۂ_cu���PncG��=�h���O|�i'�NL�Ҷ�Y��'��`�OJ�X�,�+�<oF���UYOH�l�����,�9мM�O0`��Ā'm�d��(���-�m��j ����Ox�+�^���VGփ�g�B'-*�w��1��t)�p0^�|xF�@�wp��(KhY���r)Q�����́�X�.�$�F�:S��*8�X.��_ǂ�bMX�#
j�iY��.:�/�Wp}���U	=gA�Wz�~p�v��	��~
0��H��w�V�w_�Q�W�bj*x�P��� ��Ȯ����e�������?ٌ�T� �<wp`Q��!��&�� -�&���LR�˞���^y������J%h���~4c'Ŗ���`�B*��HKߨ΅-o>�<����Se�3�lH����^Ճ�>���j��s3�P���v�@���ő���J`Д�TeFb���P�=k/�`�-�h7�I�O��X���JjFa���X��5�ԟv8|,Q���,���}Ȋ.\���Za�Ԏ2mW����/Z:�68�)+��nh���ޫ@2�E̷�dg>Zh#m�ך@��H�}��NJٙ=���z�RG�iY�I�2�GGC�;����4�����>��/��p�ƀ�X��n����:�Uf}f�a���t�,с�w�o���Q��ܖ�+�Em�����	1_�����ڟ~sn������m�݉��O_��e��ɔ���
{�`[!�S�� U'v.����g7C���� !�"��0��H��A���N �_\M&cZĚ�Td�[��-����A�V8��#�!���a?���y9�+���ۯW}�����3j6�tqgx�~��8y�B�B�@��ɔ�L.2�����B�;�DM¸X�']��=|x��O	3V���[K7�ń�y<��2�-������O
(���Ɛ��5F^_�,G�"���!���*Qo�^$�{Z96��N��4�K"�Yd�X�D�Z���9�:�~����O�вZȤ��9���U����R�51���/9g&����1&����M0��t󤙧w�Y���|V�Q��Z��pe�����bX��{��Zԗ�h�
]@�ݡ!G,�չ1��\L����w�B����;�w��b�=I/�U%��-�w�o:��)	 W�W� ����Qs��Ҁ���0��?�I}���Py����𨏚+�X��l�X_��jR�UY
a�I/N]�ɂO��9�	WUޮ�?>��3vR}�`��̼t��N/����1�&��<�"A�:�+�V	���S÷N�zD���Ֆ���;���`z�ȿ�Ы�K\�W��l��)�z�8;�HQ(n��~�T:r`4c Pmpwa�/�U �
T���P��}�v&��yQ��o�Fe�=o}�G��`��E�J&�g�����P�`S)����Fh���O�<��?���������~�i��7���~P�@B:;�3���*�z�		�f�0�c���+���f�1ޑ}ݪ�^���<���,�fv��A�d�{���v8���w�����ԅ:Z�Z�����_��ɵ��ܩ.A�8ť��F�#���������=�Jv��3)��5���M�P�\vzg��!iBh�n2�l�A4� ��G������|ZT26q�B�X��f�3�6�Xp�e]��zX��^R�����'�����ݹ��ޑ]Ze���T�	T��܎MI�Ϝ�b��d}=��G�����wO���Z�+��^2G>5�S=��$L�'���$d�5i� r�20W��t����쀩Z|&L�Q!L�Ɉ��2�f,�3�;�7�r"C��\=IK���6�;��BnjOYk������P�B&^p���+���4^@�"Bn�3�}�M�i��Dʎ�K���E�.�7�!��bEQ�uÍ���E�j���QGn��D!�-ĳLOYHm�ߝV�`X�l��i�}��1�N<v��dvţ����;�x:��4��y�\=�D"��n"pZ,��� �O\���D����R�^w]��Qr�X�>��Z�,��c��Bw�X�ห��x�\�BT_��Š�4~���5d7l����fw��3���ۏ�����¸`@�W9�k9A�J�?!ép�4�	��*/ꧠ�<+�=�$`KU4]��-Ot?�%g�K��9]�4�NFλ޲��{���M˧��&���z�i�� �U�ӵ6S��"Y r�7� ����)Ў�$�6��8�~�96�\�PSS��㆔0���EH��	��z8u'���O�%T�H5d(����4�`��~	�;�Io�~~�����C�]f�3 ��J5���z%xCr��ogkgȩA�A���lU��ð*ɚӞ?��q����VE	���;y�Nh1��{S4
���H2q{z�l��`��pdv�v|�N!�S_x�	?'��yMbڰ_p�m�D�A�<��O�,Ľ��/�T�l|zya�'�
�����CQܷ�Қ{�f�����j���R���6풦;,�:Fq�WTs�pߛ�����A���*�������{�Ƣ3g\����!\㯎�	?s)�i~�[�ݻ���˯��8`;|S�v������;���~��GMw/8b�z��`�^8��1� �]`b��T������); M,�R)���&��u@�(�~��R��p�QK��$Вp�f���W�6z��h���t]�wJ%�s?���a��_+9Y��_����_��X
��6�ijm��x:�g+*�FI�Ly3�x��'�gb�Yp;���<hl����A�y��"��N�N%��?�y�����`��E��?�Į%Q���}{�'m����?���3-�l����f��Yl5Ǜ�B��������G�B�2zH������P���K��`&�㩫B�[�\����͑���z�Y�)���#���_��}x1a7̋��X`L� ���Q�^��4�{���)*��<X�[:�5�_&��Tåi�݈Bÿ�4G�qa���;Uj�J����C�z�uu>�$ZH�4o���;N\1�ڑY�H��Oxc4bb��Z��a�)	�ʅ�b�fk��?1�M�K��-�w1�mo��>5�2��%`5��VST��2�"C���Ծ���S�39^�֪�f�]q� j11,B�"$�_P9�v��dI@$$RA��B����<Ĉl��\Cn���v�LӒ�uV�x���^����}�Q�������MY"�Q���\����O�Gq�/��JTq���}��f�2>����x�M����K��·Fg	�C�Y~{�
�P[���o$u��y(����Km���`؎�1@�Lg��(��~��/Ⱦ(��ϸ�"��N�j�H�sU�qip�a���&.5@.������..��D%�=�t-}� *ȣ��7NEߒtB_d\:��1��Z�jnDiN����0��b^8`�T�yyW��V!�r{Dh�#[ki��S�I?c��M����dZ�lv2!�1�e�BR��x@y�\�-9�^��������U�	���HZ{�6B��H���X��6�������3Ϝ�<7��ɠ�qT��cޜ2���ő� -�����:����������sJg�NC.���������(���(S�M���������rc��9����h�$�O�&a��D�s+z�#�� S��'����!�g�Ok�"�8�CG4-x��T��#�\2Z�v�*�v  ���?�]����]����Ma��>x��͉�N�%��0��F?���[�	�zL��H9\Q�.�耴r�)�M���$�Ca��.������pR�2��畁����"���Q�������˧��|���$r�ߔghm��U8C3�Y�1�Ҳ����^?�i���f��|:G/�9W8F��N�.�!x�5���Kѡ����j�%F&S�R�a8�J�!k�����79 ��V<�Wl9������8�=Z�aR|�$+��t���ֺ�`\�6�F�۔�]�++��[4�Z?bj�+E��<�]�=ײ�� *25��b��P�V�&bK0����ه�`��K��$����#�.�j�,���e�VG Ul	=����wi����J�$�����)�s*mw���Z�7�����m��")�����"����� �C�MjU�qg�����e���o�����V������θʦui5gV�s�N��֝T�3M�pm�����B�ǰ-����.����J�1�I���'4�8]A�|��%х�.�k�$MW�/W��Vx�*�x|�$�]�K/���a����Pr������Rs�)���<>�@�Y��j����&�Ï�پ�����˓��f�'S�P�\g��9�J�������bu�_�w"�,�ģ��`Q#�0��4�"S���=w�.Z>���-��@
��c�eGIǱ����.oP\A����D�m��k�yt��B�F"#����;r��b�=�T��jt����O�>�r�n��%k�(M��$��V�J�K9W2�����?g}��h���I��0`�T�rqTL��N�` ��榠��%��!�5�P������u����O˜uo���i>�رv�\�(�ŏu��[u��1Q�H7^٨f�ϱ��M'{�rX���Y���Oߏӆ$	�3r���s���A��d !
�6Ԅ�����nJ�>SX����E�U��?w��K���	VH��ZȖ�]#�ʛ^~fV�6 �d�]��]�q(�.���KFT8z{�OS@G<�dc��w�q��� n�����RʐQx5��Agj��nv'މs.q��,���ls�r~�x�k��'ĉ Sˌ��&�h"��I�G9$q��>�eY�<���P�'���w&�۔�|ithU�y3oX?�_@릞ōVyޠAR�r^�o���x׮S�G��T���F�``��\��T=��4����d0�z�_l��a�1K�7E���v�ʄ6����Z<0��Q?����*8����E�?7��D@��O�ʦPSY��f���lLc����d��L��,<��I�:���]��B�&2_'y@^�m�d�A2��`�ɥX�|�r��8�j	пAF�s�I<-u�@���9��S��g�dL�e�~��9�l�5βa?�oL�>b�L�H���9�LdF�DE��q����Wi!;�T��}z� �IX��tx:;�o"�$�� ?�X���s)����*;�4�>@�oEŕg����c^@��Y�r��(b�+\��=]_�������3�/&��b4��'���}�|���o��P-���n#���ՊL#|�C�KW�br��-[W���d�P�No<�͹r�����PW����eV��c��~���1��o��o��HF�s/�=̅o�������u8���w�YB�4DQ_o���X޷��pJ'���0Z$5F����}5����Q�M��UP���ƒ�Z��>e2�y͇��VT��i� Lx�����a8�M��-�E����Y�R��C$�$�+�\�
JPa
y!�wM���[�]�3u��H ��K�!v|s�z��)|���jN%�)��|k����Oܚ8��Fb��B�&-_o�p}˜I����ٿ)��IIɵ~���$�U�ȥt� �3SL�%<�y�>��*I"�$�X�'pT�	��g��6N��a��C���ƌꮲ˘�<�̂_�����q��(����Q@ސ��FB@����j����u:�|�I�a��EDz�����ps�����uɨN@��Hl�&|��ﰭNPˀ���2CK�f��CNU�jM�뵵������]g�k���)H +	��7�"���
�u�6�\��!z�7��B�fl4�`�rF��w�E����՜��Ř��(8K]��۵�w� �ϓ%Ys��ۈI]y)��8���q�9��r����h�/'����>�fW?5��5Ш{��DJt
�6�@�g��*��W�Z�i��6���M(+L	�1��ȗ<2evb�l��qco��c����]�p2�=9����!���������
�P�ҏ	�����t۔*tQM�&�ȂӵG�\��_�'��1Z����F�4`3�ON\~�~�y��v��?�%�a_��bC>�l$#�ڿ�d�[�
 R7���V��O&L`᥈�r7��Y���ͣ��Q�f��XK�pL96�� 7�ʶl�6 �Ԡ6�O�eU~����M'P�b�*[4�o5���d�$/O�[b�i*R4]{�ۀ��97��B �7�zU=@�˪I�/T몽0��S֙9=��,(Sv�d�*����S�ʁ���'�#��H7�ʈ����ו`��zL8���CgG��-�$�bAz�' 7����7K�l�ue+��2���|�>1?\�|�0_��_@)�<gx=Cu N���(;�
���~9�~)��aˠh��ìYH^{9*0G������/�zh<S�qH�0)����A�ת5A�Hg* �S ���yg�ܰ�s#������1�U�������'ߚ��o�Mu����^�3EE֋�H�t�7\�pyr4����	�w�1l�̆teD��K�r"F(��<��@���������X�x+m�*u�-h|���e�?�Li�Z�ϰ8�{�G��U�#T� M�ÿ_aUQ���ߔ��ͥ�i�]+��	_&_k���ʻ��F20�?�������&In�)
��_��:k_�^L^������)9��+��}@��CPL�ʫA�;���{�R���'e����&��ʭ�<��6���������)����D�ۓ�����U�~��	���NQ�L��ζ#���E$p v#�b�A�ҍ�6_F1uȒ�����H�"D��;D�_u(~�����q��K��|#�٬])��l����+���-�������n�������*C��u�_%�p?�V������C��H"����>I^��_;���i�Ot �e]�MG�? ��޷���[�4����pe0vz��۠A%�whp������˂�ީ��.����j%ђǡ)��2_�[sv�1�\`�Ќ�����+j����OA��3M*	_�."Y�2�_�����G��%��6G;P.:�C�]%:9�Oo �)�����7V��]G����#��]�8��֫u)jV6$w��
m-��9T$������>�e��Cm�<�:�I�������3�6�G�pِ��33 Czu
���i�X>�ۻ�������>L�ü�e��ܜ��Qa�U|�
��޸r����4�ri}�%�����a��P,w2�I��ìQ(�P9(X�ךѭf�(�W�Й�W"\�9�Ի�3��4oN��9�������4�U��m��C�;�9�4���d���9S5zK�����5۱�)���t�
^�܊��k�g�G�vCU�&�:�Aܣ�VO���(������X����T��%�"�=!����A��pq�&�Og>i�㙩��/�k��޷|�еj��,?T`�����^4K��Ү��['ˌ)�I�P��"WM�H���B���	�[�$��+޶p��?�I��{���Q��Q�_#x����ɘ��dd�Bn/�T������^�d��#w�u��%g��K�^?�ϕ�;<�����ĝ�P��f������N���K�!���r��n?u�|'=�ux뤳�T�ā���-f�o���?�@������x>�����ım���j��Jeg���kvQZ9�J����ln���?.�n*A�n�7p�a�$�o��,;o�1d��<ΊU�����z6�m��ּ8�X&Ek�ޢy+~���q��l��k@�_����J:���(����^�X�����ųS$�u���������\k�������ii��� ���WY}J���ݰj�$���7
3[WCO�~�R_R����� t^(�4�ܓ��c��q��ujAV�c=X�%�Q����O�r3k���:���|�W�z]CqU��
��3�=T"��<���S���Y�o�N��1�v��g�Jrt��us̍�y�,�d�(W�[!ޟ"dY/u��#b��nqA�"�����m0�Y�M����$�4����<i�� �N���bͮ@���<�z焗�& ���x�K���r]p�PB���2�B���:�;��1U7�>͆0�ǔ��G�[g��/�9#�LF)��h��KA��)��]Q�6��i�`��f��ڊ0X�8^WY���H��k�K��H%��z�;!X�l�_V�N��|���"�B�tE�m�q:"\ǘ0>���Z�t��Ǝd�?�Y�h�ۻ�!Z�g�m�Ԭc�T�@9�yP�+����C���
��Cl���5iH��Q�z2�!Y#�i���@^�hƝ;#��;�-{��aiK[����>]�P��]�ʼ��R����AV#�`�e�"�U����y�Q�|*��w.!��k��M뼒����z�i���R�Q���%�=����iG�#؋8��|�u_�`R����	�=�7��Q,S�Ԩ�Fi��I�6Z�����aR.���ke��w
Ɂi�w��`�C�A�P�FW����`�!N�	ڣ���N��T/�Z=X�1d=�5/�\�h��.�+2 ���l� V��y�7JC68�b6)�j�+d"uUr�Nt�ԥ3�	0�v�{�J��.���9ȡ�AC�mZе�<h�-��̑4!؛��(������3��$��<��te����\|�襎��5'���r]��-�ʞ�*f�,��;]n)�Vw�4S=�.����'���'�L}�{�%���vi�V��o(�c���++ISѤ�d�)j��z���s<(�u�~,�g:H��)��h�j!�h1��ޔuvp�%���O7C�Ɋ�(�{�K�����[9b7j@�_f�ˣ@��&\��#�,�G��,c��>��q8�,zh 1���G´�/Ϛd�ץ&`P���K�(+0�8:_�Es���*�̀�@�z���Z�"4�|���)$��UT�4�\(ל��Y��r"��=,iڍ\	m=���ɕ�~�3))y�q��"�}ׇ�#��"l�����Ey<��x��}$�|�/i����ű2�b>���h���7#�l���>c8�E�X������ropH��:7����Q}��JP������F�Ԙ7��e��~1�+�4�� 6�g��h��WKɷtc>��Z�I��Bvs�]:��L}�m�$���PN�wD��>fp�Fs��$L-��w�mݑ�B���# Y)�r����OE��¥mvjv�g{](�(�ïI
BW����IE�����>��<��=5���Ǌ�h�!����c�k`̿-M��m���i��S�E!�C���GOsAOd ļ��� �o^���Tc"i9}��_��u�QWVߴ&��5eHH~����X"7e��]Z�feB��nA�ќE�?;����|t�F-.�jC#�����:�.\=¸�}�{���l�q1�?���>s�A�5�G�d>lϬ�ps�[>j%��9+�z)���#�%�Ǐ*3���ɸ[�c�) y��ט~I�t��D��ݻ%�r�!�k�����Y^i���c���.6Vm�d1�� *�~3 ��X�A�j�XbW~�%���)cS�=�>E�bE0/� q�^,��W�^��X���'U�JU�R?{���T����ԑ�>�j�\���r�O�k'��4� �YC�;,���͛���60�d�al�$�c�#�­ŗ~gH��*	�|&?8�T���|ᭉ�G�h��NI	��9���o9y o0K�f��:���שE�K�l��A�)6G���и��0�����3�J䖀�C������ч93=e���M���s����C���_�����~mf�H�=c^a�c���3SY"�����ϯ�����~�'�����5DR�6'D܁�5B)�Z�.G��p\��x�S ���/Q~�l۠��_�N�ܔ�4�zd���t��t�D9�e~Ȏ���ɩ5��p#S�;
�0�7.�U�WV��]��5@�̾{xީD����u�}�|�tϮ6t
q�V�QJ=�mS9t@+��r���ٞ�XK�0Rpp�ҎZm����i�j��a�Q�YHK�p�ә��4��Ak�d�iY��0����z��n�Q�P���7�6SJ*�>�;��(��^�����xٯuT��@��L,*�(��ԚH#]�L�]�o;x=i�Q;��(�B���{�ۉ�>�yR|��	�h�(R�L��gkL�Ϗ\�,���H����� ��W�Y�wڶ�M�jl�Wnl���dj�����q��Kg�k\��NR��LYOX^U�C(���h�l���b�6`��]�������c0���㙗�+��u�L/"ЭS�w&N��Z�~X��7[�h�{���؂׷�r-=��V��u�Fxd>t���'�4�/�t[�I2�ҿ�+O'���0h�y���`�~����V�y�P(��D����7 ���-_�^۷M�)]��w VJ+%�]nޞ�������\NK�ZQ����	�߭����{�D
0ĝ� At�&���g�~��xaK3$�S��$�R�<(Qej�������ŵ�©&�Xtv�Z
۠����[�[����"�aQ���0�5��Dڹ&��\�Ӆ)�7 ��løo(�U+VG�����u�6j	YAH�U���lD\�g������B�;r��_�Ә٩s;��vއz��H�D���VQ�/~w�L�:�C9S{z�p#�뮫v�u���SF{�ʫ1C�%v[������P�/V\g��O�L������O^:Z�vj]�?o��8â�Y����;��rJ�D����G����<�߻)�� U��V�Q�V������g;"������ƶ(��F/�p�,�hoA�n�hh�5"�,-�Hx�����{������Ik�E�*�'�(�p���/s�h��tOw�?'Jsr|l}����o�c��ǃ�^�ܮ��;��3B����no�"��ĥPch����q���C��i�9I^ ԁ�I�M#�ZN(�he@�]��C>ە�������}$u'�LJYx��&9�Ƴ�[
�;���S�bD*��9,���7�5A|�ܠ +�_C]�[�F�)���r����Tj�xs�o�ۃ��~�a�zr�gP����U*	.�u�I<� $��-�4➵|~����\���?��Ǔ���كn�v䳌�8g��TM暭!?cs� ��Q��^��UHuo�`ͣ}�������d��)��g�==���o{�N��t�7�c���z/��2��-;�N*�N�N�<��x�s���|h���.x��R��.����\4x�IN|Β�isp�����~A��"+.k�dN�m�>����Q��`��/gF�jM�~���4\������a�j��Ԭ����NU�!-\O����[ӫB��Ks�m��0˫G�PT�(kۂd'v��/�Gs��⒀���i2R8��	m��p��C�� �t
�o%���]�Z��q�%U�P���6��5>oR"�ꡣ���[�~�;�γ�^��Ĵw���~ӏ3{�>Qwڛ�$�n��@a�8�5�`�t�zM�,�h�%O�|;1�ۃ��V�S�ɪ��.Ue0�������!���.�PbI+��F�֘}pl@"���~$��J
v�10~l��(��f*i2����^Az���3��6sZ����ln떯���'	4��J�����C�����j����=�'�b�̚&LMDy��kRfƨ���M�S��N5n���C�$|mE�O�{n�͠����S"rX�>$Ê���O�7�k�
|��W�Ύx�Ş~o�Њ1���c�磻f_�������5�׊-8+E��5If\�T�s�� T��B������(i�ף���2E�E� �s����� ��׎�W-c�龸�Y�ܗ�O$��d_��lƿY��BJؗD��ۘz_���N�zIh�� ٍ��T!�Q� ��D��]��#�m�=�ԩ��0�Z��K����H�~�X.'�2�K��𴆢 �	��bKN]��f$4�	��.<�%��mN�z0׿U(v!-�|,�>u:��L��E �L�K#���HY��E6Y�A�k���G�V쪤�]A�$ˊr�]�{�n�i'�aE'�#_�h" C��}���%=��6��B�@	�����������4��/��k�g�Ag����:o!��b
3}P�1L�{�Rc	�����bP��p�uwa�cthM���&� #������K<g��YG�P�ύh'Nt��$^�k��"�}�^�u��l�};�r���0e�lW3w�A�,g;�W�P��$���K�5e� A��՞TDE�5Խe��:�ō}����N?����Ez�����LH�)Ik3��ĘF���+'<]�HK�|���I̥]3\�3&P ����7����@�t&U�����P�f�n�������f	�!M$���87Tt ���gUu�Bf����-a,>�Q����p�_�h}�?}˅���]LnE�9��^�nk�n�� �ó���3=����ֺ���(�z*�����i��}0�]�p~��	s8���a���r�~P�͈Bl{��A�����7�R�(}�ӓM�|]]��!�y�C���ೡ�P���7\�I�?��F�B�_ 9� �ԏ@ަӊ����v�p�V�:2�`����3=-#�g�1l�b���T�}M�{Fg���Խ�s̪�>?�,�����r��{��%��s�D����$�x���~�r��6j�����\+r'N��*q��ㄣ�lh�b�#�ۉ�5a����(15��Y�i�m����/q��Hī�w��WH�̯~@����fqz!�����ǝJ�j�d�
u�;zP@�����H�a�6�t^C�nz�������ׁ9P��73ŉx��k�[6���͋�;]&j+[ c��3Mޣ�]'�ybδ7�]�-|S@�*�N�*��-�1o^o,�
����C.
3q?OBp''��e� �ȶ�Qg;���e�x�!g-Y8ƴFVC޺�>:���<q����y��Q��׬,�������SDs	5	��<Mop��c�;��:�K���]8�p�S����Ɨ��Mi z�_��W���Ӄ�~��W�zY�Q���8�\
��_y%�X팁L�.��0��"�*�_�o�/��@�~���=�=si]b���lf��W�9K�l��vS��L�ZGdͻ���7K�u��{q���l�����]���,���p��NXF��\��~�Ҩf9Bs��x�I3:g-j���H|B�r�c�*SzvP���� �L ��a�M���J=���k~&~	6��cU7�*ƏG�|Uz۠��D���5��?������'�o�����CB.\[��Ϟn�
C:�Q��s�"e}�ռC{��ź�4�}�\���&1��ە�a�؏��	�gr2%�6��E("�Z^�b_;���Ǒc-\��P!R��z����B$�P}�ͷ�'�`K|�-~n����=P�E����X�k̳�0�l"�aNI�ˤ���5y��#��k���� i�AE��~0i�YRZ��VмK�)[���W=L
�3������_ -�}-���#��ǯ�%Bt�u.�}���QJ��\�XJ�?��o�uQb���0ޡ����,X��X^��$ɾá�%S��2��ֶ���H.��w����؈ә�6F����R�$ �6y#��0���u�2������h8yP�T������rruB��j<�]�+Uؙ��b��{(7<}�u�c�@$��t
ݬ�ϩ��Q�eR��*�ԋ���(5���ɭ0�<�z�S�ǣ��%Gb�"x�L��`��ݵ�b?�5yd~0ӂR�1���C��y����,��=�r��Qއg�ܭoR�f&���ʏ�"(���J�Da���d��7V�$
kSw��9k ���S��tK?��&�Um7�;�xG6�pǺ�9��(�[$o!d�F�L��{O�����H6-8_��ki�	���6�칀G �)�M�YUH"�1`n�Yp� f�Lc2��FO�S�N��_���Ҝ@���%�p�|�DmY��w�W�b=��Q*^ff�cŦ)#	�_��Y�-��5������2�*�f՚��m���5��Nh�x1�v]'~&��l6��p��f��f9>�*�� ����39�Y�L�A+�9�r�O3G)1�`H�E6��]�N����8=�Z�N~6J�AJ���׈2��,m�����{��i��|���ʩ����dUTt	�V�D��_�����\NE�Y��!ʁ�l���y�/�k�ZhkE^���Eï�M�C���+�G;��)E� vш?I�Rp���mؖ@Z�^'�y,e�
������@�	U���nB!�@t�d`h.�Z}-���=Q!3������+-0��[k��p��2^����M�����	쫽3�ķ�׬͑ܲ�"��H�푆�q?�(��)�iz�]�@�6o��o �EtWpHm�
r#����P��қ�c���o4Q������K�h�J5�	�[���c��Q[��E�{��I�`!9v��&�	VLj/�X�vO\����}4wwR����x�7v#�?k�������;h�4ڸ�mm�Z���v(��J�xKX�w����*V�?����R���
�> Q:RQH���Êm�vp$%I�	�j��8��YQ{V48�?|�U�-LYť��>�o^��:�v%+<as]�5?(pW2��JO<:�"Q�*�<�����*��uq��d�\ΙHDc9��:|R��V��5�]s�+ZX��v�uX�P0Hd�9ҫ�+SJ���vҖKlj�JK�:u����m����;A'�u�Q:j����L
"(	n��	mO�]p�^�u�O�A^ǌ�U�4d�K��{�r���emw��H7X�	[�ޞ�L�q	�� I����pU�s\f�lh��f�k�	J!)�:C���e'�¶�Ү�v;����GUZ�C|�ɜ��o���e��T� �Jc^/P�/	|-�.h�2�f��|�����,���>FUv�_��Z��4��T �Zژ���c��L�"E���*�����Y;�7�Aޙ�T�V@��'�5���/����έ�i<X)�)+��V����b���(:�l1�i�9O�tޭv����A��8�� 5S��mU���0��jL�R]�5Ǌi�j9�.`*.���C�ߍ�A�|�8�9�<�Z��e��.���k������v�� )P�XbMV>�!_�۾5��#�!@�RWՙ��2�Οvԇp�\���C�ǰB��! ]�`|r�I%Ṕ}���h��K�m��5/G�D����ȝm��9�OD�H��"t=Lx�i�C��jWƞp�/u���%�&�x����]���l4뽺�(2����B+��"�nA7��iu7�"�ںa��Კ�3������X��|����>��\)5-a�Y#�l9|܂�i�P6O+���]Nh��IL�Z���^j�x -�����F��n�Q��w�b�[O�5� �t�\��� ��5f}�x9�D��'�w�9��&���xL�����Tm���?�$2*����1���'\9��5��9蹩��( ���h�4p!��N�؃�H��cf,w:��%Դ�Q��%
�T�0��To¶�A6�jk�N�\9�xT�£�7a�w-E�W~c��N] ��`�4�s�Bd���W �h�-��K���ʉ8���)��g�u��&�'����Y��}j��W~y͚3�=@���z8��GI�O�txV�=��w%kQ�&ʵZř7�<l�F:Q����Z�L�}�k����	����n2�25N�ɰ���F�ؓr�Z�����]��,�4o.� �H��)�~�z
�9yV^?���&_l�h@���*�k�4� �x����ڶ�����ە�$��Bq-�6O�-�5�l��Yt�VC=��\y���|ߏ�{H��<l��3�-l�FB�(�yQl��Bt�J�ix)���RO"��xs��O�P�ג���WLY�v7�}f4�|�Wb�鍎;���II.j���u5���I����.V6���i��r\���]y ���4_aX�mF_)ʆ$�N�����b�9���=�m3U�LvT ���p��(Ӫ;I�v��*5޿�E���]�ٔ��sh���q�����,˚P���#���aXQ[�,�0���D�m�8��q%��{��C�v��3#
L)��#G$+�a�����}7q],\6�+�(!�<0��Jl
�yd��~�;D80���z̰Ph?�-�+�ԏ[pJ����j�\�i��&s��� �D�sn#F�f�N'@�"N�[V4{��/K{uL7̏��{���)ꄹ֚�Y������v��`Z������l�6�52/��K׵zb}�i�l��Ce7��t'3�G��6vK��Y8�/�kP�eۻ�AB�)!�\�a�I/F��}2YI��〕d�c���o����~��_aQ���%R2U�� J��y��1�j^o;0R�,u0Ed-FQA�W�YM����D�\��.+��B�����L�11 `)0�v'DL���W�R��+ǆ���������*����k��j�g�@^�yaȠ�Ѣa�
E&��&�0E��H1ܷ�E	��&FG!��U��Z
H(��|�W�-��OS�0���tt)�x/5FA���ûl�)�z�b	zZ�gI���������G�˸�C;�.Q�=�~�8���9��'��Bh�o�[�����Yȗa� $m�a��#�����)����Mq�����=/}�M5Xru�"�~�E���*��ۋ�tC�i���@�D�⣵d(�yC�݇�n_r:ȅ���>ܺ���X��Hk������`����@�MH�IW`�����kv�.�B;�[R5�`H�� ev��0xt�:W�©�8��ome[���%���`�@d��2dp���9ou,�7�Y�������˱�ȼ�@��jㅊŪ�F	Ϙ YO-(��Ȝ��5E�ZB=�!x�5���E��z��ŉo�=��"Yc�����Ճ̴cJ����a*��K�+]�� �vmRm��z&nXOr�X6�с�8�7���F�'z���[W���w%�/x�{=7EP��W�����(�bt�	`[J�*�<#ӣ�9�Q�o8C3T���V~z���n������j��~_2B�L�e�m�k�?ra��	����<`�'o��C����:��8.�%�
di�u�Sn
�eЉ!�|��Vo��Hf�8�&ML'w�Xu_g��%�S�5��i�m�-xJ���V��/��O��9b��6*�p
y�&,�#��'�/�h��s��������^D��=��d�d��ʀ��� ������ی�P�����fuZ�.��Q��xAl�P��X6�oY�.|�j�KO��'<P#��Ȝ��أ��s�����XI����@�imbU>�u�$�%���� �����ΰ�;�8a�a?����BS�-�Lz�/�f]=+ЏӔ���C�֠�̝~�ʳ�l*�ERt��=ւ�������fw�����1�ům��hyG����Xy��]x�P�M8�B=��H���9Ԡt9�(^uq�:�b�u+vB�ҟ]{U̕�F�pd��޸�ǭ {*��as�Q,�Z)iGHP5���˚�Ak aMP�Z"^l��kA�s����f�EQ>'�V��qEk�>r���+�ݭ����!��2!v�zO'��:]����D��c}�#����Gk�-<�����;C%������������'�]�54�R��z�X?8/[��G���.��8[�'�"�N�8�����9L;y�~������Ҋ^����(&�ˢ.L�=|n��Wl(��d�
� �Eg�lg�[�b����2��q[ba������f���N2�XJ}�(��b@ ��8S�A�\�P}"�N�~|���F�a���l�y�y�'�=�Y����mK$�Ke%�,a���[�\b���,E��8�d�1V�(�`�"�j��