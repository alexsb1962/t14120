��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����pn�R��}�t�  ",�N<��;���Z��4d��{�
��|��Ȋ)zo1���á-�w~��d�<4��ˌ�ň��h����mo����/~.)��3\�R�F*}�c}��uO�������3�����U���T���딣0&_���X0���2|	p��rw@	@us������q�P.�U��h�`.yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\����vg������W�a���R���⪘����t�켻�S���c, '�yN�����8��U�7�+fja�ԈE�/T��  �ݘ��`��О������/��^���4!����Y�f��a�Z��Vv�c
����7(�(���2���oK���j��J"/��B������0�M�be8Wg��5F��(	��������E2ܠ�􋒥)��Hi+�3��������*��pcg�%�э�|�8��,\�x�j؀O��.��;��/�Ԯ)1~�w�i��y��}��@�dB���8`���ı���Nq� ,DEEN�� ƃ�J-;��;�]?Yr/r��\���7��(�z]ɗ���1H#�b!��u፮�[k�#χ������e���2��㓵@L�d�~�z7	9짎�����6K�_����6H��ź���f���ϹS �b�6��+V�	¾�-�t�3�K�O9��l����!k��T-�02bt�T���AH'i�P�EZo�]�$�ʫ�)���Uڀ;p�x�6B�ʏwU�'*\�y4dT>
k�����a�М�V����YD�i��]6�
�F��T�g��������yl��A�x铞E���  �_FE�:����d,��>{�i�C�˩���.|��β��o�W��Ls�Fޣ�����jF[s�AD�CJ�O��~���$�X 
�����&��T� [����0�Ee!J�nx!����%�>��~
EF���3��p^G��斻$�÷8=G�𿦗��0I$�o���M��m�'��q���E,�^����2$6�sI䮡"�N$Q/���7ތ�m�[;S�񊠓`�9w��{���鞘�؏���o���̄\�2��s��9������	]�k��,>&S�XQ��N���x�[oI��У��Z#`nVtȣ�2$6�sI�O��$�[9�S8a�bY#J;���A�\�2��s���|s�h���?��Ϙꛤ).�޽�c& �� dJ��l��
�%�э�3@�%���+�Mrt���448@��N��5I0��J��Z�']��%����j�?4{R�H�^9�?o��U;mG�ٓܣ�h�� 7��ӊ���n�\ӑ��:,i_�����7����˅EΩ���CY�樐 ��c�Euޚ$d��H'-������a�Ň�bos��n��I8� NLDY�P|�1�ljg�wʢ�E��S_��� ��o�}a�C��k(����`7і^�������w=��[�+� ���*5�$�Z�G�:y�}�zY'\(/�3��R�d�3M�$��fF�:aw#bࡸ_$�E�#s�l���{�	p!���?\����8���f��>zrd>�T�����V��߹�_$�O
�iC���Kʺ+c��"?pH�Z,R%��3�}���R�n)z�Z����2>�dƆ�Q;�����AOP(|VJ�m�<����LR<dV�kJ�e
aZ�Ბ���݊>8��/9���-F.8��-��b��(��[c�-�-n`���=m�K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|n����f�Y!�1��8�h�� ����f�#�eM�f<�,=K�F��N��j��D���s��e�IC�_�\H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���%	v3�t�  ",�ri�y�!�3]o��in�m��+�<4��ˌ�ň��h��j�V��v"�却G�Ct�z&��â&�3ݾw�����$G⃍����,ԯ���gn��Ab�%^�;-оk�	ܷ�4D�Ps��܇�`5��\�vňu�,�s�?�/�2@V�����*�P�1ߒg�A�/�����%>%�����2 � ,w	����[7�d|���XP��� �vBX�y�E�e����KoϬ�ί��#�ڊ<?@��[	J��;I<��fҮ�w�Z�M�_F�k-�!�`�(i3�E����F��j��\w��0]��0�&�ͭ�h�O�0Y%T��BPe.��xu	�>��l%i�-Kp(����2�����VcƮ��.J� ���rqϟ<�^�5��q�\E��0!�`�(i3�E����F��j���0z�cUL�2�c�L��lC��U�T�\ ���A����u�#�$IXe���b���|g�Y�'���Xwd�n]N��F�dH����y���	ܷ�4D�P�r|�֖j��T�\ �͘�f��p�b�z'hۉ)��d�7�qĕ%t̓�@�H�\�{\�"�f'�gܜ�]���>����C����Wj4��⍽аN�By3��<�]�!����M[��Ǣ�K�&�a���i|�l5R�]2�y�Z鎬����x�#w���Ƀ�?PA�c��|[��|g�Y�'���Xwd�n]N�/��A����Q[R�7Kp(����2�����Vc;��2h�����	�rl0�G�ņrŀ!0���!�I%H3�j�V��v�˩��*��c��Et��q���U���V9{)����0��G5���S)��TD��ό���.�^	QW�Q!r�#✲�@���K�*� �7G#+�Ǘ0z�cUL�2�c�L��lC��U�T�\ ��oR��m��%�э�g��L�*������
L'���Xwd�n]N��F�dH����y���	ܷ�4D�P�r|�֖j��T�\ ��oR��m��%�э�ghR�P�����
L'���Xwd�n]N�/��A����Q[R�7��+g^l���v�Z�"B��$I��w��,>����C�x�j؀O���ўC�k�Yl���#�]�!���D��L#���W���ͽ�ʇTf�\kJ���I�?g�f���\X�<����8��UWJ��)�# DY��Wa�b����y�E�nwE��S��}|��XH�����,>$+W��� j/~.)��3\�R�F*}�c}��uO�������R;�{m�B�p)�,)!�G�Ḁ�T"h�p��晬@�1�˓JHn��z��p�Sg�3 ���t��!Z`x-���ˇy�.�`L⯹:������m�5��C�F�=)��A\E#�SX��J|�%eP�� ����Og�r���d��Z�J��|���`�47�q���Z��c��:KYЙMǿI?���V����P�n�lx�k��V�4����,D�H�p0�����}�S�'�d�6�91|�!��3��zl����b!��u�|��sQ�GD��P��Z���+�J���q���U��@����gG��s 1����FE��E����FZ鎬������_�,��T:���V�ÿ�����!�`�(i3�d�٣���N N�S����6�vhW�2�w����g���<%�n`5�fK�\w��0]b!��uፄ\�2��s�pRF�E���_�S�
utY�{'%s�ui�铨g��U-�ez�r�6��g#j�V��v��=�����n`5�fK�\w��0]b!��uፄ\�2��s�5irAz.l���+�J���q���U��@����gGm��s&}o�+��\���Z�n�f��Z鎬������_�,�� ʔ.te`�\1^O�0Ox�%�d�٣���N N�S���g#j�V��v�1�8*#�$�H>+�w�\w��0]b!��uፄ\�2��s���1�, �ޡ.pz�Lۘq���U��@����gG=%� g�Vv�܋�n焞�a�W�Z鎬������_�,�[/�cWM���Xy|�Wn��[��Lp�d�٣���N N�S���c��:KYЙMǿI?B����\��n`5�fK�\w��0]b!��u���_~s�8�c�kg�����+�J���q���U�h}Nw���U�m#j[�E�`JcU!�`�(i3��Q]� _�rs�i��s�٭���lC��U�T�\ ��i3�|)sՀ�T:���V�r>�[I��:!�`�(i3���+�J��Y�{'%s�Ǹ2���;�¬pX��g��U-�e,%�0g���[�=�5x��,����I!�`�(i3зq8�Ј'���Xw���,DU�m#j[�n>���w^Ċ`���Q]� _ό���.�}�
�?�&����(Au.$���!�`�(i37s�9���o>��l%i�-����n9�&+��[N3Y��P4"�,�>E���]�!��	Ǹ�y85��3}�@�7"j���b7|#9���b!��uፇ,��7-K:ٖ�i��!�`�(i3�d�٣���N N�S��+\�g����)e��r>�[I��:�E����FZ鎬������_�,�n�j�<�� �e�d����V�%�1�d6�[aI�q���U��@����gG�F��o�F�M��:�j�%�֒�n`5�fK�\w��0]b!��uፇ,��7-��v
�Mˆ· ���4�d�٣���N N�S���DP֞ �'��L���Υ�d[g�E����FZ鎬�������(���:���U��^"4/���°������R�wX��}�
�?�{U�����?9�׈(!�`�(i37s�9���o��S8�:��Q�Z��"u��������f�՜�T�\ ��i3�|)sՀ�T:���V�9mh��n��V�%�1�d6�[aIY�{'%s�rOw����ZU2h�d�+�q�Q`����"X��[��Q[R�7ݓ��E� ��A�Y�����N�"�,�>E���#�ڊ<?@���,D\X��!��z�>(n��LT��8C��x z�Jm]�#�;� ݓ��E�0]��2�O2/�]]��"�,�>E���#�ڊ<?@���,D}p$_~RSwx�x�K_Dk�����Q]� _�rs�i���Ӧ�am�T�\ ��i3�|)sՀ�=��b�!��&����k�%�֒���+�J���q���U�ԡ/�f�<�i�L<v�<���f0� �ؔe"���3�^"4/���F���ˏ��Z����V9{)�K�&�a�M����*���ic)�̩ƍ2���lĄ\�2��s�(7�QЄ��UJaB)P<�ܓ�YC�4M/�S�@9m����1!�`�(i3�+�)���A�qIp��K��y���=��+g^l��~��w3*)+ZtD��q9+t�}��V9{)=�?��3�����3���b�l��Ƀ�?PA%�G�Q�W�/w1z��ӊo�*H��&�C��|u��%>%��/w1z��ӊ�[�0�7��I����~u��%>%��(@X~�H:��}�S�74/����ch>[G�
 �_FE�:�	^���y ��-O$U1���~!�`�(i3!�`�(i3�#�-�p��q�$x=���P�z�1�rݓ�r���n��뾦��.�g3ZrZ�0m�\�O�W,�P d��s+K�T�=qއ*|8�TO����aF<��[��CC��z>9�R��d���!it�td���5o� c �����v1��k�5l����w����7,������Z�ש���&��[�=�5x�������n�c%ij��d�3F�
����{<�����]I�3Ԩg��U-�e�,���6+���èVuD�*'��>E-�N\��be�����E8�c�r%�t^sRK1сF}���V6�Fc�45'7���ˇ��2���xx��"u����ù]�����b�38ܽ!�`�(i3!�`�(i3!�`�(i3�������l�X%�;���H����_��`:,��� �e�d�����^��U�&�j�G�ZbyBH�}�x�Va�ir�,��7-�B�9��-|�]�[�����k$ !�`�(i3!�`�(i3'����t���}Dq�f��c�r%����:���P"G�wk�>_� �Z���`���`b����d�V��l/�#⃓a���80�iN�
_�Ƞ��ղ]��nF��kJ2������n�'��4e��ޠ���!�`�(i3!�`�(i3!�`�(i3w�HjW��ǟ,����In�h�u׆\���>��S&Q�f���fa����xy�ˉSbT��;�k
��R/�fcXy��q;If�b��_�1����!�`�(i3!�`�(i39�O��F���{S'���.�g3Z�)V��B�1�N�'t�c�I��q�o� c ���r3����MPd�)T}|�qx2�Cm�w���i���Z�ש���&��[�=�5x�������n�c%ij��d���0y�	�B�e�X�}�f�����AӶ�H�Da(􆿳����^�����8-|�D�����y'l/7w|]e:q|+�������{U����ƻ��W\Dܬ��P�|T�|N��+#$|��o\U|~^��zu�D(���B����V_���07��i:���_�1����!�`�(i3!�`�(i3!�`�(i3��%>%�������y�?g�j�P\��be�����E8�c�r%�����!(Ƒ��jVѭ@!�`�(i3!�`�(i3پ[���-[�g�DPp�T�=qއ*|�X�G[����t�T��?E-h���U���e�&�2����{y����i�q,?5q�E�a�8�X�G[��ݚ�Н��r$ɓǉ�.y�U=������&G!�`�(i3{U����ơ_�;+�}�{_8�Y��=�}�Vݨ��}Dq�f��k��^�1��dc�@c�����h��-����!�`�(i3��;��L��-q+�u�M�Һ��;��Cٯu��U`�PW}��[��o}B��!f%��ݚ�Н�?V��j�c������n�|M�U��b�z'hۉ)��MgWĪW)��� ��O(� ���}Dq�f��߆�p�hع��)/^��>&S�XQ�u�j�fKÀ�:����j�V��v�Gj7�uz�Va�irw�+ʝ�lQ�T���������*��ޫ�8�Wp��;�{��!�`�(i3q�\E��0�X�G[�v{��lw	�X�G[��ԝy'�
�:qEp_f���$'l/7w|]�o
�Z����b=�W!�`�(i3q�\E��0�X�G[�E�g�������(ӈ���m�r����
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��φ��<�6�i�:`�+P�� �R�}�	76�&�;��|B�8@0]�¯��^�Hmr�C�4M/�S�@9m����1K�VSƅ��	^���y�<�8ҟ��Ƀ�?PA�b�'�wJ:������������-��{��ڥ����Ⱦ�$�������_j������bg�GM�(R\֎u��w�`L�\܈�X�;� ��;՟��}�S���/d�m��]�e�!�`�(i3!�`�(i3��7I��٪�E�d�똚H
�=�Gs]k�WM��q.��5jDh�Ҭ����j�V��v���"���%�э�=1�5����!�`�(i3!�`�(i3!�`�(i3!�`�(i3uD�*'��>E-�N;
�����I�xѴ����C2�����NۥUn��<�ry^�!�`�(i3!�`�(i3!�`�(i3�q�9�ͭ�Ƀ�?PAC�A�η�=A�qIp��K�ܼ8��v��� �f�?ǉ�=!�`�(i3!�`�(i3!�`�(i3����a��҉�)e��W�3o���)e��,qh��_�G!�`�(i3!�`�(i3!�`�(i3!�`�(i3T#�3�["�",oMG~��Abh��)e�������?�y�Mu�O.C�U��B��-g>C$����i��T^���M�ｂ g���=����tc�.�u�v��� ���`UNP�G�&ց�*�#�vzR5�<���>e`���*1����l��-4fV���d�ވQ�:�G��Hb� h�ҩι�+�t2�4��A妡��M/*�3���X�zK;��t��:!�`�(i3��+g^l��~��w3*)/�k�2�i�:`�+Py�b�G2!�`�(i3T#�3�["���'(��Ь3Ǽ��)P<�ܓ�Y!�`�(i3T#�3�["�7#1=��*�Ь3Ǽ��״$(�>g�!�`�(i3��jVѭ@!�`�(i3��+g^l��+��\���,�����b+}y[!�`�(i3��+g^l��~��w3*)/�k�2�n�)�� �g!�`�(i3H�%�sw��)e������e�r/�1�Va�ir�zO;_�bZ�`� ��f��>�X6�j~�'�:�w�x�j؀O��)����bXe�Ɵ�s��H�RtV�^!�`�(i3�$�������_j���H^�h���i��}Dq�f�!�`�(i3�\�2��s������x~>#�+#��]��}Dq�f�՝� s�#���k$ !�`�(i3�(R\֎u��w�`L����Y� ��q�$x=��!�`�(i3T#�3�["���'(��Cw�Hm��/��kOT!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �m�ڨ�hծ�ݓ�W���Mh��S(����>e`���*1����l��-4fV���d�ވQ�:�G��Hb� h�ҩι�+�t2�4��A妡��M/*�3���X�zK;��t��:!�`�(i3��+g^l��~��w3*)/�k�2�i�:`�+Py�b�G2!�`�(i3T#�3�["���'(��Ь3Ǽ��)P<�ܓ�Y!�`�(i3T#�3�["�7#1=��*�Ь3Ǽ��״$(�>g�!�`�(i3��jVѭ@!�`�(i3��+g^l��~��w3*)/�k�2�n�)�� �g!�`�(i3T#�3�["�7#1=��*�Ь3Ǽ��)P<�ܓ�Y!�`�(i3���g!h!j�V��veK�	�$V�#o�]�ʄ�	]�k��,���^���'ƃ�3�Y۶&��L�H��>E-�N�Ӗ�����#���T�!�`�(i3;�jmT�#��h��G�@�/�Hp����6O!�`�(i3!�`�(i3�$�������_j���QCH�9#G�>������!�`�(i3��jVѭ@!�`�(i3��l�^!Fڸ�>P��=����h�ӸK)~� �ݚ�Н�
�:qEp�;�P�t�5!�`�(i3��F���K�&�a��i
�i�w)P<�ܓ�Y!�`�(i3�̢k���b$��ڣV���^���'ƃ�3�Y*���k� |�;�Ojz�$�AՁ�Va�ir���J�sy�V��R"�+�e�* q��j�J^!�`�(i3�x=��oQ2w���B}0/0`9N15s�FF'l/7w|]�o
�Z�0Qxj���;R{��J:� �e�d�� L#_/�e�܌��!��!�`�(i3(@X~�H:��}�S�k�:6FY̆�a�݌3)�!�`�(i3�_��>νrj�V��vN#~8"�Z�*\�x9?&�8���&�!�`�(i3x�j؀O��(�\G�@�L^�?����NM���!�`�(i3T#�3�["���'(��Ь3Ǽ��)P<�ܓ�Y!�`�(i3��w�w:�!�`�(i3��l�^!Fڸ�>P��=����h�5���`�!�`�(i3�_��>νrj�V��v��=����n��뾦�!�`�(i3HN��R��bP�63Z�t���%>�rG�@�	������6���WW	�Ec�&U�)j�S�_��>νrj�V��v��=����%��v���ݚ�Н���V�?z<�2�w����r%�4¼�k�����&G!�`�(i3(@X~�H:��}�S�k�:6FY̆�,�F��P��}Dq�f��_��>νrj�V��vN#~8"�Z��wH�/�A�qIp��K�=@'ѥ���'T���+�%�э��8�>�}�D9��ɰ���|e"�Ra])n#���r����;�jmT�#b$��ڣV���^���'ƃ�3�Y*���k� |�;�Ojz�$�AՁ�Va�ir���J�sy�V��R"�+�e�* q��j�J^!�`�(i3�x=��oQ2w���B}0/0`9N15s�FF'l/7w|]�o
�Z�0Qxj���;R{��J:� �e�d�� L#_/�e�܌��!��!�`�(i3(@X~�H:��}�S�k�:6FY̆�a�݌3)�!�`�(i3�_��>νrj�V��vN#~8"�Z�*\�x9?&�8���&�!�`�(i3x�j؀O��(�\G�@�L^�?����NM���!�`�(i3��jVѭ@!�`�(i3���̰�!��U`�PW}D��ɍ�ٝ'�j
/��ݚ�Н���'T���+�%�э�X6و�cµ���(A�,"T�z�D�R!�`�(i3��+g^l��+��\���,�����b+}y[!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�t�mJ�0�6���6��Ͳ�h"QU-�\��������l��-4fV���d�ވQ�:�G��Hb� h�ҩι�+�t2�4��A妡��M/*�3���X�zK;��t��:!�`�(i3��+g^l��~��w3*)/�k�2�i�:`�+Py�b�G2!�`�(i3T#�3�["���'(��Ь3Ǽ��)P<�ܓ�Y!�`�(i3T#�3�["�7#1=��*�Ь3Ǽ��״$(�>g�!�`�(i3��jVѭ@!�`�(i3��+g^l��~��w3*)/�k�2�n�)�� �g!�`�(i3���g!h!j�V��veK�	�$V�#o�]�ʄ����n�0R�0�iN�
_�{ݮƻ�@T��6�F���N�DNlvr5�Dѯ���-����!�`�(i3���̰�!��U`�PW}�Y��{�D�~���!�`�(i3^	QW�Q!r�����g��Mt���"��ӌ�r!�`�(i3^	QW�Q!r�\1^O���Mt�꾸b+}y[!�`�(i3�k��^�1�\�2��s���1�, �y�`��vN*���k� ��$J�L�l:�
d������&G!�`�(i3ݑ���&�d��ҟw����f�\%���}��ݚ�Н���'T���+�%�эȈ]Z�����q9+t�}�ݚ�Н���'T���+�%�э��8�>�}��q9+t�}�ݚ�Н��Ra])n#���r����!�`�(i3�$�������_j���=n��c��>������!�`�(i3x�j؀O��%c5#	�.� ����7����|e"!�`�(i3x�j؀O��(�\G�@�LX��ͷ(�-���|e"
�:qEp�;�P�t�5!�`�(i3���F��O��ݚ�Н�t�td���5G�&ց�*�3QAZ
0��3��Y$���F���K�&�a��i
�i�w)P<�ܓ�Y!�`�(i3x�j؀O��(�\G�@�L ����7����|e"�H�����J�g�*�7�~�k�_�mS8<�n�ݚ�Н�ݑ���&�d��ҟw���Z9�+	����3��[<�m��I�!�`�(i3�\�2��s�pRF�E����4�'��'�Ƀ�?PA������B
�:qEp'{w#/ B!�`�(i3�$�������_j�����ur�?lqT7u��2�!�`�(i3��+g^l��~��w3*)/�k�2�n�)�� �g!�`�(i3���F��O��ݚ�Н���O�������ϒ!�`�(i3�%t̓�@���{
Be���C���������ݚ�Н�T#�3�["���'(��Ь3Ǽ��)P<�ܓ�Y!�`�(i3x�j؀O��(�\G�@�L^�?����NM�����'T���+�%�э�X6و�cµd���2��C��C&���mJ�0�6�fĉ>99��|��3�W?�;�끶���A��Vx���_>
xM�v.���e\:"t��Q� �_tt��`���`����=�˨6�o8:4�I���c�90Mj�dL�d�G}%����3f�;�C�f��wFlE� ��xjzӝ���w3��׍�&�U��f�!�`�(i3�c�r%���32��B�dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H����|��sQ�GGE�"RM?��y�!�`�(i3Q� �_tt��`���`v{��lw	�Jw��3�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��jO.�x�����'��L��ʮ�X��:�4��}�<��'��L��[���	�p'�,A��89��A$�P��O�@י����z��q�`���φ��<�6�3�;5 M�|#HK�����qD��=a�^7�1tSjv�?V��j�c<o�;)�y�7u�T�M#dK7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩ�yo���_$���Uŗ�4�=+��-����!�`�(i3�c�r%�{q^:� ,��rQ�f��1.X
�:qEp�;�P�t�5fĉ>99��A0ok�׹�S�C��-<o�;)�y���:W���4��}�<��'��L�������U�k�
�{U�����%ϨEѠ��nF��kJ2�,����Iwl53�e�'{w#/ B!�`�(i3!�`�(i3!�`�(i3EOJ�uxmNۥUn���&UX�{6j�"Hs,�%+���S�$?1fs5��S	JZ�_��=�q���\�rҖ�A$�P��O�@יߌ��omq�:Fa�7�����PϾ���"sS<GYqcHTX�';��#jx��7�֕iK�D�b=k	䶙%T7u��2��k��^�1Aj��t�35L��$
8��2�ֈe1tSjv�(@X~�H:-q+�ۢ	:j���}�S���k�{����Ě����ڻC�i�φ��<�6��(R\֎u����ȫ_V��ˀ�!e�˼S������
�\!6�o8:4�I���c�90Mj�dL�{y����i�q,?5q}�P�|��U���e��d9=���u��r�助+g^l�h����M�E�g�������(ӈ���m�r������$���͜P_�_S:g�RMm�o��'����u��r���_��*��jC��6�g���'����u��r��^	QW�Q!r�#✲�@�e*��@O�/�B���aږ<�#�;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�8���SY�N��&Y��V�Y|�#�)�(�X)��#��Eo�3�IX0F�MV�ҁGG�K�BN
\����8-|�D���"sS<GYqcHTX�';��#j�������%�э��5)��Z^�q9+t�}cp6Dq���e������/��$ʖT�q9+t�}cp6Dq���e������L�$�K�d�q9+t�}ȓM�Me��1���{KB�u.$���k������8���[{/;tiND�S���/9�=eSe.��a��o���H�RtV�^�\�2��s���1�, ��4��'������0��G�|G�N.�N��}Dq�f��,��7-K:ٖ�i��	d���fcXy��q;|X�����N��W��fcXy��q;ko�����2��h��M��:�j��T��hf���3mx��Y�-�_{sxJ�a$�Y ��M�
QC7�T���Ek���,��5ߧE4��Fr��jj,;P�j�x�j؀O��w���B}?�4V�I|�;�Ojz�#�,t��B��?g��>��W�.��A$�P��O�@יߌ��omq��.��|ȃ����qD��=a�^7�1tSjv�T#�3�["���'(���#QSU:��8���[{/;tiND�S���/9�=eSe.��a��o���H�RtV�^�\�2��s�5irAz.l����Z��R��'(�����W���Ě���aT��3G4�����љ%��t�C�G����]'\gWg��	�Z�kfcj��r���(&�L��'ž1�|��P�:k& ��-����^	QW�Q!r�\1^O�Z�_v(��ƍ2���l��Ro�G/]%�z�-uͺ�s�η3G��Hb� h�ҩ�x�j؀O��`�����?�4V�I�\1^O������$f��_Ub���uQL+��φ��<�6�v���Y,���K�&�a���R"`s�]j�V��v~q�z���x�j؀O���}�Ͷ�,*�����<�+��\��]N� ����sp���#��JeW{o\��6�o8:4�I���c�90Mj�dL���èVxjzӝ���w3��׍�&�U��f��_��>νrj�V��v�.R�n�)�� �g�̢k���"��w6�0��ɗ��zi#Y)M���Fe��-����^	QW�Q!r�{F��#�P.`�]3��%�э�X6و�cµW���b�0��5ߧE4��Fr��ja�U�ے
��=m緒x���LU��x}���cB8��I�G�p�PP��#��s�'	�?��[n8�A�A��Xf��&�W��	]�	�U��)���Y;e�iK-pm!9�>������y�:Fa�7��׏�����Xf��&���Aɘ%;�jmT�#�U���e��d9=���u��r��^	QW�Q!r�fN�ї�;m*�z߶�{_8�Y��=�}�Vݨ��}Dq�f��Ro�G/]%�z�-uͺ�s�η3G��Hb� h�ҩ�yo���_$���U���LQ�/81tSjv���'T���+�%�э�g��L�*�v{��lw	9mh��n��V�%�1�D"!���gfĉ>99��A0ok��$f��_Ub��7��G_��$�)�vxK���q
�֥g>i�
�bvxc�V��	��yM����O�LǞg61 ��y3ĝ���l��%�'�M�
�oz˸�%�7�� ��x�壃�5���g!��*ȑs;��|B�Sa���7j�V��v�f0� ���nF���<�W�.�P��'�h�.6j�"HsP����x�S�ӄz4S���2�S�&+��[N��J��ۍb�o��_�Rv�䩲$����E)e|A��`���φ��<�6�3�;5 M�7�癆cgR������������ h�ҩ΅��'�u��'DV���b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-����u?�:�H���z��l t�w�@�������&G�wӨj]h��;o�� ������8�~�;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6����'�u��O��\����'�u�W��is�φ��<�6�@a� ����C�'�ąd�G}%����3f�;�C�f��wFlE� ��'ž1�|��P�:k& ��-����q�\E��0����V_�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^���ըR��Bft>��G��Hb� h�ҩ�EOJ�uxm�7u�T�M#d��+�T[nHN��R��bP�63Z�t�5ߧE4��Fr��jO.�x�������X�ƫD���'$�}��u@:b����d�+4��8�ڙ�^W7�}}��%v�\���ۭXX���X��O���r����!�`�(i3!�`�(i3���'�u�j>��_&�M��)e�������U�k�
�\���>����!�|D�nF��kJ2�,����I�m���Ar)���r����!�`�(i3!�`�(i3��+p��qR��e�����#9xf��g�!�`�(i3!�`�(i3�p}8����%�#�"_����Ӵ����	 �e�d��t`!��K���)e��x��Ca���x�j؀O��w���B}���$�Gv�A���A��Q\�_qd*���φ��<�6�. t��/B�M��:�jq��i7����M��:�jo�YmHA�",oMG~�ǘgl�ف�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�A���A3�p��(�7w��\�Z��N�DNl�S�k�l}
@Ŧ�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3���̰�!w���B}r��x�~�iK�D�b=�E|=#���!�`�(i3!�`�(i3!�`�(i3!�`�(i3�%t̓�@��܋�n焞�*Dѐ�Q�-l�;���P�����=���R���8-|�D_dW����w� �O[s���?8�F���`UNP��Yw���ӥra����!�`�(i3!�`�(i3M�����\���Pi&BL�ѹ�+�t2��iK�D�b=G�6�!~�%��v��!�`�(i3|��sQ�G�չ�Ad��q9+t�}!�`�(i3Gu�b��	�_a��jPG��ݚ�Н���B/�w���B}/�%�� ;̃Va�ir��_~s�8	0X��f*������&G!�`�(i3;�j����E�
 �՛yS�RD���y��lD��{���4bz��26��*��;�ݚ�Н���jVѭ@!�`�(i3|��sQ�G����7E�/��kOTfĉ>99��A0ok��?V��j�cC��6�g���8���$��}Dq�f��W.���f�̰\�!�`�(i3!�`�(i3��LD��C� �\Yy��Z����/����r<�X�!�`�(i3��;��L�ז�1�, ��0in�p����2+m�ᾣ4��L!�`�(i3�K�&�a������kO�q9+t�}"WK�o9z�!�`�(i3y�7a�; !�`�(i3���̰�!�Xy|�WCw�Hm��´M��sȸ�"rR$f��_Ub�F�S�1 �(@X~�H:����dܟz�-��h���`|M���b��i����H���u�(�,�˒�gɀ�X�Z��Zj���
����0��G��e�������5��X���+���b�6��R����VPYu��r���2��}�����U��f���0z8#һ����~���U���O@���zxC5�h3]�< :�՝� s�#���k$ ?V��j�cC��6�g��3��	cA霯}Dq�f���Ě�����}Dq�f���M2ϼI�)�ݳ�1���S�Y��� .�P�2�`W������|C&&v	����B��´�<�p��GeY�?V��j�cC��6�g���8���$��}Dq�f���!J�"�f�̰\�!�`�(i3!�`�(i3��LD��C� �\Yy����S�	RN&c�@N� ��H�����\�2��s��W��7=G��Hb� h�ҩ�?V��j�cC��6�g��'�^�����ݚ�Н���jVѭ@!�`�(i3|��sQ�G��*(H=�ƍ2���l�HN��R��bP�63Z�t��#�a�Ą|�;�Ojz���)e���d��-��!M�2*详p*�з=8k��.ͥ�H�RtV�^q�\E��0�p[nۈ'�^����!�`�(i3ϵ�֚��e���B���&��;H��wFlE� ��;�jmT�#x�j؀O��w���B}�����z��>!XM�#�yP��C��?�T'����M?��y�!�`�(i3���̰�!�Xy|�WCw�Hm��/��kOT
�:qEp'{w#/ B!�`�(i3�K�&�a������kO'�^�����ݚ�Н�$f��_Ub�F�S�1 ���w�w:�!�`�(i3��M2�!m�vINk���������|e"ݑ���&�d�����l9�̪=����b+}y[���%>�rGO�D mWN�2��}�����U!�R�-�_���|e" 0,�{��ϰ/����_�!�`�(i3!�`�(i3�[�H���,�}d��̷mq�a�G�p�k��M�,�˳�*CyP��C��?�T'����M?��y�!�`�(i3���#�cQfcXy��q;�˹�+�[�G���Kg�>x��:�XH�J�#�������J1	�R]�B �ݚ�Н��H�����X%�;���H����_��1tSjv�!�`�(i3~BĿ���N����dܟz�-��h���?D�8��.Y΄�l�j��M2χ����a�)P<�ܓ�Y!�`�(i3?V��j�cC��6�g���8���$��}Dq�f��\�*:.����k$ !�`�(i3�(R\֎u�=7�7K�P�"ª�����}Dq�f�!�`�(i3|��sQ�G���I:)�/��kOT!�`�(i3�c5ew�|�;�Ojz���)e���d��-��!M�2*详p*�з=V�Q�� h�ҩ�!�`�(i3EOJ�uxm�}�Z��yn��뾦�!�`�(i3՝� s�#���k$ !�`�(i3EOJ�uxm�}�Z��y%��v��!�`�(i3���%>�rGO�D mWN!�`�(i3��Ě�����}Dq�f��mJ�0�6�!�`�(i3��|YOF@ܗ�6���L�~�[_.H Pu>�<~K!�`�(i3�%t̓�@��܋�n焞 ����7����|e"�wӨj]h���z��l 2�����4ƍ2���l�!�`�(i3ns0mWw���B}/�%�� ;̃Va�ir��_~s�8	0X��f*�x{^4��*m!�`�(i3�2��}�����U��f���0z���|e"
�:qEp'{w#/ B!�`�(i3��M2χ����a�)P<�ܓ�Y!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok���wӨj]h���z��l .+�N�R����|e"��w�w:�!�`�(i3�%t̓�@��܋�n焞X��ͷ(�-���|e"�H�����,��7-u��Y�rG��Hb�H��
J��!�`�(i3|��sQ�G���I:)�/��kOT
�:qEp'{w#/ B;�jmT�#�(R\֎u�,��7-� �9�!�Q��s�s�{��ҽ��d9=���u��r��!�`�(i3|��sQ�G���I:)򊎆NM���
�:qEp'{w#/ B!�`�(i3|��sQ�G���I:)�/��kOT
�:qEp�;�P�t�5!�`�(i3���F��O��ݚ�Н�EOJ�uxm��M����%��v��!�`�(i3��M2χ����a�)P<�ܓ�Y
�:qEp�;�P�t�5ʁ���Mյ$��Q��@&U�)j�S���̰�!�Xy|�WCw�Hm��/��kOT?V��j�cC��6�g������;q��b+}y[�2��}�����U��!]o���)P<�ܓ�Y�wӨj]h���z��l (�?qE��w%��v��HN��R���
�Ŏ����ܐ�}�JX ����D��
@�F_���k����1�����瑨R����Fҫ�5Ymg�CT�\U�d�#�bp�z�E��':5,:b
m;�E,	P�QUH6"�w��B�j���;�����cl���,��7-�B�9��-4�@	�u�a��4	_��%�э��XW�G�<v"��1^�!�`�(i3!�`�(i3?Q�@X>#�D�ʵ�b�����"��Ϙ;�b��t�|K�mb�˿�Mq��M�!'B�}<��}�t����*��1�&p��)e�����FV\���;z#�����UyP��C��?�T'���� ��F2�!�`�(i3��7I����bȱ>�Ѥ+�Ä��#��Eo�3�IX0F�MV�ҁGG�K�BN
\����8-|�D���"sS<GYqcHTX�';��#j�@��v{�G��4AL���c����L�{�q9+t�}����@|��璓�c�������t �[l;M?��y�;�jmT�#b$��ڣV>&S�XQ�u�j�fKÀ�:����j�V��vi$'�vu���эp��6+q><�ah��e��������*��ot5^ݿ牴)e�����FV��:����j�V��v�/�/�r&l������y����jSAB<�L�V_�I����~u�X%�;���|�W�믜�}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ��RL� `����f�nd羬U	�`�o��_�Rv�䩲$����E)e|A�յ[+8��r$ɓǉ�.y�U=������&Gݑ���&�d�����l���}ϴ�%��v�ڵ��R��Q�-l�;�zigzA=v)�q9+t�}����@|��璓�c�������t �[l;M?��y���l�^!ЙMǿI?��t?�@����}o��Xy|�W����W���#�a�Ą�iK�D�b=`u0�F��a�Va�irmyC�0kc��g���Qrf�R�}S��,��z��l ��΂����-�������R��Q�-l�;����p
v��}Dq�f�����Mp�ЙMǿI?��g�F��6&�U��f�!�`�(i3��_~s�8�c�1���7�`|M���b!�`�(i3沙���A�0q�#术}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍн�Js�������lIR!	=�^/���'�i��y��숕iK�D�b=��L4��Մ����XF������lP�y��WZ��iK�D�b=l�rx��E���ŕpO" �e�d��Q"���_�p�@OM.Ir��yb�	�����u��
�b~*��s�!*Ĭ�����|�x@�iK�D�b=`u0�F��aȗ۰�=!�`�(i3!�`�(i3�F���ᘮz��l t�w�@�Ԁ����2|Q�-l�;��5��t�;��Cٯu�Xy|�W�����z��s)l໶�,!�`�(i3!�`�(i3[:���[}�p[nۈ�d��-��!M�2*详p*�з=I�^$D����(R\֎u�{��b�b�*���";Yy\'{w#/ B!�`�(i3!�`�(i3�H&&��+�O�XÁÿ�����#o�]�ʄǃ1a�Hj���Z���m�����a�,��7-�B�9��-Ho{�0!�`�(i3!�`�(i3!�`�(i33��0��|��sQ�GGE�"R�V(MH��C��|���j�֎��](g���������l4N�J�ףǅ)�'�N7�����\fcXy��q;_��y���ݚ�Н�!�`�(i3!�`�(i3!�`�(i3�$�������_j���W�TU�-��`�2!�`�(i3!�`�(i3����a��҉�)e������WՇ,��7-��v
�M��⍇���!+�+$�����z��l Ю��U������2|Q�-l�;�Kͽ<\��;��Cٯu�Xy|�W0/0`9N1s)l໶�,!�`�(i3!�`�(i3kǿ�E�Q�C��6�g���7t��'����+���b�6��R#o�]�ʄ�;4�zu%��0q�#�<���H�
nЯ�O�!�`�(i3!�`�(i3���>���Bft>��#o�]�ʄ�< �SS@�
�رjwc�gVdxQ,�K�&�a�/�dI{�W��j�[O��!޽�d�E;4�zu%��0q�#��?�iZ"x,!�`�(i3!�`�(i3����(��e
� <"w���U���LQ�/8��u��m�byBH�}�xf���fa��myC�0kc���Ø��4��Va�ir��_~s�8� ���3�<<��lpЙMǿI?��g�F��6�5掼�s��ݚ�Н�!�`�(i3!�`�(i3�,��7-�K��*\*����d'��",oMG~��i�*O���2�H����ϕ��r�^|�;�Ojz�$�AՁ�Va�ir�\�2��s��W��7=#o�]�ʄ���wK�;� �e�d��}��NY��}vރ�d�,����I�<d��{�v. t��/B�M��:�j��/���+��u��m�byBH�}�x�6�[��y_�e�������{
BfxQ�-V�N|~�.�u���r����!�`�(i3!�`�(i3~���e��?5��wnj���)e��e���N�Sc?0G.{T�2��8��Ս��%�r� �7���U�� �e�d�������km�������.����px��=Uy�,�$ک��&����k �Ģ��|���jVѭ@!�`�(i3!�`�(i3��'T���+�%�э��5)��Z^׆p�9��+:��0	��