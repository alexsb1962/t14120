��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~�/�gXŨB�>KK�z?�������=�O�+8&6�ͿN��}�����nE4!}Bj�Ɍ���+|cˤ��f )���V3��3BY��֟���FG�jA���0�0��[pJۡ{��V2�����֪��:} ��:I
���p������C���n��CG�o�8e�f�.(܌���q�����Q�S��֟�]Ž(��M��Q�C$�"+�0dN�D�L@?�`za�Tn��Q8.�fJ�D��L�䞸�yvSH�H0K!���"���;f���"~���{�^��V���������3q�e�@���J�rHgv)�� Dl��-��JB���U��&�H�r���N��?�BO�pǖ�-��"�c��.(�PA&�"��00CV b�gj�G��w�y�=�b��p2=[��Q�b�\�I�5���P%���P�����G��b@|��.uF��������i�S���G�y_�wVu龛��<�u�5�����Ɏ��YZ�+������/��o>!�E�Q.�$�����p�;m��CTJ����s�&*�A��RB��CpAH�f�/v�\���H}����F�&�pE�r���k0�l'��6�a��
�,� ��A��R�����'0Xz�C�A���MO���}��ہV�Ƥ?�~�F��w�~淿�q�.!��Z��ۑG��^���=��܁�L�M���<My�9�qT�Qo�6Ȣh}�h2��<P^��lGo����w��	H�Z��+^>���C��q�L1��?աJ;u�k�~H��6[�c鼭�е�w�?�S�8��
��Y�0��z(����|���R3=�8�k����gK���jJ�[NUEr�-�I-o��M�8[��$�R��q�ne©���Ζ����3��C9$�������wR���)��sbI���\#B���ѶJ:���UH��Ca�t0*~k�#=�T��Unr����R��Y��0I|+�Nע�⥰F�6�-��m�K��31Nc�R�W]��)��qͥ9M� eu��DyO�t�� �v�o5pa�n������ކu3W��ǊKr"���8�
�nf�_�t������?�n0�#5�nv_Qf�{`b���W�TwZaɖb=�[��QJ,�L��d�wS�/�ޫiB���J�,�=���a�"E�LR�*�>�9�&��	� �bMh��f���"��ɂ�>�� ��i$�Ф� W/d@f����}�Gul�Jt(����v�4ҙw�0v߰�P��n6Գ\�B��[�r �L����
���&����m�B���dRej��)*��H�ґ�=Fplu�1��'4���u[x��4�h�p���(ƥ�m{�3w��>�1Ld�[=����t��XmϭuL>�����n!�d��hG�;����F�P<��y����.b�4�q0>�u��_�����a��9�Wʼ���΃\���ҏ�܀5콍"y�k֨ʨ�RI��|��*�CL4�\'��9�C�d�لGI�.m+���p��!��汧n�_���3�&�3�M4�a3b@z���_\N9�<��T�}���x �X�u�{G;��j�C���MZ�l�q�=�,�((�;�A�'aD�����:�-��T 4��J�&I&�� ������x*���ͤ�^�;o�o��b�]af>�<�(a1Iȵ~֍B�9W�L]���cb�.��`�+>W���%�J�0�ڙLm�gN�EO�����d�@�42�9��7S�7��ڧSZ�]n�.A�����v���\��=��=Nhcq_=��a��[E��2"M���]#�ȝ?��VO�{�̟����PQ��vD�ӊ@�����(���a��8,�Cu�~�h?���ە����T� �`l��
���ۊ���I�I�"�¡��6��2ԯ�4�`��3��4X:4U�Ti�#r���]*�Y��?�O傿B��A0�с��:���u�O����a��d��}9��I�ګ�{�1̢T.����@���8|�GT_��˃	ɱ�+�����i������B	C?��|��Y�0�j%%0����p��R���%A��xs$~}SnC��_�R���;�Ax�&�B��I�#�:g��zc)RX�V�̈��6�`@��1�-��Ľy�K�4��5���Y�T��ki�s��_??iD�N�;�|�И[�1�0��~V��r���sW)m��'��q��_�2W ���BZN�&t*n���(��L�K[7@"�5��kS*��)�Lyz2ۗ\Md���M�(u:2���?#iҮuː�����<���h�u�r/�d�(�4C�QD@�(@�@�3f�s�9CWВ��X�;jaj�v������W.2�Ħ/�N��h���I0����aEW���4�96��x!�ʅB}ʎf�Q�)�go�M���dӹ��_#�
־lJ��z�759,�_&�v̦��F����Eh�
��`Ŀ�!(*?.�{����G�&���`�+/���WH!]+.J�� �~�?�K����S�kgދ6�5�&�}T�an��[ީ˿gT�,��5v���}{u� h��?��*<x藷p��o#���X���b�?ej�}��?�B7%[s������x�g'�ɟN�ˌD�b�,����+�\kx:��P:�:8%�n�'.��D����˔�k���D�%�5�4 }�z����0��^����j�c��C������w��X4uW�h,-�E*�/�/o�'	�� �'����^���S�òEo�c�V?�L\\���c!��7k��(K�xx�����Z0�Y�\���Q
�v�D) ]=�I�2�\���p�h�-�'�A�M�i:������BG�m�~�rk7֝ ��Q�i��������7���o�X�!�{6��� bf�?�&����6t�fhB�HO2.zLTg�=`��!wƊ�',cV�Y�o�0�w���y#�ɓ�����I��L�|�c����|����IgG�H��Yfu��i
��^4t����cc�H/삄�˜�����/�m�!�	���dg��2��ז3��YΩH�B|�s�[Zx�
�):r��fa7z�F��[��R�΍������njC5��a|I
�Q^2�A��k!W|˽V�`z���f��r�j�g?nY�_��+�>D ��z��ϛ#�Qy5��5|�w�N�����H���eV,+.L�Kz��M��)⬆��ʃ=֍���=~Un���M�s�Q��c*��h���\�����1���[�b¤嶽���mg�	��k^�^#��t 2	*��'\��oK�����6���\�P吮ѳ>��ͺ�K;���y��n��쑨N�Xϻ�a��3�ؽ�k�NU|�r����
j��v��lMa�Uc�g����0��A��x:����kMD�?����B��NV�� R��:$ߐ�j�����ۮ��5���)����g�q�|����@�������?s����v'p3�'>��J�F��@�����9�ū�i������E�;<U��.qп6������[��1��ID��uE#��Kd�F��>ᅌLωZL��*i�Fd��^�ؐa*��e	��e�����
�V��=�C������(Z.Z��
2 >��-�g�ԍ�� +�6(ٍa�����Ss��`�z��GǴu��򢝡�o��Z��������C�;�Sl"��|fz�Ʉ��� [vj�S=�K����r�V_���م��]-clWP�l�����\JuO ��AA���I�39u�ܗj ��鲧W�G)��M$}��goj9�dn�T����AS��ؓ���Κ��}u��-ۼ\�����0��Z��W�E��868î����p�
\_�|ʔ����<����cƿ���1�%��#y� O�H�$���sEm� 6�TIuroN��H����&��.��Q8���#jv�6=��j�7�|D��ʀ�y�1i4�띥kF�EޕAB���q�n��j 6o�d�w�ڒ[_� �T7d	E>��u	��5�/�p��nH�
�
Y����O־H��s�Bfv��|% ��Ÿ�`�.z�HUc\��6�6����zK��z�Wc��@�1�����H|�*F
���F>Qg�='��xB�/��U=��<˧�׋�����P�\�����QB����sf�3c�p7D�h\~V\�Xם�67��DcL�q��J-LV�X܀rZ��,+������i�aڛ4�1���S
:(���?�ڡ��
J&��t�}0B���Ï��|����4��C�N�n%��5�L��S�4ˀ�ˆv5]�\��&
�𮖤�d�l!#��xEUs��n����<�C��ĉ ����&=������R��P@n��w%�b�4C�����=��׻y��<�M5�zO�C5�>�lj���
H&��c}�,9;����a�^�
�\ EH���0��
�{>��=1�ߑ>�궒ps�A�KtPd����G ���&]�<�NGT��%�����Ӓ��� U?�К�s���]����'XW���y���_���J=Zk�x��1�5{��,�A�A���l�8���j0�����K�R8*��jlس�W�j�L/u�3G_����3��ɼ�F+���m���/�x�]�d��z��s�c��==��B[��^�a(��LN�I�Yp�4֤B�\�m�w�x� y��~�8��r�]E ����>	Q��/ń��$�QM4a��Zf}����
���o�c�g��.��W�d��Vd@�ff�n��/���.h��_����d!�/HL8�Bx^�w1�1|�������T'Z�z's������b+;��6踋aua$��n�vhw�m�Ʋl&�0�zF��a����B�DG�o���]���g$�0'�	;)_0嗵�����wD�E�N�SQN��u�[َ%��n.���R{�
�}�z٨f�9��c���t�2������^��Tm!o�ka����"<.�P����Ȥ�����p.@;#�VP��-�g������qڐ}{����[!��|q�B=���>����r�#I���%�Ry�����������^������
�X���}�EU��e�*$�����w�0<]+_�LL��n�ru}JBGG�+ �*�t;6�*#bW�J�u��i�7X�a��%6K0v�^:P暒sq8����Ub@k��Q�!�J�3����_�2ͯ���
h��oǞ��CJ�m-rx@kѸ�V��Nˣ`�ȣs��o��k��2�9����7��f��	#�1J`B ����I�� �P�N��U����_��nW��b=���c*~C=qR}�Xz���(΁��m�+�'�ƭ�7��Ճ? �-|<�\_�[�Q�kuɜ�� ��^�2�8[�3{�n7�/4�C|>u�E�Xӹ���`����N��I�a����-R�R�-�(���{��t��6gͬԝ���Ҋ�4���!)�`����>�Ε#�;
�)�����oۻIK$�^����)��H`�8ҧ���$�k᷽LI�-@)�[T`��k m1�I{����d�3\�ۜ�Xu��տQyug�e H�N�O0 L�\�T�Qqvv:���>qu㞤V!�2���p�1d2�Mt��(�G冴�����폼�YE�EQe7�����_�4���P�S��@s'U2�_I�BU�͖����$RC �K�����`ھ��,NS�#9
%!�6[qH�5��v?��<
����K8{8����\�%�#�ݗ&�~lt��-c�AK���� �o}�l.�D��t�n���mќ B��Xw��W��S�t8�|3l,�ZЙ	�x�{��H���*��[w]��CMᎮl�O[2�*}�#x�R&����z �N���QU�$�kũV���)ѭ�qp��F��0��.�dG���
f�1���>ڨ�x�W� U��o%?�����z��=5TDZۧ�q�A�]�W��)ŏ�_8�d\/��,��O�G"z��$�����|��L ��*�5 ��ZjB�#)G�*��#E����}ڌ��L�S�1D���jd�Tb��͝�~���\�Ӻֻg^�3�z����A�k����������ɢH7|�\KW�y�+w���B5ZZ���� ���64 ~	�.L֫���vMޤ�>b!1�^+kH6��5�f�V31#�8@�'P���V��M�t�M�)	rp�+���${�}�EP)UX�����1&H�ނ�)\8ێ��Caݓ��G�;:b�><�7�t4#��O�R�~H�K��U�߿��(� �S��&�V�{O���Ôs�$4��%�vON��Axsz����O�`�d-�u`ˠo��)��@i����z��b�7��٩�&�s��mn��F����ZQ�&g�Lz�Î��� �[h�@i��1��N+� Mex���ɱ �R0O��tJJ	z�fa���P��s�� ��<���w���S� �������ToW��.�O�8�[�hN��Ǘ+v	j�O:��v����K��N�&-�6p����YBg���ib���z���o'ƺa�p�x�[��c�/	�0���abV��^I���\ɂ�(�o盰�[%a��!h�8���R�U���0J�Di��X�x#.��A��e��nł*[��oZ�<ʀI�O4���f<y0������F��մ�ھ���%�x�eka��uaE�C�Au�Z	?:�g���2���[�cX@�=W��ԭ!KF�Gg���
�qt@؊O%�j݋L�c��7�r��Fz�)�e#�Hk�7 �Az�W@a։Pƺ��3�&&A�F��su�I���%��q�"d��,M9׶ͨ^if`z,P����z�	�a��5@M�X�.��������%�9Gl�������ɲN���,������&��x��n����@.�T�1	ȹ,�L)�m��;���P��[�y{�Q%Rh"�S@)��C�"#�������b���3NA���u\��Ѓ��^��e���f�1]U���_�j��7�@"E]�� S�A���D�����T�F[��zF����
�V��pW,�����1�|�;��ZNq�������(2�"�D��Yɝ1�ѵ�M�?U�n���VR��:��������E	{t�.��wD�����,bz�[ңm��u�tZ-�%Hp����]@u��1H-����u��tw�5Q2�B��|�xcqí *�'A��N�:���dw�r��'٦#�6�H,���P�A�ط0ҏX���u�x	��T��l_��9LDq��oH�o���o��cc���uN�^�J|������ŀw+�+gl��Xe��%x'h�&���n,�1B�bN^��3���Blnk&v���A'��
E��v@tLk>%tͰt`�hE
Gp�e:Ǟ�F�&�����N���$��15�<{��~�B��
� ��ė����nɈ��;������p��wMU,:R�A�����ر8~F���c6��Z����PO|n�T��\_�6l䰭K��O�۽z��K�*qq�?�I��U��pZk�]���j�(�ԙ��cc�tYXAF�&���>w�T	g�~����(�L��R飼�1«WÓ�xBh�f�r������	����y�U��W/�KD�����{
5��r��i{��P):��yJ��6|k@�������z"��3y[���Pe�=;v��]=O�V�\e_Q�NY{+��
z:(_'��h��W[6�T��HK6z��V�G�5�T~�5��$S���/K뇀Ҫ�������zR��#Е��E<��@l�&�0@���fŗ�>��ݗN24k��iϷ�i��������~�k����B�I ����0o�c��N��D6om��Q�^��ӗ������*U;5Ѻ�,~8���|T
~�� gs���>��jѯ��i���A��Ĺ[��\(�]|���蘻�tN�z����f��ܗa����W1oU���_:�@�ϸ$��T�-7!������I���=���#�G�R�T�Al��R�Lz��i�=�X+o���ʞz-gk:�X�!9�f���p�.�❼ �tb\�ە��/�m������P`@J��i-�ӛx}ꝧ��8��Fa�!v���,sb5��/��\?�C�$�F�Ѳ�+��pz4Y�>s��P�cFR�ݚo�|ŉgǑ?��p�?TNTݩb�	6���j��A��k$ ����}5��gm�9�
eK �tTa�p����R{J��'-�Y��0D��t	���m�F[~v���[_�����C�y��k��4U�[O�ǣ��.W�5�>7�ݙ����W����ߎ�H�畴6[�+~6�\�?v�9�����3r�r�f�B�瑿�Ц�}�0?W���C$�N���=�?9_�~�/UVw�-x�=�Ο�%s��ڭ�@`���������?���b2�Ԙ�+ J<GOG�T�f�n �/��`�$�6�[��Y��6�.�s�²�ޡ�.�F���ŀE'6[���[4l�CX���� ��v�՛�T����e�B�_��?��N��	1�|J0�UN�Lx���b���8��W!�gYzal]�x~����wBZ�9oo�������@=9>��:�^]q7SW����2�#��6��>��Ol���F�@��/�z)*��ý����&�zV�V��K�!���w8���$����]^�'���d�6.��Hb�{^����UH�]q#ځa�]_�uJ;D�{��D�MM2�.b���(��tU�Ca',�i��HR�v?]5�@U��q�O�Kw�1�vIv�C�����<�,��T;�,ʁ{°��������&�Zck���'"�ɪ��h䍴� �GMHR���x���#|�y%��NU`
J��7��5�o���+T)�VV����2���o���!/�fJ��	:"Āgt��"P�dior9��_z����էG\�����M��ߞ�z�R/���s�+���.�x��?D��"ش)��U��f�̋�/�_ߤR̟�(� ������,��������]7!��x���p�I���~���]4���N���=j��rB0;�}���I�W��C幽j��3E�e!|R�v��2�Nw;�M�lӉS6M�S|� �qa��YdZ*�[|�'���!���������w��8Τ��F���k$�I����!�[�åu��A޸g��Q�zн�g���wBx�	6�)� ���b�����v̛:ܚ�|��݂�H/KDW�����^�J�Q�i��?5W�H
���d)fv<{u�_q�0��9�=�fg�T��C�1|��_��������v�cnIt��W�;��`��<������+u~NS%>���<S�b� �k��P	�ɟ0����Ni]����'�������3�}3����;�e�Il���%�E�`���	�/ި}��3\UǛ�.2��F��E�a_c�G���Xo;�;��ԃ�	d m������*˫ȞjDj�ġ�vP,�/�G3d`�;I
���JA�����l�D����vD9rL+��mr7��A'=�	�i�EH�c��$��¬�"� F�u�LJ�|�LEh�;����N5��\ցg�P*�\A��<D����>���`�L���9>��k �m4��}�y�Ғ/�॒�ڈ�
�B��6:D��n����XlÆD��FϲS)�c��ZA�4LŹb���v�Y%A��1"��f,�H��ϐ2t{���';��a&��&���SVt���O��,�KMx���E���z�r����sXQ?�đ�vr�,R�ߞ�>6}.�+Xbk���_EV��:��`����ڳO�~-�)Ꮥ-z[]R�d�8u>s��'����^�h¤�"���'���Ǝ"Ģ�d3�;-��>�9R��az�����3cl�%"e1�7=�"r�<>|�D��Ţ���J:_4�v�ٷ8!�9�mm���ܝ�(�����O�6۠�g�$��d|4_� �0����ܴ8iVYE�;'Oej�(��{�-Yf,�˨H�j�o�eUX�.h�."�|�.mLR�wk: �TL75�������:�Z����**�T"�5Ǣ�RqM�%���G;��("�i�F�_�~����_��no��������	ǤU�O�i0f�^g��XGF��w6O�qQ�SI�� ��A;{�K�H��R kt��^����&�bvD7��=4�K�7��((�+��@Xs��xZ��mMg3��/���;�s��[���W�<���v^�R�Q�(��"�|����$u�Z�:ڔ)wIr����¨��k�
{=�i�V��}��P/���u�EW��{}��=P��x�V��gl��S(;��fA�O��eWc�iy�ll���fE*���d~����� Ǵ��C_;|djΊͮa�1�	K?�q������K*�7@�$�;��*���/���{�՘�~cr�R�!���E�����J�k�{�Uo��9%u3��\ҷ��"���[Z�f�}-����%�g���v՛P�m�) )r�l���~����bbdQ��o�im�^���ӏoM���s,ve�Djd���]\��k �s�L؝ �0�H:sY��㟔a9T��?��eau��`@o�">�� ׅ�&l��#�-�;G���%&Ҧ2r��t�V�\<kc��֍ǃuj�\yo��Us}��p�RK��J���Xt���-�)i���{�P~[(d�:�a��_���t�E���eۛ,�.N�2;�ꑻ���(�ؓ�� %�2�|����Q���e���G�0���If-�:���]��K�}��{.�PbWAͩV=�0+_���1�xY�K��<��l��B�<t�!�I?��lmD�j]׊�9�B~R���@���)opH��6q�bЦ�����3�5�L��#JKG)��M�[�S�53M+��η�����}D��'C��rS0-�>OW�^?8f��z�$�*�3��t�u�؇��%>��܋�� �u�n��98����m��_�Ƈ�޾X֕�DRP�%�������~��r���z��E��\:HJU��o�oJdKrg�\Ԉ����=;8?�{X�Q �C�>	��:��xC�j��0�4�CtfU��]��\�59СHЂ��N�G���9��h�q�E�*'f	������l�%$�@w��-���yL,N�����]^dnQ6X�xy�ƿ+���<���_.n
$�?j I�Սc1CJR7+�b��4���p�*�+�3�?���9Qd��,�"Ҵ�n�ff��?��W{\MDo�7���kk��{��G�{o���:�R_�9�{#n��Vfk�(x5<�D��f*1Yh��ݫ�Y��xp[J�6��4�9����o&�v9@���ٿ��}�-���2nY'�g�)�&�l'��_�D��S괵񏺇�6�{���L���|��-;�o��e��:_�a�)�d;�*^���� �������,����R��^(ǈ�:�}}5'�jq)l�Ԛ��?�褦�5�'.	�E�[��� �_��D4E���=�ЛC&d�_����֢]:�3i�.1�ݪU��yD���_9l�P��(����b���8��Cl�����<y��&GHc��#Ef,���өϗSI��`���J��^�`���Zt�I��{J4��%��pa��yf��A��x�դ��C��pD�\w٣mw�[n��^X�	-�6FB����Y�Ղ��p� �^��QX~$�Z�~��?�bM"R;6��$�Pl��u�,�Es��Dy�g^ОX��^�`���qO�N��"��j����hC���[�T0h�퐇���%��g�(���^�	=�s��,\�zkp�����0�<�������9��r��!Y��QٿoGJ�jF^Ɵ/�dQi�g8�c���d˛Ue�� H����c�;E!�%^�v)�U��e�D��-��z�Az)�p�-!�����x�U���wEBS[Y/_Ł,�� �%�������l��m9��Qv:�F"Y�}ʕT2��T 2�{:�>�|��{��B��R�>���̊�⺵B0�v!��'g�r�xi.ILj�m�͸r+��/��q�㔐�+`d@eh��(�t8Wh����`��co��pjLC*�ʲ��q�A2ĎL4Z��%Tq	,tQ]��:7�J"��JGj�2��~�<���,�$8b�:'�3;b���_����FT�u��<t�����!�A ���qS��n: `=qF�=6�*�aޱ|�}��0�Dt3I��$/;�2�0���M�z���]�Y���F�����~3����jC:W����<~�M	˃A�ˈ7ZT,U�Pe�z����&)��lF��o	��x�����ƏD�l���8 74@!������V9�$X�9�P�dY!eF�©#��7)7(���	�9�e�͹+��F�9�c��ϒ���+��ֽ�J����'��;@����"_5ȼǵ삶)���b�1|�Lc�܅k�ܱ�g�]���g}���H`��Dם�'Q[���6[~�
xɈ�;n-l~�1��D��q/J�f���-���ٲ�k�gk_ѐ\����v~����f��pLW3�� ����YOۓGw�}��ݏ|�#e��UN+�������e�xN��dՄ舋��\������|0@r=��Ke"%�) �[��>n��v}��4����ṅ��:.�wFI���)@_�����j�f�@�e��(q�z��b�ƫ�$Wf��0���(�!�كI;f��9!��=�g�. ㊅�05�eg;E�T��:0�F�$��L1��vs��:��aR�t!���b�����i�殅���D��ݕ�`֕ZC�~���L��I-���I\1#��k��If�F�HC���i҈�=���W�O�wo�1�3|��� �MMT�c^fY�����i��\Ʉ.|(#҃X#C�z)`ف����,��iEv���<(r
���2D�A������c 6(�=�]ǋ欔�X�2w��TZc��H�k�b9@���g�ֽ���1g��x���\ FGmm�-��vm$����z.)OH���6p�������7Ͷ��t���P�
�w+ }{%S��)8�s����;��s��J�K߼]��	g���c�X�'q��Kk��t��!����䅑�$��{��O���*��y?A֦��*�"^���Q��|��f��`6��O�����6'G�5��")*�PL��b|<h���m[#C&hu�$�42���
7�F�eX;G��"#
�)#ވ^�C�i*�:U�@~i'#�]���yf�Ku��h{��6�gsfCY��"N�v�E/P͇�)@.g�R�Y#�Q���ŵ��C�z��,�5F}4B1mA�i�����>:��~/�Cϩ���oۭ���qˬ����j��D^�lJUS�<oKU��t�{[l�ƲȺ�b:�|����89��-ga|�߲tkoP�]"W����~�5Ϛ�Q�Nd��몓ge{*��:��	���N�BVW\HW.���Z�ѵ4]&�2Bu��D�Ϗٙ��g�f�CY$OIL����yr>B~@�3}7���~���TذO%6m�I�7��ŷ�*�!��)���E�$���0�,J��T&H��/f���i22�g�7�a��q����^��J"�ɓ�
�2}�K��"�g瘕�T@�V���v��4j��;�>5�٩���*c�H-��2�3]Z�X�N�gز ��D�ԧ��K
m�I�}�=���4�wݓ��&�.:�t���8C)�(�������<��Z�� Mg�uP�v��%[�Lդu~�X�����ĠߒvA����e*�O���.?�X_v2�E4Y�.H�N��#ܫ��m�縋Z`�7�JT7��j�!�ܖ7.v^���F�%�x,|��#��,�ٛ���ͪ��6�Ѭ<�R}*��,���'��n�������������!`͏��{*q��T�]r�붇�]hӀ����bZZ1��nV!b�EH�O�<��+oh�[���h-���z���a��#b��)F{T-� ���@��Y�6"��I����2f4�ty%��m���jX�j�C�ljYxG��iۏ��łlI���1U&�q�o"����q��L!N�:b�|�U��<�AIU���ŭ��ˬd�r�.��f<�$��1���S�
s�`]�bs���o$�J��\�l}�6|y����&J��$g� (S������ph����}C��/��w~�s~}P�뿂�[��ۜqi�Α��zʣ�47�y��HY�Z�;T.��z��Mw����3�j��
��U�d�mS�nN��x�R0D>=�=�K�&45��Mj���AY�6�G������Ĵ�R�#U�tz>��0@*L�a�48�iY������rʏ��⤜�}��Qx	oݛ`�v�4l�!l�f�r�n.�����5ɿ�[���V _2Lp�opn�9��� �s��#���[��b�������.�47"������A?�ǆYs	�Z�[;R� �e��v%�WI�[Wa(x1�ݒ��ߍ��dU~�Ȉ��>���	��
�3Nl�m<@#�/�:�<1��T�?`E ��.L��[�=��f'
Ju�"�1�%�H�8M`�O��3��;|�SDϥ���7��C��m�s��Gs�}��!�˵&�Lf�a3�&����B��٧7�gHo�����>��<BjFTG����9�[�*�<v����
e!}`�= ���6�k ���ʣ��9��&@��X�}���3ζ@�9\\`[�X��H����d�C����+tUF�ɢ/�_�	k�<��כ�o� ����*��f�څXˎIֲQ��qf.#���ޣ�m�Xm��\'x@و�\qwL�ן�}n���Rﯮ�5��G.�����V��T�jc�TB<�E{K�� ����8��V�I�wh��W��&�s�~��V?t���R_Λ�E!H�-
��=�`��R�N*���賬-�������:�9����Uy�j#��� �'>"|���
>����j��e5N;�ol�j�%X�,N>�闞"��X誊����ֺ^�3�ʏ8�f�s~/�}�r�#PS��t�c����M!��Fg��ݱ+���1zS������u�f���xW�wЧ{����߾A����0��Td{_�߱'QEՠF�>�׌n��;V���ݍM�X{�*}�a��iS�Rؽ��+å�d��&�3q��'5+BHN�fOs��'~��X��M�5Xn��M�� ����ֹ���N�8�G>�vh�d�8)��k�Օ�sG�g�{G��[N��>�G�Q�%��Wm���:%ڥ'�އִ�w�WT>k*7�����|����%ė��|�rz�p�����>O� ?�FKu�N��-�p{��9��<���CN%�q�g��_\��];��u���KВ,��G{5�	\�c�9!�µg�U����}Z[H���k�]	׻=�w�	��ۅD��`*oM_8�2�KJXs�lu���H� ���,V�B��q�t����'k����es�=��#��b�LÈ���85Iы	�A>�n�O뾀_G6�^R!�t�bC�d׭`F���3qd��TŨ�7>�)�^�A׌I�^>��M�}Eb�.�ׯ�'�S��K��E�Ɉ��my��[j�����+����8�[
�N���*���o��w��'�b����1Ŭ�2�}Z%2~q�?j�\z5�P����C�6��#�*\�R�Uh�C���M|�8~W7K�S��B���) ;�ނm��֫����-�Wa�hI�.nx�*�W�I�cЫ��&@Q��l��!�(nt�3}�<��k�������)Na��)�y]g!�:<��U ��[�W��"U��B��7��az8Y; :���`�b��w2�wp�h��^R���W�b<�j���6�,�Ƣ��G(�����%0��^�p ]F5��M�"0�6`ϡ/�:-%����)�f����,��ڹ��i��B��%� �|sW-�S�@����b�p��j��uu샹S�E�"�DK��qO���9 ��Lѱ�p�W���q*�9�I��eMX��6�B��w���(z-d�2�3�0�-= "6��;H�A�RYK���)�/�����=N���L�����6G6���-�>\�v�ڎ�=ԃ�G(?�
����1��}9v���'�#�� ��Z- Y(EY>����-.�ҷ���Z+��� ހ��?I��`j�%ˋk9������N�,��I����I�����Lk2��(g9��h�ۢj��K���OBx:2�pp��'����$T���xȕe<�M��N/�s�3d���RGh��EO�m(i�ho�����1�`�
���1ܷ���.�g~�O(�86�!��Fzъ?b��R��;5��2����Z��)��312�:;H�[G�%�����ɮSy9� ��T��"˝y���AdT�CS9&[�ծnٱ���q�`c=`�����Ě� ��$��zw���>�����|��eT���D��cO �RT!���R�xA>o�c��8-83�#z��6���_G����jB�r��x$�$,VLy�fM�HE֘U"��:�x�PNo	�}!8){-���5[ٹ���j$����fo���b��&Kɜ��k�L
�/����R���7�gǤ�teuu\�L��R�o��wr�_���$�s#@>v��͑V*��J�b�"R�ʀZ�т��g�sɆ�0��I��>�Z3�	�?,�bD;w���,��J�*�5�F���M�;{�]�����LdT��u�Ը�ș��Z�0s��V��{�-����,6ua�nq�k,]��հ��g�<n�cN�Rۏ����=r�U�]ù�h"��|����n�M�{��
@�z�:p�W���7!~��xQ��@0�7�<��Y���C�De� q@.����o���P]��ָ�ض�='��d�æ�mP?A��;�0�����A/Z4ú�� �����o��9��ƴؔ�77���oF���E�A�шi�K%��*�����P���o9�w�"<u����m����unY��휁ao6�oe�rl,n���co�#����,�_���(+�S��\	����^Z@O�8���>�BKE�Ձ'���۳�es,Ҫ�P�afQ�o�aM�\?�(bKD�|����4��fsw�����|_t+^!GKh��p^OŞߴ?�*����e�smY-p�M�IӀ��6�
x�ˤ�"$Pv���%�eȤ�{��B��D�2N���L��|�J�����ǧQ:+o�b��*P���@�״͇�-b�CF�R% �>jt0,����x�K�4"��[%F�(��x|Q<R�W�\��g�b2t" 郉����gc�iA���B~��:����i�zj�Rw2X���� r�x�Y��#�����&vm3e�Ó�BS&1&"l�6ĝ�n�э�Q�2���>*����g_��*���gMyI��B���{Y2��*��^3�HN����B)'�^��8$6]j}���lW��.}DXo�4E��W�F�}q���3�AfTG�	>,׭7�Ab���	Jf�t'(3��k)P�k�M@,Ph ݩ�A˰�"'w��Y��B"�R�mQ��1:U 27���W\���T���P��`0���qE���q���!$^�"@_��R�
l����XH6����Ƈ���b�R��4x�NP/���b�Y�������jd%�9z��.����Fޥ�ɱJ~OjsR��u�h�������/�Z��I�i�Ӥ����Tn������ղo��zk�r�F3g�i�@ڴՔ	n�y6���7J9��4��H���/Q��Ci{g\Csf�П���Π��7[~/#�4+��]��*�Ȧ� ��nS�@:����K�u�<�ڞ��~3JR��rt�1�؛���>�M�Դ;s�%��}�G��yT73M��o�.�/�2i:L�(�9�nӛ��y�E}�����%�mE�㣧��wS��zo�~~�E"��_$:�h[r��$�T7�*�]�����r;L��ު��oH�D��nTF���r+KH��s1[�Ŝ'� !���.?j�tni;�V�7��1�ԭ:���Q����&(�~�g�}�.[S�HV�K:�x�]�h9�}���R.��?	�2�Kb+�ǿT��,&_Io�7���&��'A5<E�� �*������.�+���f���{�_�(
��B���W��
��vI2�����:�"�����>�A��'��&�1�_]6Z�*?B9�bS%��:i�C��~��Q�[	����{����r�B(��{��5��l��!�O�����9�/�a��$s-1m��T��aN^�#����,��GΤ�j����)��gb�����w,���H�s�����ځ�n�:���М��\�d��K�h}���+Ln���v��s 6��gW9�>^��N�k���E�Δ""=K��%�$�����uΫ^���n�J�U�-*;��,�}r�%��͙�pl}�ðO�&4��Rs���ٙ���XT�@K�Ԃ�tR�v�C?��oK&>�G��Ԟ�Rxtvς��%�B엣Ŕ���z�g�� $����f~x�8J��\@M�Zp,ujC�M!��W�ߓo׭	O|dɘ�G-s;�<pq6_��,�>��F��'_�݆~?Z�8�����b4l��Kq����[-�ڪRe� lUs�B�͋��kY��#�0\�ÆO�ί�2=G�xP��C����x.�v���eJ7o��U�V,-X�0 E�s��'�e���]2MD�""�7�O��Gi�U��`rN���{��r�����'�m�+m/v�����_WK��+�fkS�;�hLw�WV[��>�k����V [WqX��t�R��e�����[k�(\k	���W�Rᧁ�[Ǣ�'7顱��_��đ	���&T��ז���V>FU
š�#U�tC7�%^|Õ��rQ�,%h�,(�Y�:�fJ�璄���A'[3#J���sUi��&W�y���	�듨���Vt�)�^�fN@ q��_�}� i�+�����s�+Ι�J���}�������ј��բM�9��� �����
ɨT�7,���^�Q�۝؆fe=����8�0Y�)^b6Y�O�M��'�]"��n���	ݕFD}��%��}i�������ے�T�Y�2qSv�Hp=9ۋ�y��R��ի#g�1����Ug�e�q���3��OUЕn�#�M��Nflα�AX���ϭ�:��2�]���	
A�v�i�*�P4��o?�t�\�f!P��BB��f$��R���6aۧ�9U���ٞ��Gq<5��C�46�̭V����v�'�-��!8@�W��ٯ���)l>��V�P��}[�{J,�N��y�]O}J���r$do��%n�q��Io0�iB�r�! z�N�v�+xX�x�BtBPfԅB���h���(SW\;~�i��.�7y
��J0=�֫��@�-�9�n���=ܨ�z����G��#$]m�es��n��Ku��Av��\H�?7�1�y�$�	���=/)p���pjh]ˮ�a?����j����F6&XL�|:)���T��5��
M����ў�9תu�ů#��}���1��@#u,�"8>�1NÃA�I/t��J�?s8�ϊ*!�f�F̏�ua���u��y��*�e�*���5��*�!��W�kNH�ԅ�Ȝ�?LD-FN��G$�M�ܦF	-m�A��(N���~J��:=�GV��JCF�"Qc��gl�ܿ��g8�a���6u
��.(!�t94���}r��BmUO��wiٗ`��2[������G	�x�!��j���A��>I~~�Ox�MA����H��}&�	\����v��C���M2gll�	$��fDC��$�r#%).�
���0���e�J�jW�۔� flI��{�G�5������/�b��pXV!(�׎l˄��j�|MrU�Ż\��ڕ^." ���q���[�,H�xv �v�#�ϐgR�HL>��L]�#�j�X= /���e<�8H���8���7�������AP�����0m���0��m 
֫�3jj�+�����7_���������+�R�z-�6���5q��)�'0��gQł�F�a?��Yɚ�K;�������Q�,m�\�nl��zA���!�)J���dFN�,����ˁQ\i����D�BU�tE�����jd����@]ʫ����C�=�]b������Xp��UQ߫=;=��o����4���3�O��L��P��F~���@n�5iAAL3�,�q�k�9����:}�+�Ep�]�w),w[�i�� �Ѐ���V3Ӟ���]{� ���)��V)�ƵI;UzXI�Y�&��fzQ'���y\�Iy��(N�e��X��u���.<��0����*=?Ɗ,F����bZfA�2g��ȉ��k�oa�����j�)aF3��7���ľ$B�s�ٗY]ʹ��"��q�K���Q����s(���[7�uNJLݘ�k����|[)�/��P��\�°,�ɻ7�v�7��R��Y���Qށ�vk���n�Ԁ�������դ	���[�#[.�UPuc�[�� ����`Ta�m��_'�cs��P���sm�dmż$q[�b�!� \Dpr��b�	e(���ak7k�����fD�MӲc#�/�;���7�#\1�d�4�Av�5A�8Y<9#�\sA�|��^���nw�&�V$p<C'Ý��fa�Y�cie�j�EPU��������<��GɠhS{3:�p�X�Rǋ�Ta{}jnm}8P��*�g��2@;��2	~���V�,��1�ZEMP"z
m����v�y�*��Ts�����R�.O�O*4���ǂY�� ����ݬw�g;%_T����s��Kf�Ӑ?�\�D�ύ����[�,��ȕ��5Z^��J���+��1?�Alɕ������b�"�Ȅ�<"�wp�&}g`e_~�]u��J���x��,�60W��`+��sʇ��f� N-*SS�K���*�� q�D	T E4���IKj>�.E�7��V�@�1j5N��<K�oD{���]�[���%�=!�D���v���B�
�4w`�lV"B(\�"�j6FM"���6]���ޝ�:�4 �CL�B������]���m��ϢB��v�K������ӽWG�>Ows�C�*�E��ҝ�@�ր^1=�󶟱cDm�����F+�;H4\��eO&^���b�+�/��;{�����$4����=��\=��M��I�������?q�+���.��8K�K7� �4���{k��l�b��&�Id�S� �F�ű0)ar&�/h���Z��P��ZH1­��ў��D$��q'��ݼd��}e�>
8�H$U�W� �Ջ��ݸUt#Az�1z�y�wT ���ZZ�~�� ��Y� �}^��"X��E�����6��sl�����SV@I��U�����,�m����5"���ڽ�%g�J̞��ʫ���u0e�d�����F��3���]x�M�	ČHFKC�فa�L����h��������R��I���eq>�y�H��%�fzZ��]�^���Gr����L,�����B�6�xz��%O��<%O�{���L{t?��6	��$��K\©2��C�[w���ݞ\)���-bO�gW�?�0��-&�A�k+<����#	�Z��,3�۷ǢF���c�IuJ˹��Cc3c�-���een�)���z��
��Ӊd����c7^�2�/����:�6����K=�L��9;��z��I��~��F�ox�Q#�9�Ћq����0~��g L����_��(JS��g�e����ќ�r9Y��7�@|�|±��M���z^��Յ(�ca<�m��O!�҂g^b+1�w���d�SM�:7�I��jaA�ϦRb!V�[]���{{*����B�˷%�߰eˆ��ݑS	�TkMף���A��sS)߿q����:�WOSp��r�E���#��C���&��$̂��d�к�tQl�ϑD�����8˃/�� ��s���yv������i='l>":���=��(]���o:ry�G y��b	��}`�KcQo��Z�d�ɳ�X�!���!�a��Y'��VHp�ޙ����b�|E @OY�q�%�W�������;b�ߢ2})�V��|��[����T0z��l%a?��q��s�W��ݔT�	e�DWvڑ0�|po��������d��WT=8��@ސʴ�{Pq�\�v�����9^�����`�̄����SV���t�F
�4ov&{JM�@���=#^��z@0��95L��v��Pew���g]lJ��*"�ɺm"*���l�7?F�y��T�ś�>q�3|N�//%9F$��}k ��7����Ӄ��[#�8��3ǚ�\Q1\�N�W��������1�5f6F�����Lt�j,h�p��T���G��<��Η6Ӌ�/��3���]��#8�/,�5�,�FX� �b(��|�N|��޼���ú�w���jJ�U�!��p���6_�j$p��?�G��J{HyX%�S����"��ԍ�t03H+E��M�Ŷ��L(m��;捧��G��F�R<(�Z9X��+]���܃P���ud}�Z8>��x�.֥�M7�3j��ж]����4s8�콙�e�3�~�IjN�g��'�	��-$?��x�)+p�2�*1J�����.�g�.��)�Y��hHB�G���8��6�"[V�v;-ǛC���$;"��HJ��:l�B[���"��	�Q��}��$��C/Iw�k�Ntm�~^]���r�5��ޘ��Z2�˼����F�H�A�.�a�(N�{A6��"kUlD�^/P�AGdO#5�7ÇHBcS����\{IRgK��h��M�N�1+~ �S���63�S�_.b�&���<��1������i1{.�t�#����RU���+E�lɐ�Wh�[4�����/��-E]d���v�� ���\�/Q�ؙ�x��\��p�e �(����sc����UL�����}��vC�-��t�
������nY�Nq������k96ЪJ
\���ʋ������	�=�r��f������!F�����R</b
i�mq̒�:���/�+�����h�{��:^"!��bg6�^G�1�m�c95�`G�:����֜�?��+�L&`iZ�+}]3Ӓ��<����G�?�C�t�R��k��~"��pd 7�f��Rp[���i��el��Ȍ�,�_Z�[Kj�ڪ�Fx��zb� ��҈*RｙW�;��(Ҁ7�ލ.,5�n�@Nw_Gޡ�����a>��FB&� �}�s���_�`��?�ҕq��ؘ�iԊ�K����	7���uyo��+��Q�5P���K��KL����p�E��'�As6�'~�+�la��,�U��L�}'�.��L�IYҥ�1�D��6�C��Z"�p���	[ĝ�Cp�s'[&�Q��FY^�L���'�YXhM�1�q�}��ڦ_�2��X��ɥ>�7���8�c ԓ�垲�2z���d��sA
�HP �?_�XO���JrK%R�w�;��"C˟*�����zb��[_.o	ڶ��6�� �ݣ��.���#p&��Y��C�MK��j��TY�ڈ�c���k~�
Vib˕�2�ՕQ�p��ZoL���`w��t������v�{]oA��9"+�s��:@@��Fz���N�ݧ�B��N	n<`���0���Ԑ��F��Z�.�q��c�O\a��2L��ğ
NO"L�p�2�VS�2��r�5�%?S&0��x�5�xkG�!�78%�6��I2s�;`S�1Qq��c���pP�%d��5�!b��/	�I��f�L��r�Y�K�����;�L�I�-j=\���]��u�RL�ΰ��P���\�i ���;yd��wk��8o�a��w83dgMufi�/�H��ځ�Za T ���i��&)ܻ�T�ùȘC4���~�к>y�܍$�+2H]���{�1�iy�t�#b`V�l~�ͿH����6��ZG>��E�5A�Ls�;��u�\K���b�bRGCYFE8�|��C�T:/^ey����.��3�� /zpp���tNO�ya�q����6�`luK�d����E5x�:�=����sf���TY	��mCB\a�2��<`�bT�(ee�o�	������dd�`M� ��Q�*�񇎺zߐr<�|υlX�k����n�9�0y��$Ǫ#�o׏;���|��%%�R�Q�㲲��z�և���ԯE��f&<o_-�A,�9�d��Eh�X����^'��)���b��"PNn��Pl�a�{=�E�?�)��5J��H1��9rդ��&�N�ոE�Z�՚�[mUV�0���=	���98R�qe�+x�������
z:��%�׍;X�QϾ���`s�a����9(�i��d����2����0�����n:U��8Q�������8��\���(�Tm3�����צg���+��- �߹�&�B�ώ&��a�6AN�;p3��aKڡ��0S��C�'�_GF�zq���L��c��ֈx���[ř��v���r=�\�G��F��r[v�R���|�X
�f-ڛ������U�%HX4L�5N�x]B�_�F&�j�y�^����(� �0ؐ���bz�i]���&��5�>�t,�v��$k(��ew�
���R]�4s�y�(���U���H���OR�����fq�wmu���R$:���#��󵯅$��Z��Ű�E�`���8��F�Aw�E{;\UYM��{�y�!x㤶d���k�|b��"l7�^´MI�?����E�N-6��P%�p8�\�)�>858/p>1q<��ѩ�;�#.9B�o�#����(��5~��~�����!�ƞ{
��N�G���ڊ��ABo�~{��ᶸ����s}灚!�����af��1_�64��#WXc��s#X;i��h�sYާ��B�B��&��I��c)gV!uO�z����������B���߮+���2��Ju0tT��E��������� �!b�Ů}%$����U���/�&�ݥE�h,M`N��k�1�4����7jފ����]OP��Wj��K���i渍��鴫��;N�����MZ=VMs�i4���]*@'&��w��A�^�&�M -�ߛR^K��P0�����&*��.����@��S`|J�#��e���'�<И��2�\��B����l����vd��^��C���I��٩��	�AYYF�O~�� M��VmL؅"۴�v� �p��J�{v�P���~�.�=�n�ե(�o�I��
�y���r5k��˥`!�������c�&�;���+�Z�TU���<�s�F�@#��g�@L@e��>G�%���4b����+�[�̜&6c������ۋE:��.��zqI��ۼ���I�l�7�/�����)�
��&��t���c�q`��a�g�\�,��� ���e}��8�H�x�#����R�a6{ip�&��c��%G9ԈG�m�$�j�gl��;�M)����(��!�/ņ�KQ��MxJ�~�ڍ���m�v�Cn\k4��,½J׹�gA�լ����1�����.QRFc�`����A�-������h�V���|3���[-�
T�y�-��u`N����b��-��K�3��P�W傧�t�S�:�*[ɗ3��4qI����J�'&�1 e��i��90�<bL��8qgj
6Z��^�lV��u_M�v�Y���XU�r=�f{+]b��nk�v�:|��c��܅��å��hsU��{xAػd`��[-A]*��D��r6u�Pa��
����-7 [S��e����Ű\�"�.��O�ޡJ��簘�*�R$$���>L䥾@I��-;en-�!�WҒ�w��X�m��E���vD���$��<�'P[i�Җ��
�Y�רh��V���d��\�y����CNܠ��TA�E���/�pV+��Ը�. ry��$�[h�s��7j�(|ɪ�2����G��Y��!�9=��2P������ٹB��Mj�m�5	����@e?=�W6���k[�3�&"n(�,��Dh��L=���[ȃA����j�}zQ�q�wih}��<�����&�ř&�� fb��>��kc�&�3`1�+\�ׄ��3
�B�A\B	^ �tU��J2:��D��@m�r��P�>��
��A�w������D������KԄ���#���5N��`��>�~W*|H��KC{fr;e3�w�a׋Vz?�ً֝�"�RɎ��Tɛ��xP�W�e5�qf%��lڜ�Giь�i��!q��u��+�:�ω�B0��7P#D�m���{|�8���|�10� D��\9Œ�F5�)NP��T�QpZ�E�<�"�@9��\Ҙ�\R���rUIi,�>5�A�#��Kq�����>Nm\�ٿ� ��u0kx�'×/a~��RN�&sB���`O^�%wVX�B�a��)��Ѓf�5m����A�CWh� _�9S_IT3A�<�J���j��g���I!���Ԉ$p���\+���ē?-I��{G�u=�ݶ�jti��ˉ�k�ȴ��Q4Հ�eY����#7"q;��ŕt�1S& e����0y�W�S���@��� ���Ɍ�'Rq��-����^����.���͍r0߽�]q��l
�B8[�yy��n�e�E0ힺ��F-�����p�쮞�Eŀڀ=�8����W����P��%
���ꤥ�pK0xw��]a�@�w
Id�7�ֶ4������)�+�l�k��
��m���J������Kb����>ת��^P�nz0t��?.b���`^�t$��Ѣ�B> p����������d��+
���.�ิ��N��h��s�q5^/^=X� w u�Y�����nxO<�*�XX�\���{�}���'�腆�#����*��Zd�H�N���Zշ4�D�9�R���j����}��)����ΤyƫeF���P�2������φ�}������ ����>3�m2+ҔE��ݞ�#��8�����h���6-��Dk�)��"KPHOʉ�?g �������� �����$=�Ѽ��a��ęy�Ԍ�F���3i�t���W���]�h�V|,���Qi�Q�{�(��k��X;j�%���8��ൡ8e)�ЕW�5��>>����4���d�?�Y:ƻ������1	�o_0]�]�k��^���\
���G������2�%TS�h3هC�ۚ������&����<~�5;D����m�������Ő�����v5*�KMdK����ni������r�WI��3x7Bi�:��6�5���&�f���3/XI��z���p�%l�v���6�rsV�V��[*k���Qw
D��i�*ӿY\����n��T���g�Sg�xi���%'kX>e�Ҷ�Hϋ����w'�z�Fn�9��e��Ю���<T���E�_��D<QL��2�L�o:d�k.�& �F�k�y��9�͈J�ҟ�)���i����`���.�#Z�����]���t�r�(�U�e�Q���� k
�uX\=��,�$��M!���c��ͭy��~[�����a�^��g����e��d�e�L5�p���S���Dr�w���	���A "���Yc����JAu}hO�7&�㇄61w���Ap���tΩ&/]{�=P=��.��県��F��If�b�m�	E�L^��?��xD��>�hv`�+k�;$�����|������?V Q9�Q��@U�u�Q,�����2�ѩ�t�l&)9*�N�H^7=���@Ź��M��`�=$��5�4���ڨ���SO��Qw���e����`�}d$$���1-~�[G<��c�-�P��A-�����[@��$�K�l+�M�ٝ
�]��5I�uX?��!��~A���޲���=G�5*�{�>�����Gj��iEX���IƳ����I�+�'�m��a`r� e��|N�҂ Z`2ϣ�v�Dڡ�3�n�����ƜƬ��WF���0��4| �O���R���d=��G�yb��Y������lN?��D�Kis}��P�^<M�~h{O��f|iV�Q���Z ҂�݂�����0ò�=�7/�,{IM�@�%V3��s����8����f���'PW�UɲG1����,?�R|=ОjٮK[�p(`	+�Q�ߧ���cB�9���d�Ra
�d�O�h)�2�^�R�r��R�d|r����ҫ�챙ȯ5s���8&����s�˂>%��M~N���!<��"��WP�H(N��̀bA�g��ouaF�`�Q8v%T�8)䫧m
�m�����P�|���e(�gR�p5�	�{�Wy��=��+���Z���(m�V�sפ(A&��^n�ax����2������v���7]G��itX�'ݷ����`�q{T��r�b��F@�SA;mF�.��3D�5�܂�'�i��G��:t]����r�|w��5B_(����wt��7�x*��۝�F���}?:Z����! �T@oܡ�!�|$��K�zs)��xsK����!1���2�z��5v�iǩ�W9�Er�r��,vE�>^������ �R�~�Ml�bZ5��k�jãؤ���w�M֫����[N_��^Pq���MR�r����L]Cq� �\�%PX���l���89���ĮJ:FH��i��#�SmRf-�E�L�$%���N~ǆ��'~M37	�z@�g�q���ey#�vAm׽��y�����a�������_�A�}��-�W�re���҅i "�����u��:�`�{֦�p�~�є|�
�$):C�S'�Kzj�7v6|L���i���:-���#�����2��P+�ǒ��O�YU�1����H>ٸ�]�3e��I�x,s����f��u���&�/�@R�\���i�w�#^^� ��$��d��ͺ�Y�p��kdl��I�H�K*�+}��L����	E;��Iɺ�
�?���F�mR�#�|���(+����s�����R��b����e��î���^�:9��P[:]��Z&��¯dE��u+�A���p�^|�-i$[�%[
�A���a��^���S�'i���������&h+��BiB�V�K��ZtH�w|'m�U�3� M`�2�r4�Eχaa3�$���8���N�c�Ё*.�_M` ��!/������L�:�܌"6��I��e.�E1�Ŏ��m�oPY�����o1�0�%�O*o#���K�~�W�vl�H�G�`)U7|c��|���3�p�M]��Zt��dT�\�R�专�Ŭw��WU�z8b�r����Y :��&���
�ٮ�Jg�
��]�+1RT��֡��Hĳ܂>�aƖ�)@�>�C:ڎ_�~�U㉡ZA��F�ј`z.�f.����KǬ���2#i^��Єe(恅YQ�NC��gk+�4ۈ`�9�	�1ގ�s���'S��I��f�i�%\?{�g;c�E*6�jb�1��S��>�[�	vЀ��6����zr���v�����a�\"z��F��5���G���e��v��}�h�rL�Q�E�q��O�q�'C���d.mDc��|�vQ*!2��~��J±e/��K���Ѷ?�}H �!m�^���V��Z�'�D��/Y��Ԁ��υ1�JU�l��d��V����jb�j����y��}�գ�+OD" ���3GDkP:/�bDQ��p����[�7\KW�|\����^�n��k]�`P�Ȥa�����Gʹ#������Җ_���'u:��,��Z-Р��ή5�����n�o�E��g�ㆴqO���P����)��ym0�b���g=c���If�	��؞��Y5%��)N� �#�5�2����٧-�r��.8h��y{C�lcU��iG�R����ّ[G%�޹⢇^z�Kט\u &A�QI�!DC`���ü��ў�ߝ}^��G�vS{[:'իM#���혽zI�uG�(/rQ����C�4���ӡ ϶S<��� ��1�sX��;�:�,�4(KF�������=5���i!gR��S�foD�:9#����k���I룺�4�����P����r~�KH�i٘���W��Z\�a��B�z�x!^i���t���?*�8=�$�f�(��*�',��]�E�[;/���X��^g��%y�<��Z��h�aJ�z��{͌)�U;�(�m�}���eI��YC:o˩U�����D�l(�͢*��e��b�V��+@	�7���^4�b��9|1>���I���9y�[[�e'��:�#�AW����_S��������A�sp[���y���0�:����u�G7�E��ʲZ�m�����&$k+����#�L�f6��
����[E�(����J��5v���(En?ʵ�&��`.�)йS��z$јg0$��$�7�S��Tкs�짰�4ɬ�+F�e������k��=�X���6UY�Ƒ�=A_o�NE����ꪈ�}1
��?$W��U� ˣ�@���OZZ�\Ǹ�q1u�I�N��e�S$u��s8�ѭ��%m����b4��,O,��C)��.����k������	��TNX����^��C=I�d8�א�M�dd���R�_�p�]��62 w�O�����gjq��VU`��0s�'�PZ�����=�h���#� �Vo�R�+8����CC^��pߊ���i�*�#�կ�dKj8B��BȗP���	��i�������!����L��.}�k�M��݌8�> *�۶����{ؕ���?�	�C�p��ȹO��Q�BE�th?�1Z��l��ռ�Hc���h�1fb�``s�_f��͖�z��iާ��E���/�E�������U�Б�+�@��u=5�B�zۙ�ZZ��^}p�B��c[�����MH��*[.�@��a� �~��C��o���<ًh?��t��n�Qώf���]
O�ru�%ȍ�o0�)�O�.�Y'�f��h/�'�). �&OM�,���`�u~�Tx0����A�!L*��)��Y�hP�����v��5�sλ]���ӄ2�N�E�n��8�P��核;��c(�g ���7�J�@$k��J ��/Z�)C�s���zYTl�;1[��f������c_�����F	������u�����0���X�s�S�_m��E=��3+{����<��C� d.�O�˙f�u�ʘÃ�|�T��O���R=+��u�EY>�9$ ��'������U����@���+B��*$a�f��pM��h&����Ø���̩̙҃P�e"&p��85��I��w���G[�F?~=�t+��v�M+Y|��}���Jl(u��qT�^+�k�Y?�٠* (��hj���I����V;�3FNp�j�S-Bf�9؋�l����]ӎ���K��2�x�$��'�t���m1��ڐ��LrNo���|�\pl����m��M�+�z�۞����N���uf����ٝ�W�z��`�1�)	�H3��8ߠt>�Vhpx�0�e����Zs�Q��ϛ���-��j��M���8"��@_6��p2o��W�;�;��B��~��.r)���3��b�G����rK�fA�܄�W@I栚��d��m�p�j���<|�|�*z\)�s>�����uk\:���`8�1�T�CP��OY�s4�]�VB���tm�l"��}37�k��"��Ӫn;�>B�'	ڥ�t� �hDd����KU�;=�Z���&g	��M�F�(�Ӎ�[�^��x"`2$O���UR~���C�s#&�����c����>R�+:s�<p3�O�h	/q\\&�5��J�@�IQ��!]��+Րx�Em?Yzl�B8O*�Tw��)���ʌc&�_�f������ǧď,Tn�;뇊n�V�t���ʮ�b�X�Q�Ä�-�U<��K[j?/g��lR�6�O��.{4?H2���	4�p®�э�g����M<E�M��Y4w|5J�f�pBcۺ�
������
a�:Lf��+�7<ꤧ�ݔtJP�!摒<�h`���XL*gC��
��`F�ϻ*�NO�FG�a`�Q��B��;��,��Z�������F��%�/��9�$��?�%?��H��J���.�8�s�Eb|�E&�FK����3Ϟ�
��I��t���O�Ӭ,p���3�+�4�B��"���� ��Wr����D�D=4I^
}��d{*�Ӌ�4���=?��`�FX��vO���2D��/���+�[�$�BN��Ʃ��7����������R��Xb���U�C
J��)�f&����:��1�k�8i�A������c_T��v�2���ֽU�M+��k�1���y��2��l/���R�%?vK�JC��(0��W*.%wg�6��T�6�-nښH�b u�D�-@��+k
CqLؼ����=ծyz��[M\��V���A�I����V7��1��G�����H��T�G-f*�n�'.d�r@�׈"��C�X��=����Y5�i �g�q(vz�K�=4aw=�ZS�"<�{�X!�8I�UP���4+i���{��p�n�����&B\>%)m;��x�: G���ɍ_�V�C�=�E�]��΀}ym����KǱ�Ԋ=/��B'��Ҧ=�.x�#���p�h��3;x0�cm)4W�
auE6STě$��D�׾��i�7I�QƓ�!���&!��u�<?�p�O���>��ا��Y�`Vo�SOEQ�c@��`���CW��a��bH���ZD��g���]f���k:1�jpGRj��)QpB����$�ڭ����9��Ɖ���4nƹM{P*! �\��}m�N�
�@1Wk���c��3�:M1�-d̃-C�������:uL�{@�Y���+�� 3��f��,�0$+h������Oz��rRպk[���F&nȆO�1�jQ��&��{r�⣏��C����/��G�/�!j�  �d��lT��1Ļ��x�~�W8���Ő��i/�aQ��}FpS�z��Z��9DM�-|J��Q5,5�s�\���P�r����������\���L�˞���>�vtJw��r�@����}���#��g��D����LQ�腁,�OS��6|Q�DG�_n<,��:ǇH��oZ��`��DX��*譱�v��6�s����N>���2;�E�J�?���r�5-:g�]a�.+s�W�c��ώ�'8��|�w�4>�'�<3�Kh����,��//6�8oO�,�K&�aˊ���p TC���S�f�D+G2�-�\Yq7���f#�F��95�m�c[FC� ��Ce��u�tBQmj�E9t�R 8���%�-5M�a���UC]����՝��ie���t^k��\��I��J�^̈��Z�Tv�H�� e�^�������{I�b|��ҁI�c^�i��$���С4��믋W�5���t+�����L��NӬ��~��i�j���|�C�n)���udR��aV&=��6ʴ�|i{��e�№`�#�1ʿ�6u ��1�6����A�H��v��`,�̚�)�����Yzz�87Aa0� �3��<�����ʴ�B�F�R��/��I34����v��R��y?A�z���>�ToG�S4Ĥi.ڜ��ڱ,U-k�ة晃��礗�`Ǝ��LA�r) ��M�����|�	+��v:l[���g܃Ӡ�

"K��q,Os��F%-����l��:J�JV�ct�Ϭ@)�d���2�������/�uh�2���rߴ�[��=\{�S1�b��<L����Z)�$�!��f�+�x"��&Zr��)Rh#�K����?RD^�B���䖸"����e����nļ��u��,�G򢞌��'_:P�֍����:�ր�z�?�v�_��r������[��W�'�ѮJ�+k�rX�.�>~f���䇉:閛'���?.\�S�
��K�tp�
m���QJ�L��Ԭ������é�˃���'\iE�;H��@u7+���e��y=�j�z>���1̼��m՟�zӐ�����u���F��cM�ȋ�H�ገ�R72����fH�,� �8	4����/f��9���9�m[ޝ��"�����I7T�ڪD�0#X�����[vF��i�H�%���-H�jt�Ԣ�sD)���N O�����?��oG�d�+�h��3��7��,M�?;,���H�?A����T�Ł��W�u+W���嫟ӫ�P�ŧ�g��"����@C;.P2�D5�S�\�ف��A͕�I�H�����'���,�=���1����+��a��Σ�w�{��Sxk��%�!3������������+�M��h؟ζϭ�]�hu���mE�JM!�u�u��N���0���9��+X{y���:��g1L�^�H�ÛN�\)wuBc���e��p��OO���׏�ql�N�'J�g�f���6��s�4����L�Q(�{��3auNS����P(�u'y�p]+(��懮�#��.B��r��#C^���G�����{"�x�?���hIOne�o";��tqW��u��=�����Q;�zPG�M�a`ˬy��TS��[6�T�I]��fu\b�,��� �=sJİ�=Hr0G{)�� �� 
���=�W�IO��su�P���F��ꀚR�{p�~kv���KN�
�X��ݐD
�~�7	�\Yqb�M�pu9�\~g��Y�P�_m牎��2iG;��)��h#%����J�\��L�'z��(��f�5_v�n�\/��Fc^ '�]�g����	G��-T�W���>D��.���kXҒ	ًr��ٿ�Itz�����ޟ�&2@]�lT�J?�.$��Jo��{:����'�����*�E��-;�ה�Ҩ�ҁp��j�\T��B�� ˀ����(Qfr�"V|@�H�5~F	]u�!{���}AW:�T)��Ǜ�����F�4�&��"*���O50�5����T� j[7p'"�H	���fe��dP�-[�W�c��@�ml��#���[]%\b3Y��NXlǿ$EՔ\=.P
>���x�lS��?h��stN)�;sv��@z��I�O2�9�ó���v1q��=��{���i?�k�e�)��S&��Y������]N�ױ�?󾕛�<=���ъ������e�^���f��k���OGt�YX45)>aڏ6�$f�Q"]w?s�⾼n������M�.Z����-�?�_`�!�?nyc]7��%b�H����YV�]��aW�J���:����V8.qe[�I$���f��faM����~	�e�������Z��d�V�B5qbb��:�\�_���P�R=z��|�sf����o�j~��mtN��}تc�h�������ۖZ�<��ZǷ���!<a��7V�CW�����r�W��Ύ����ѓ=z�G�Į�	k�]��3�Ʈ0\ڒ�Bt��*���j�:M��1�iA�����UK��dz�%���z2vb�xH��=��u̦?�j�"Er�=����߸�(*���3�׋�ĐF�_�r�+��4�ck0c+frYu��?߸y��A>g~.��hK��p�\�͛F��/<�|8[����(Z�:�t��fs�|f��
����R0Q�%|�[�<a��$j��������8̈9��F���b��x0`LQ)ȓ)W�t�{t���(�]}�,�7�˜0�\�1�K����G=�{Je��tJ�4�3��9�PZ�o#(��ީJ�	}�Ђ�z���T;���:�V��O�V��(��p 5��-�y$'������w͓��[og�+�r L3�C=���{�� ��b�Yˮ�uJ�!��T��煃RA�8�������&��<n�vA�W݁�	�t��
�I���=��3~�4f�'������M����<�L��'6�l�~�ʁy�����|�#fVQ�7&���D�(��^��nQi��UL��?��[Y!���m�@�<6s����dQ�m_��ƙ���?�\��t���WsD=)]�>�0w�4X7.n�1�|HݘdsO��+��lX���ʾg�����f̋v*�B*��Y�o����,a��%; ~U��Ռ-DhD��X���!��|�Z��h�5�m��B�<����N�C���6B��7����b�`�@�_.�2�j����CIu��WZ�{�Q=�E�27	0�ri���Q��,=K� ��P���<O�G�ў®�A����i��I���iK�����4tE�(p��95�x^	vPH�!�lw�T��*�:�R�l��s��ql�<RW1G\4 g7�VJ���x��`��x4��v�����a=Y��d��o���y�c�u�SŐ ��[Z�%5^�X�١�-"z1�Ѡ�e�)����}^#��f
-it�&_�!���n^���Z˓��!G�?��>..k�S���v��^:�&���o����P(�y�_�TY��'ѝ*��AE�3�ی����,��N����7�P���D#�A�f!:��	�i�t��9�a��"x�y:�R1�D|��A?��N'���ȩ�����W�����ď#�s�費��w��uj_���JDF�+���
��%J�,|q�%���L����/�H1L�������y�w�͜��_�Q� �+|��v%Te=��=`S��D��껑,"����&�%/�|�<��M����9a�\/��F�]=]��qn�(�m�*	�=;��f�;tU��%VZp} 	�����XFz�`�ڟ�ΎŁ��wG4�_����k5��u�p�n����S�:�\�7d�S$Y��d��t?"����q��+���j���{\pE�DX�F���򄩆��	~�}�����W�@�{s�N"|��3Y�a�Ч^��u>pu��UZ�� �V�.!���v#A�:z�~R����݈�E�q�l�}�|bXT�9j�ѫsS7xѧb!{j���D�k�׸SoZT�^ʰf��i�Y�&7aSZ4H��Ӏ����
�pV���_.��<���O�04\`h�sq�����{?ȸZ�6M6��r~Ji<�����݃�[*���0������细�ϑ��EcL)�A�ל6�j &���C-��H F�׿�8-������D��{����.�[~�/�����~B��5�)��s�b��C1Hr5kB�2�+���f�
RW�>-�'�X�Dz8F���I�lR�S�v|���l~��p����,��A�fk4#�%��\���P��:��a]C�S�kr?.u�һ��v�9��w�пK��`���0��\�6��9���S�󥔓�N��w�G�ԓ�p�J��Rjnk�<\���Nɕ\'����A �Q�r�7���=��e5ܷ�*X��Zt��>O�},���	�^Q�k:%���C`��=V��\�<C�jm���/��Vb�9 @
I�fY��%�����g�XG�ZF��5H���غ줝j�k���*%%��z�OB�"Zp��M�or�K���\޼d��e�cu�%�1b�a��1�yq]�b��d����_�����W�R<��:��oY+�s|p�/xMy)����P�ȴ^Kp��l Q�K�r�7yF���s�KS��	c:5�s4K=�<����x~���3�G�	Ň"&����>���4>MݹS���"l#u�,�;�ow��j8R���^��]f	�^�o
�ZB�Ϡ��6Q5��|�wP�� !&�B@y��^��������,�S+��z� �u�ݽ����y��w�ڠz�3���3�^���e���̒?= ����EB[�'[�)d�3��PY��B���P�m��[@���%z:��(���UMQ8�"¤nJy�;ś���`��I����Q��q�=�j'=�x�@��P��J2���?�*gh�YK;l_Z�iwsp���L���u[)x�T˹�e6�o"b=JA��1j��Р�9ڨ�>��)�`�\�/�q�8C��R��挬�`��,b�dC�<�&g���*V�`Z����T��Z��_�2NaLA�bv�v���yȎ����ޜ�#VS,ED6 ����GwOfP=�����(�dY2~��n�Pn?Y_Hd*�� S\��ԃ�ű7r�۠��wO����C^��	h�U{j��κ�d�n�s��U#c~S>��tz�!�2�ovU�K-}@��p�Z`��Ǫ��Ո9"=þ�е��ĺ��
���9?J�
�\h����Y�����\�����~���pU�v36��D����M�{i��\W}�}V$N���q�쮢؝��l��A���2�U�^��e��3����c������6��C�$�_ୡտ��O���Ȅ��w���؂���ơ��5�X��Dp�:��R�b�Qe�Ĕ{���I��W��V�B�[:�9�G�sM�a������I�v����O�e���NkK����SFB��<i�,��N�M��/
����+?9�&�y�]3��qb����q%�	�:���?f�޿�'{|��V'��/���Pk�RS�\==�W=(��\�f�=�?�6���a�M�B�X��3�f���s���o7�HiO�ŋ}Wd��F��\FV*-g�Ã���۟��g���@�	��	�T�a��7Wͳ��a�:�1�r[�������tC�3�e��Aj�<��̕�q�=�}^_�p!��!���)(��W7v`�xM�ٹ�w(+�$X��܈���N̾�h�atDtl��ti��Þ���<|8m��]�`|���*�p����?eM���F�������c݋��DYI�cA�K��8� ��2�!���!�{<Y�Ol�����B��͊-� )g�UN#���2�6:�.�_�Yk�쬌�Ყ��sʈѰ��.Ѳ��>��x���U4Q�, L���jK� _nZx��o����v�w
$N)���.S���Hp�Tf���s�=a��j��?�>q_u�m��:�A�`}�e��Qc,�4�X�A�vk�����3��Y���\��ۜJ-���s��aL�\Ը��f�|Td���<�D���qx���Z�%�4:0�/��|�r�yd;�W�'�$j�*��A�6.�k�4����RrD�;Xu��cM8 �o�N=$��N]6����A�Y�u'0Dfi���S_v҃\���R8��l㜫ن�����B�L�L�+1���k2�4��c���-X�I��j�PV��}�Ib��*��B�-M@�Ii�O�8�����W�|Y C����.n�F@�����j�ջ�����o�Z0�\X5�����o8|�	i��B�G�p���h���{�v;EHp��tjO����X��K`J�Y`^�E��1x���U���ijכH%�;��'�2�׿�zc��|��v[,�ݪQ���`g�U:,�37+�p� ʼ��q�=pk;P��j���GQO�V��|�Ŀv5��2�M��lI�R>A�Pyip�ԏA��=r�P�D��Ȳ"!{���.iWB��b��	o�����]:Sܧ���н���}�+�5	�KH%�?��F���w2��>k�[���!�W#��mi�m�<<H�KĶ�t/�������J��so&>�Nj����>��T3Q�.GƉ7�w��
D�U�ȕh��E8L�-��l�Ҿ�u�3��W(�|���lu���V���[oy��O.x�(Ho�z;�YQ��^�'hg�1�S�Geӻ��e�������E8vn���B�3ѵ��C�"xKcI\�:����yt��TOhrHH���.8a����z�zY(�`*AZ�����Y�?[|���n��z�s�x�Z��0�}#u�/�tb�À���}>�|eő�p�u^=<��ԛk�?!�{��Ó�k:8�J�k��ft�Ʉ��Y�����O [ ��n߼='z�XUps�>O�� �N���/��V�Z ���d[�V��(�Y�@s�������@=ę��<�$i�LȦ~{�v%��!1%u~���QҲ�^ȥ��z������Ϻ�i�^1	��ώ� V	�.6�,�Ĉ̢	�����S>H[�)a���t@���q	�Qޔ�xz[#�B�ad�����$��1Ԫ�Mf���#e��	�`)hq7�*�4o���.j���ޛ2]�o(���x�H�2��ց�q�����&1v]4Aؽ�jnZ�:U;`�'$��B��?�Y�<�bfb2��]�D2� Q^��L�&��y��������S�x�s�������Zbzх�۟�,ڌ�����ztK����GC�e�0����t����v�1i&��^��$��J0��)�PvWH�@M�>}z�X�b������X=ט{�n�B=m�\|��z��Sv�4_hX�\��-� �p�뺅>�A��f�Z[GK�634�]%��C�@&!�*����?D������� ��OK�h�Q*��I�g���n��*�;u�P'�lk��1g���$Lp�k	I/���u&Y�?�\�=�ے�^3Gߴ�vzceu�:SV�P)�Z�/���w�����6c��I�O C���E�(LBѮ)�\�Y������i�6�i�FG�����1O��]Sg��|c_��F�r}�\YS��
�x<�1M.�˳�kr��ѼRO�1�3%��dx�(�=	I���]*�Ch_����!�#��I�������_���P˾/���@��|0k&�̦	��W� ���b �7���/~�_/qqn{���2W�D�sxn5�n�Jf$.��,.�۩k��bT�
脷p�O�Q� ��,���/�E�r�f�^ H���!�Ԯ��*�C�@W�j�W-�S�]�8~&��"��T`���>:��պ�k�C�n�gK�M2T0W��ڝdG�����\Ix�yO}%
e�DY��ً�]����t�1Lz�~�F%�e�^�ڟC ���ES½oG�&�v>���	���A!
�}�U1�L�FW-bg��>I�cŭ�jFެ��ˍ)��k��̭��'��!���u�<����m�_��%^TϴN�W����b���G����A��G�Y���~�z�WD�<$j:c�bߔz6X�4j��WY#�-_Ó��3��*�L�ҍ�f�V�a�r�Сn!����[J�aP�d��T�%��
Y��Z�D�P�o�&n�2�z��)}���3z��KL�z��`8��0������s�7���R{��%�2h��h.#��=��W��O�2�ɞ�=��vb< 2HK$��oO[�o�ea_5���H�]AOnk���P�G�$NW؇�C�LDE��x���H��e�=�6��NY��]��@��K�?�K�5���N�|�N_�[�� ��Ld�~$k��0�}�j��N���%9�����s�l�I���/U*�]��!I����G�Ì�l����H�~Zy����)z��F^ޖ�坖 T �]�LPm�3�x��i�?ۚ��2��Kq*�����h�;Q���,e&do`}Ag�5g�*䬱RD;K+�/~�2���ǋ����J\T&.f@6� ���x�*i&2�q7��i�u]!1O^�\�+�<����j���
��p뼽�"J� ���~5�&���un����1�e�a����8ć�Py�i�'>����@�9$�����G�:��; �m���A�	�_6�H�$9@�u����5`1,j�5��7�x�c�L��8��<Tf-Oޛ�~�f/�ߎ�|�%��Wz����ŕ	2kbKь8�g�������2�
�.g�렩�}�ir��!É�f)હN�L]����"f3��Zz�K��V�s��lƌ������_��'A�@�a����������S�Z:ye���j�,z��T�\y�4-hɼ�@�	T�*!n��Š��,p9q��թ�zg˘K�ٔ��&ƐS�����o~��?4ۀ\!T{e�%����h�}e�%?0.�x��@��(�D��a��S�$5PM�z[l0w�\������O��XT5?�.�VM!X���hv�����$YG�.�/p�l���ψ�_*�" �^8�j.�r�mj0�̺�1=f�a &���d�P#��ڃ< �p�XѶ�{�D���{����M@�Ge=��q�c2Қ�w֟&��(@� �u��uJw�*!��\��E9�nnfL˴S?�� *ȕ�����^h�lA���`�>:�s���ڳg',��]q�T%AO3�*����Kp�rV�ƫ�Ű��H��[Me� ��WWM��� �b�`�*�2�F�~��I`O�ВE��4�}T�\��s�ڄ����j�$N���OkS���;,H�\�+�����E�ӕ���nN"���i��^[��������L:�E��dد?��� �O�(��.S�'��I�E����Fz$�|����Q����>�#��]�lz�o���\�VS�G(��5���|4^�;�~�&�Vx���� �;&	�ڰ�>����w�7� ���_��uy#�d���I�n���,��^ 7.����3�n���'�3a0l3�JV��3�V�(�д��Ux��a�3��������҇C��<��C}���mLPq~&��#�6�F�yH���,����-�V�/.!t���o�R���2q�"��	��A�n��ĕ�G5��c��ȩ�:<�VL��gs��c�7�.��_ٰ�� �	�9[��ܢ,�s�-E|th�#��ʾ���i�ܓ�o񶱀#�=S��s����F�Bԩ������zV�>`f8��N=��&n���5*>+���7֏��Rs���֛}8a<�>6���Vө_�w�k��r�R�yG_�<���Uϛ^����i�.l^ʀ���j���}�5���������q�c�7�hQr^|-����[̺��*-Mu����w'[���X���Ю5~q�Thz �,�&�H��]"���Hi$��n	�Q��+�`}�Q�R�LP<6����>ЋU^z��_Pu���3�!��a�pV��t��G�"��?��g������ڍD�zzC�F��{g�f]W#�0�؍{�w�n�mj˓��~�lP��/�dt�J���w�/�O$�m���� �����Ұ�M�߮�Z��%0���y��&�vv���_�gb��
��&�jc����� uQ���a�꜐�;]�35n��h��yJ簑xܰ�^�遚��+,2�E;�?�mN|���f"P�� C�t��\��0o��K�Q����vY^�o<y�Ա8��?��fVPh�UQ<�QzN�
��S��'�}�+K+�iy�`��o��ӦU�y]�A`n�{�'V���a��`!
�'���?��Y�[\f��k5ͳ+X�L&@y��褠k�ߵ�R4�{c>a�$�l[��>�3��4��P�\m���[(<�yY�o��a�{m�q��?�UG"�0�e��F���"����/��G��V�,k��eV�-�����M�W�5�ޡ��nX)�݀	!D�ƀV��F��A�$q��,\e�5�J����O�zŐ`lA`�4���N}C�����_���Ӽ��W;ȿ�"�EH#�g����e;1W0����v��@�nkG�,�Ȁ�s�}c�'��q�`h]Wv��a�P~7t�g`����R�n���U�F�g�x��앴��i�L��H��lO�z��(�UR�Ee��9���=ONι��i�´%e����W�
�<�wkӟ��1�h�y���a�6O�"��˥��bׂ��:���/矴p6��x���5�,��
�^a,�+2�2L�Vd�I�K�JM��n-��d|n�P�J�yz��Ք�/Ly��7����ɅB�->h��X"�!-��Vޕt7�]�PW{z�6��նV͙֐f���"�)�:��ᣎ�6W�y�	c�@�:O��B����"~]��G�i���̮���� BA{y��3U}8��c󓆏��1ϩz�-!}�
a_~�G���N_����%pq�߁Nm��p?���%�Y��� ��U�����K�-;9�$�m��ޠ�Hk�VD�"��y��z���ꗸ�e9�ݥ]�~ky>x>�d�3��p9r�6S��Sy���-ΡN0�b!J���ZE�'7y���vӌa���ؙ�y)��:.�~�Ҏ�L��Z� ζp��8�	�6���t
�֮��s�@)��������C��p�� %N�UZ'u�v	-�1Y��M�AZ���7ǐTC�G.���1w�Э�~�q�ǉ�ԧ$��<��3{;�Vh�>UfaH�̦��t��i#���%�*��B6�P�[T��OA�O�:��ZR::����V����|.��&9\�i�.�՞t|�o*%G�W>��a:�\/���ޮ�I����)�^�Qy��-�ƸAS�}V^D5���]����'�B�*�(ܫ�{K6�1�l�h2��N"��u��qm2�i�+�bh�5|ϪNt��AC$y��o��{�}P�\�5:��Nuh _|v����T���#�,\i.C�o�+A17�+6�������;9T�"�m�J��ɟS�.��t�k��W���A:�,��R#��ċn���Y4-�������I���a��V(��@�������qǽ�i��7�4o�$p8�i�Xȩ�9�ջ֜ �
�-�����ݐp�鸞a����C'��\��嘦�!�O�DZKh������j˥D��8��D�D^A%y����4Q7���i�r�";�WF�G�����ه��.�mh�aBw�^�	P�1��0���𔆣r�9]�>zƵH���*�"&?7�E��dI4v[J��j
�b�����s��)b��J�Fip�Q�C~��$��w���-���\%Z ��~�`f��kj�T��ۧ��t{A��a)Δ����S/�!�{���6��;��- k�������9
�q�G�&x֨þ�A��:l0�"Ѩ�B��y;%�H������]x�S�|�m�x`�4t�]]����4�����j��� @Q�L��|+��U�i�wW��j5���5�`�=j<��2����5ԫ;xlr��Y���G+Wj��������,-߾}0yJZ��c}7ڃ謀�׷�+��3��s�B���Ȝ
�H�^�f���$_Gb����өs�����z�7�q<i���zA�����[�h�h��^�ƈWw�����/D}k���[mT#g4���|FH%2�t6-qKgZ�|8���:>�9�����s~]3McMw#]��U�VƯ���z��F�Т8T������,���5�j�Q��)b��Ȳ���8/���� ���{3�oӄ�[g2�j�#x��U��������Ar$�3�p��,�56d���fҪ(f.��=d�J;鶧�6/{�uP	w����쓫�dq�K��?��Ӏ@�0N{@����K����AZ3�J�F�q�ΆTQA�ϴ�9��X~�ӽO�T�&��VG�X�����gY�IyE��+���C^�=����D�/�����T,�Y�-�/7jr��5����+|)��,�����+��d{����ۊ�{�"r�T���Z����.��D�J�v��ǜa�h5�^��a���rG�w>6'X��N��٬I�B�XF�+#ֿ�,\�E���㙕(Z�U��G�V�Q�4��d�g�T
� �Ԅ�Sm����gQ%�Y`�'yK8�.K*(ܝ���"f�䗃D�LA�vYe1�LՈ�4�5�ˏ!�!�� ��BW��Ӧ�6���������.�}J]^lUDlM�Q���W����dN�2U�A���U��ԩ�������zyk���5B���^�Y�X9:è�1u%m5���a0�$ ��)/����'Ӱ�"���f�g3�e�D+��ۃy��"�(Z%"v�~Tt��T�Շ��	
���n] �|d.)^�V���|�ֲa��,���1�U(֌�Õ��]���F��Ѫ�����P��юJA �<w�f^,خ9�����\vyW=r�vwڵ�so�O������{+�Nt���!}3e�]~<Բ���b|`ۋ+=��<��z/�{�NuX�8l� x����OXW�}����K�_�DP!-u@J`��tfQ�K��"B��Y k6�#9�Gmw��e_�NU���2J�)��hF�Pل��S*8)�Z�L��B��ǭ����I�J�2�x��Lb_�9��
R�H8OV�$f���lA�?{~�{o�Va�Lv��&��}8\)�o{@�Ђ�E{
����ԖW���pJ����(L}�ȋ��;��~�taj10�!��������ވ�FO͚��=)��և��zF��(F�ࢺDjדm�7C|F(�N��������{�N?��d7��:�!�2d�y�F�՗�����MI�Y
񮑚"�ġ;i'TeE�	��1�S�������b)�!|���k�$ʐ���׮���Gu��9�b8�̀1W�ep��|(<�ٰ���]����)�V�r��Q�k��n�u o�:@�,z�cq;ԾZw�˨�V���hٖ'Rŏ�s���"�!4N1�v��y�+��@�J���	4��Lн�AN����	Έ臾���� ֓��㧥v]�qd���W�*��Ea�p�:>E%�B�1Z��{�.�3�ֹ�$Q��&/$!r�
�h+wp�B�m��r���8D��%�qNbc�ͦ�o�#�I��p#��^�rjT��|�.��z_3 `;ak�k�4��O�zb����Åd'��%i�)���s(*�=��˘���zF��ʹ>���{?m>ҳ� q.@L�h;הm������{�[}���0�1�W_���ԃAC���WR7�����w��}}�)���CP/��x���:�f:O�|_A�/�97,��$6���*�n��~�q#�@m�y���&�e��\[d-"�z�a~�^+FP�0�I�l���q&������"�n��ƙ�q�#;�܄��~��F�E��U�*����̽�X8C���f�a�W˧������QLu�[aP)'O,�禐����q�����t������j	��$D���L����٢�~Ļ�Cv3k��^�1���3�픭�F�@�� '569��;�$�}��t�E--�6�dF�Fb��
?-�4h�3^���h�wϘ�n�5%\�����aW�=�m� >Fg�C����S�Q̞�Q�.c��;{*U��۳r��Lb⑃����9%�G̶C�;g�rR�8�F��HM��9�@X&_��D�w��L!qV�	�A��GW����L�y
Ƙ��,2T�v�6�XG��^kхz���D���2o�0�glw�ǿa0 ����KK	��i����E�S]�A�n����q}�]I Y?xޅ�����%�ՊC@m�ϏL'B�1�Xⷚf&�m���O���>o������VZC�W�0m��N蓏��K;�p	���yeC�	��z�o�0����^�sx�
&9�A��ϒ�f&U��C	�ȴ�zi2r�O�����2�	�xݦw�;uNit�/�광�����}���PE`U4��^?+ ����R/
W���sY㐖���I��r4Kr\P�1D���o	��V5�����">=b8���RW��5V]�$��s��ڣb���9˞ AcPl.z�Q�a#�xL#�{{�b���;d�r`�cp�& �G���I� �OPˌ$��osmU�	m�=�la1�Up��K&�	��'"'fK!�v���~6�l���Ξ�Kl�R�*��������R}�1R��<����bS��ʈ���ʈL���D��Zɭ ���"��)�O�<��G���iA�Mg��'Q�K��(���H�t�]�zn��w�ڭ��{��-�uc�h��.Y{�0[(�u@0]���F�Dh�n��?y�p���(�a���zm�B��r��~v�p��ǟ�m(�;-��Yc��8�P�0R"�KnDܡ�x��ܶӥgM�1���9��:�X�����z����Q�8��,~R3�1���w��z�i�p6��'l��4;�*�8k̏o	�-�N&k�������be<\7���:yUʛ}�UE�,��L�d��S�4���Y#G��v����r�׺H�����/���8,���S75������J%=��Խ��Gi�l&[�7�iY�jHmw�0\�	�g��_�%�a�e����2�Y��ۃ����V!~��� �%���vH��S}�qo�VO�s�7g{��b�}X?�$����p���&t����d=�!�����IJ�Q�#�%�`9��2.0`gc��9k���jr�%.~F;���	�`RC�aΑL.�Y�y߂O�*�Z��[��s���]�o,�+U>�8c���;*ٛ�"8v�Z��#|&?����mIt��0�6���{r�F����Dt�8!�e焷b�v�!ni�x�@�N�|n�Vѕ�Ud����!(�I }is�J����#ft���+���Z7,N���J�Xg��/Z��)�ä���3�5�cZ؍�-������6ٔ��������"�t"�Y�c?Rж��SD���vŀ��"� ��H�u���?����LC���h�r��[C��7�[�UH9ܗ���jm,V?Y�44R��_��a�w��R%�"�}�P���3�D��g���F�ܳ�'P�n !`�?��w�?��V�+�O�`�X{�Eg��5&9�(�o�-L�%N:��ú:��������M�g�-*Y\��2��Dk�:��������d�yMɐ���!p��:,;�{��@ڙ�Q�i6^������Q桖�hǠ+J�;$��Ƿ����(V3¯��1�ĺ*�l�����W����)�5~1�Փ%,�P��t�'�mfb�ϊ�i}(��$��pd�#��oc�*����� ]��� V�2�敁��!}���@�g�	V�*;7��!s���-�A؀�ݯh��gJ�{6c}�� �,smE�| � ���+�R��#�2WB��i�I�[�� �`4V7ME�(F�ؗ!\�<�2��
h���d�$�|�y����&�e�:\���7��:!��9�x6�����>��r�����@-�\�-���~�ԑ�j�����C��7�5O�&��Q�J0Ez�c�U�9H�Tj���>5�6C1������z��į`�#"p��c��U���sp&�!���}�#����P��\�� �Q��T[�����X�+1'VV(���O~7��b�P{�(r�A�K*E�Fp���j����s�qߑ��MVE�9��O�_��2���
ٶ��7
˲P�8�*5��������-s�.L����������H���:�X����l2�w���4A`� ]b�J�>^S=4��'��a����H"�㧾&����=[�p���`����F2��g�"��1��pѐ r��u�W� ���a� o�:�v�š����܏Ʀ?F�E�
m ��1��s4�X�'�ŔaC������8��ut|�@A��M��K/"��}����IX5+M�[(h��ӕ�+��s�'t+�!�1qLAx�˸�y�0+������)7���� �qG�������P���^�^�����ss�^T�b�
'���q��fe��@�Eݲ�p*)��ˇ^��O�E�GOv��$`�I���Mz���G��	pN����n���q��}�����ι��~uE�L�� ��4{�����Y0t$QJ�m���0͍�Jcf͝�������t�+��2	�B�Mأ�.ܣ��2d�N�a���M��1De-.y�-�[8g�fb����6͈��~
�%g������Tm�B{�D8�?0r�L�1@�����z���쒓5�0����L��= X������-�����ee�7���@�r�v\��$�[�Ċ0\Z����~�\"���	��R�]p_T~ބ��\ܮ�@»hd��K��,XB��t��ﻓ�� X_�9�a��g���e���g,��V�BzJ8��a#���b�[���2�5��ݥB�+W�
�����#()���of�iŤ����,ވ���O#�c��vû����k�j+����,t\�g��T�Cu��j �"wz3���iu<��~�c��N��*�OM���d/%�9��yφ��r��,�_�@��]x/�=��P��8{�v�ȄgI�}�i��H��bg�g���Dz�p�t|��y�.�и���a�[<�C�H��Tq-�����C�e�ϗ�&��J7����o@��>2^�3H#|2T���8�\OJ�����'��"���M�G�#I`�~%*ʋ,���̑��2�)�J�Q܀�.��T[7���:e෫��͗����'%{r΢]a����a ��1\���H�n�MY4���t�Ԥ�(2����0s�4��# 5"�r��3�ܸ��?��8�����>e��
G��<=)�mP�Ig�s cd���4|��X���1��T�LԄ��J��]գ�IW"����w;{iE�c��4�H�kP�l��T���G
7"��@�3x"��bI��_�C�jL.VqZEN�]�³�Τ_�����=�����0��+Y5O���A�<�E�����uż�e	�U$����gO��n�h/�ލUI|�E��Ư�6n��jU�U+@����L��'�v�]1����y��cSH7,Q���&#Xx�Tg�2����&�5BZi4+�8������3�yP���/<�>�	˵<�*���J^x���6`��鍘4�&��W��K ����'�(	�" 4�� y8��eHP�Fb�*��+5䰴��_�&��F�A��f��B5��P1�`$P�#�Hi,�H丌QI��(8��+ֻ3�~)�����,#z�+��h]^ ����W��}�!a�X�=9�����t ��>�T��n"m>Tn!��a�U��n ��YM�w۫d��Q� uYw�.z��u���5Ja�����4�A[ ��WW��=7~ĉ��9܂�F����X*�/g�5�Pl����;�\c�\����;�)��)��Ҹ�Ic��!㕩lb���&m��vp�ފ��h`T������b<K���9�.D�܇n8JP�<J��"���N�^�Je������(XQT�Kŕ�rJv�=T���{���}\"��)�\l����$*�	CH+��D2��߮j�v��|�'`%��VC��e�~:�]�0-0����Np��t�.���MG�UN�޴��97���F�'��Z,�O@9� �z�#/���q��%�
�p
��m͆@t���|�H\2�V����)~�$��ɻ*-4��\�;-�r~?��OL�sO��uRFBE��ncm ��]R��+e�Y�-��2�0B&D��ɵ��H��g+M�5����We.��i�B& �u]�'י;��'"_x�Mz��R��t��(Վ�x�_��UF��ė*��4��- �c~jXE~�Vl8N�9��	�\~?Kf�[�+�
}���؍�7��F�hvu^z�Kk�U#E�G)�oz��~�b�L�}��RcWf�-$K?Z��##���ͣ�`���M�eJ:J�~������[��<��BkiUfzW�W*�IR�`$;�#�G2A	����b>�{��=3���um�*�aпҌ#YFPs7}ȳXp��x�rY"���U6��Z�j�Q
r!d�\���8�ԛ|�JP�ȍ�إ�}�K}�i��Kܕ8e!ﰿ�iL�q��nv.�lJܹ���C�U�U{T>W�O���ֳܕ��,��]F{��4k��{e����"�b�L46@��dlz蟲�m���~�\y��R����(9�i6�}6�XA�m�w�6�3�D>��}C��ͨ�\ɹ]}&%7��'c�T������a�8�ސ��E���!:�(ܮ�^�A2)��G�u���αG�G/�����M��.��:ӳ r�&N�M�six��|�,���d&�b��7�<r�j?l�4_Nz���~�:x��xi�����f﫞^�U�o"�&1�ƚ��-㉕bjM<;�'�G'ӫ��I$��M������d�A�'#�Q�E<�]JH�����zA"q�\�B��1�U�'���[4��a�>�bP�.��Q��B�����;d�GV@�2k�>�!6�O���j�ӆ2�ƄnY�V)��Կ��2�	��_��*��G��/?���`�Bڝ���I�6X��MM՚_�5���b	��[����!�h�Lr�X�`����^��*;uKU���c�Ɵ��2�]�/�bf?e��7�g����\d;
k
��K�e�Uf?#=��O�������@M�e"9�ٌ�"ڷ, �0�E:�1�����%k��&����,rj(~�5dgi�k.7�Ă�W��d�����Q���|2��[j �� �-�ܜ�0��^����8��I���__�zuJ��Ѕ���!��
큱GhQ�.˗��h�䠼p��N���XJ��P\�M�����eI�i���t\˞r�3�Dǃ�qD~���~z�;u"X�x*��,�5��SZ1�D�$\�S�՛����.��r(0S/ts
��dK��1达P�����I���vy�A`���`O�w�]⢀a�>����2�K�ͬ� NL�EX�W�^�ۍf��(q�)�oc2�2����5X͞�(��tϸC�>�/�p�+�m�}�YM�/�7-��s�ou�1�j�Zbn�T��|f�ܕ�����v�'��ή|
�,i����,��{�ڽ<�����d�A�7�6�g�<�JF{sQH�k<�&*�S9�=M���_��J�p��V���Dc�~}�^ }v��<�@�ca��$��X_�?�~�9�u52�~���pw�t?O%r��ʼjL�����f�w	��TabU��պIz:�lYL���4\gb	���@w8\�I�ؑ~B@N��ߚر��:O�#��ൂ��,�?��-ߗ�.��'g!;=H�<,"t8��u	�'��`y����p+�K5D(�Mя��D��șeؘQ&Wm�OC���{0Y�鱇�k��^��q?�k�6�J��Ƕ�Ҧ���<|���TK+�����8�1��CT���|�Y����S
��C�+���x������+ө�^Z�«��5f�C�ބ4:�D����>�{��)��ҟ��78H"��Zh�$\/ݪ���'w\�J���V�З����R��hk�� �?��y���.�cc&{�'5�w�l̮����Bu!4�b�W��ݦ�눺��f�����`�����f�a��v�z����()ĩ
�4IWx���E��}'�ͪ�MI��o.���3i.d�:�WV�����iM��A?�D:�&��i��˂*}l�߁��-.����˶
��t�(kC&��R�t�)]^c:�^���Ѻ�hB��}�E8~�d�Br��&�k�3,���=�Y ���U>�HVMY���Z[I,U.��t\	�#��F��x��[㜍Mi���-`��|#Y(���x:P�ktR^ {uWB�-T�-��<X����p�l����%��Y"B����x�M��t���7�Ę�B��8�e����a)��[D+�<�T�~G��Rb���57����uޯ������TĆ"j_� G��Ä��e2�Q�T��V��z��=0V�sK ��w�`cxY�N%�_=��+��ڭE坂Q1%Z���{'�4�Rٻ�R����}�������97{�.���/�a����hv@R�e�/�1Ѝ�0��he���7�	k�t���nƠcQ[سw�^��Y���|�w���q��<�r*V0��f�H����z����0.�k얹�y�%�����%�ho4�`�R�L3t ��B������dI2Hz@���a����݃hYDB���{p�<(>�ր���XXF��/�B�Z��G����J�I����}��G$͂���F�����A2�%�f!���Ʃ�#k����5���y�WU�k̤9[S��D�Y�$�		B��C�d�K�j.�����cS/��W����B���:>H��>4����k����侙{)���sغ|��t^w�U�,o�[���ׅX����$ɡ�L׮���:�O7�+���h��WH���@Y���솽+�-$�/�����S��zMx��U�c�B��wM��
Q�9</��l�{�e�v�Xȍ�CS��g��[*|K��Q//�7�<}�.�B���7��6�	��50�o�ۅ���ޛ%����*	/M� ���9$���1���+�K2!3T��Y�L#�Z������qO�/�$���+޳�� ��S׽�Z��S�K��ČUE\2�	����KCr[;nw���6=��O���_y����e08���YF��"�\ ���Ō�̛��5(���)�:��,�8�N��ܯ�����l�דV��	��,���=��x�2��nA���҄�Uի���6���d�CM#Qh�m��;/»�����!E���Mޜ�c��)=^�'Xpq���9���H�;<�~�m�$��a����<���'�IoyO_���ʡaV̶�_iyz2d�(;�����ݘp�k3����&|t��G�M4G�
A���+S��|e�YH[?��T�I�F���s	Hl+�Y�Zx��Q7
����'	*��в��;��7����*��U�f��mA����9�6)nM�H�~�&Eh?�����;үv>΅zC�)� Q���=��.���� ������wPH��OWP4���9��x/em���g�'�S8��>�G0���ql�!a��45�r-�L�����H�S;�w����묮��]�� `��'e�8Gg����S�_^��%C�h�h�j��c�s���`��(Dhq.������BQ�8���:c݀�s���Xi�d�Taso�^���K��=��i��)(e7P!6�k��yQ>���ct�iv��oy����7�5��$�=����wf��88w�]fF�E��BxP��Kѷx�3S�锱�Q�xf�A�I��)
\t�.�Cܖy���|A&U, ��a�6�k�m@^��<I���zU�ڱ��~2�U�F��W��h�2Ù����'���"'�U��YZ�rn).�x+���1����i��	 �4U^���Y~�r��*ak�T����{�-v܇�$#Y�qܢ}ty{����-33���᚞�΍����]�i�$��R�Nw���1P?�Ǽ�ߢ��I�RU�f�{����ȼ:��/������yC��ںi:@��1�*}�ԆÖ�'u+��a�1��.�L	�`_�]1�Ӥ��o3p`isq�G�
����������M�Y�U��sn�K��=W%Θ�� �Y�����'9D�;����P����p�!/�cസ��q	l����h[���;��0�^'����`�cDp�໩�b}��cOz�-�=�P�Z�dl6�2�I�I3Q\�c Olm�1Q�9�0'�/T�#K�!�m
�д񼞶�$ʣ�CD�xE-��6�K���^s��e.v���T�ac�|��RZ��| ��HRp�"w��?]��Xzf��5c�H{�u�%%�܂�&5���uWdͨ���E���h� ��'7P|zJ�F�_q�E����8��m��(����h���8�G�rW_ٕ{���^����F�G���Ĕ�*��nha�{��H~>���0�;-5֓���{�u-J���bXøC�Ə�e
-D���DtubBu�QRފ�ί�C����mA��qS.�?���%|�ٵ�쏅��డ��
�x�'4*3��s|���h��e�1�Ũ�����Pd�B4�,�u���>hBwLt�-�]����QW.�V�*@��M+��V��Wy+"(��!���W8��0�6�EG%�۹x�7�H�ج
V� �T\B7���!ݣ�A��h���@����TF=z?���b��)��6C�f�s9��s����I�O�p�Sū�r�P�@��&fn�}�ɫ��-i������ 5�4除�h�.�i�:U�#���[�J*�0br�������e,�[�y�T�@)I���=K�>H� -�ZJ���r�!� E<���!�A�agW��ƖsY0r����Z�K4{�cr{��P��e��窩\L�l�5v�6#��j�34�e%���z�!��y� �lled{�(Rt;���K�	�a�k�mo<}f?О�PMq��"�i��CHA`Lߊ�XʁJ�9$Ku�Ԥ������s~�+�OsD:�������<��9���?h�]��r��){�����RI^�v���n�B��D�S�´O�z&ߋO<�-�=�)^�~�m&�`ľ, �����ړ�.-\�4<iM�H�
�O�⵨fW���3.�r�Ù���s�G3g�(ᐠ@-c���j`�l�;���)Z1�
i]�G�	"��:���#�&V��3�!��5�̀� e29���V��[B]����}�ZG�\�#��y�\�2=w�r�,@l�����2ZVl�Wp.t���`-�L�0�^�*��� �E��I��W5\yӐyY����Rwݍ�񖾣�_#?ԈpEQl�V�
�{�_$���Kz�'@�y�Cֵ��Ϸ#K
՞/��w�)E��i�O:R	��L�NtZU>Ր�h�����>�^����#G\�h�i.�^f�K'0i��%�.&{��������Bמ�xHϻa���
E�ZU�t �64�*|}C-��$�2+(����JK�#g�س�0#&*u�H��x�+�8��(!"0㐜h����bR�8��;��rv5c��6�N������XU~�	ʂ֊eGPM��Xw=e�"���c�|(��`�p�**|<�g!�G�I��U�R3����MDNزy?=oQ|�"�8b��΂Ӛ��c���J��z0^�[�Cs`�`�L����P�������8Kcۘ3�G^�L{**��HG.���9Vy���J���g{�LC~h2̠ؐF���o��z�������'��~�F=q}����d))H���_�q4�Q �u��s����҂e����d��`H�D�HJ#fS���Y�U
�W���"�}	r0э1ͩT#X�0�=Qa�,�Kd_�%ԫz�cV�#��x���1	N!�K��r�q��)� ��yP��ugz��E��͸7o �z��#�+q��D�S��tf:��.�3�^w���Q8\h�:���!aٿAj5}���2*�2�

�u��O��s\���S��R�cX荘_��Xh��B�h��D֢�;�1���l�ڱ/��Fɧ}�����#���o����/6#��� �?��]�︙'cY�g:'G�?)��cx��S��+q܎��کe��B�+�5�4�`���PzR�a�/�χ/eY[���,�0� /�pn��Jt̳�2�h$��~J��v`���1� &hLR )X�K��`��u3>���W^��4��$a���YMg���_w�(���k��2y�_yJ�Yy�_G޿�y�g/��1��¿�{��A+
U�	�7��h0>�LU�WRN���2Mcw��z�y���n��H��tc�t�JP0�]����֜�=��R���N;�d��TT����tG��0��@\�MaS�F[?'7 {S8���5!z;f�bn)y,���3�WG)�����v�@��u���X��E~��v�+�(^?cW��(��'`Vgg��ȟ�ޘ��%�FeS�1AJ�f�l����@��.����L/�)��*.�-c6���i���܀Q�a;:	I�'K�ʠ$Js)\0*�R���	�Ȁ+r5��H�cІ
���M��5�s	�����;�:8-�i�|	���)M=�H��M�s��=��d[�2>���d�k?Cݑx�RO����q�@#��qs������Sd8��4ӽ��.�
���o�$���E�Yƽ�8��*��}	���t���/�GJ`-#�XL�]u����T��q�Z�J[��(�������K�:���`�6[D$qC�o�D[>���Cn�ݱ2Q> ��Z$> S�AI�D��y�]����V���Z�� �g|�FM�����u� 7JC!�5%\a^Y#��6=9��yԏl�K�5�c���Nk	���^!}���¨�ٽ��+�PYmS�S��9>	���"���{����O�B^�w�~�2+��`ې�h��y�}�Ъ�`�a|�́�}"{��#���J'�9S�!�y^��R&���\���7���A)y�m���NW/�$Ń{;a�=�PҀ��d��
'A�����2�9�jzr�C�P��v9�sꧯ�[�b*�hO�2��mj�b��*��-��\f��>.7���ia�D��h�3j�y���*�M��q�02�ҥkE0m#t��0�	��ЕV���H:�˸e�0P�kw�|^C��$o�@~�M$�{D��#�v���asO�I{M�>�K���{=n}IPG��#�r���i3��p��"]��s ��fU|g�.�#�~��l�>�'��,4ֿ�%�T��̗S� ��&\=mV��ϪҐ���Ai��#"��B������j�kP�.婢����5�`�I��J�0���6��$ml<��gu�Q�|M��u�B��[$LQ��(*����_F��C����q�Fܧy�;����B"�M3�#���?`o���k�^1ա5UfL����
?�C|�rah�x�--<B;
����C?���I�K�������w��ݹ5Tb�f��9������d��.(l*ok;�ƺ�7q�y��J2���תunb;4��3����n��`4B��z�}1F*
UĦ.��Grk^{Ŏw�9n�}�͐��υԍ�9XC�Q�-��q50�o~ϛa��dT�1�A�uk�̀�}�JÑfq�A7{,jmv��;�!�ZN*��Pv��nhMǫ�Qd%�,�YTW�@j��O��c�������y��@�@��?1v*���S	�ԯp��%Y����Zk��� _r��|^�3����J�AP\9�V�va��6	a/�M��*{��\�M���j���σ{��6�z֡2���	�H��0��ݶԈ�C���啛H�QPz�����O�^O��f�Z,n�SEϟa=Qŗ�6��oY;d���);ʾ_��H�g-�[���'�k8���Q�|v�.���u� ��>f�sW�<q��N�7�ո������?l-�u��*����9ۦ��Q�2��j菩}���Fa���OB���/�$g!�ׅ<5x�pA�"�>J�X�f&��l~ U٤���a`�Kw��R%T6Ϣ�x�Re>�@gA���L� #h)��ߣ�e��퓭3�\֣č�=Y�P�R6r�rݫ�4��_/kW6���mv�3����'&��@@�g�~G*@�8�����a��P�}C���\�6+kg�S%.Z5��	ux{Q5���'Ҫ'Sh&O��;��h^�sR��tJ�({����"��]���{���ͧ��\�c���a��E&����q�1�GF�4��$��*��.*kq*�K`\�!YP{�u�'c�	EҢ�l�,R�G���"KտȺzB��>�����S8��Z)k� ��e�����ʹ�-��B	�l��Od<B��]��c�����W�;Ԋ�/�F���Ѧ��;Mxu����"O�X�uQ>�?P����ήE}9����bG���}����_~�����[���ӹZY��'�Z`�Zrۖ���o+�̭�. 8����D�r���ixk�kӉ�b�q�>=�_�c$oue���(�m�*���J�'���
_�m�x0�Բقi�
��m%��	�UHK�\e�"����6���/��O�f�-�}-��{���qo^��	q}Ӻ�DE�EkfZ���޹&�� ��~�Lj[��G]��\��}�l�jǛ{�b��$Ү����`w�݅)]ɀ�b�͞��.�b��bQ�+��<�M�n��~n�i�dے�<okq�}N�n����gЦxb��.}����НL#TS�}`lX������N�:KL�Έ��Q�N�}m�K�y%�O��8�I/]������r�)��U���V+f��_TBM|���V�&^7Ӆ]��&M�Cm���mJ����Fvj����/��C�����H������`0Q�8G2�@8K��p�S`�lJ/��5��q�;��J3�U|������g]&vM?�ĝ>QQ��*��6{��0�#�"F�A�W�썉���1�A�=rmϯ�'��7ysԕ=V\�+�Z�dzM�XO�Y�2ȼWH�:�>�m�5���V�0'{k��_���{aL/>+���~j;I����k�.���dh��S��U���;l ��Tݙ���M�X GJ ����յ���Z$��+�O�QeМJ#&Y�A��(}eY+��
̞���N�<(,О�+���bՁ���������&�c��.z����S5L0}�� ��Mm�)�3���؍��Y�O�q��'�K�W�Bᙐ�~��K��֒��d>HTC���Hq��ת�D�99�h�q�'�_� Of>o��z_X�ʾN�$Jes���@\�ֳg���)L���h��B�k������TbJ��$���M˄��*G/	�h�վ��#<�JNϺ$	�8�drff��[@R����<����{�z�F�a9���8�v�Qؖz��}�|X�j ��~��|�8��S��F��;lm�]�T�͊�w74���BGsD����y1�]~m��Go�X$`e.���ǔ^ 
�B�5l\|��5.�[:�XV}��\ڼ���Mf7&נ]�E��x�&tCP>7ն2b�Y�71ؘ��j�L�+��a���r��[�v`V�� � �o�틀w�y��*ґIf��s�����M>%'2��߳�?٩T!��$&.Pp��i�x��
	���)�{���O=
�%wi[Q��U-@w��-ί����u1�@k����1�T�8怿��2�~;9,��C�E����
��T���p�}���e� �EW&�����6��t���X�;dh'�v8c����i����z~��gbv<X�� ��h�j����y��8�Q�`�N��wE�#���_��L>�=�������󠱮�N�"�'�������:m�S��,2����Kі��1�ӱ�xs� �0��_6���&YEW��W�=Θ.U�����cҤd�P�&���Sɑu���4�rf���a��rL�y����@�ܬ9��%)�	M�l���7F����ۭ��Q ��+E������F���R��W��ffhe�E����g͝=ʄ7s�Уuu�'m.9F)����cjs*�d���ǝ�^M�\�W�nCH4� ����A�����/�^����aěd�BO���?%W��ܲSh�\W��bLܼi��q�����j��E�t�y�?*n����4�&��t,2f�Nʜ\�
�b��@-B�7�	�<h�JK=����g�}H'��}�!r��pGq��g�48�ǅ�NQO"�����se?8��谪��W:,����e�
 Z �����"P��k:�Q��F:7Q�N}����!B�#� [�SΫX������#8�蜧dK"��Ш�]]Q<�����u���������H	���4ZO�]_�+�4��|�<��Z*L; �DFJx��R��R�0n���:z���jY�{��'�m��h ���I�p��k)g�Hi9�|-�L���
�i-��Od�f�h{���UC�����Wt��l��L��9�gn#kpg6C����
A}!�v>(b�T2��L�8�2>��ñ^�Zw٪^��9�1�+�i^����\K����TM��K~�Pݪ���LE��u�k7���#̙���}�`��PN�&)�

: ܜ �̧ê�M��隣ǻ�Q�����NسxΖ�J��#���,��M�T�A��b&r&��w��I� n]�w:'�~3ޭ��m�Q�I�k��ɟ=w�fo�/)o��=�dKjfc��R5f��?c�kf�uXD�
}�a⤠(،��	��u�2��#:�&z֑�	�R�>3��V��=�����W,�C:j�K$�b��v�x ���-�Ou6��X�x�mk�Vÿ�aK�w�ZF�Y�F�?����Kq����Z��X�O�DT� ���t�ʽ�\��(檅'vw�\��e��3���	�y��9������=6(�^e����7Mi��a.ވL�7���H4��R�ޣy]�ݘ���B����7AN�����ʙ[p�ֿZM�i�.9;,�u"�P�\)��Q����3/�2���Z�@<tAœC^��i����	��
~t�l�^��ՋSHM�L�*?O�4���G�ٙ@�f)�:Wr��4�j%4�1��G�%�uV��^X���l����S�����P2��([m<�)������j�D������釰GQ�,U:���=����f�a����N�Z3�m���A��x�ET�]A��߸��:�C�Z/�B�!zq�(�5��"}C*��j�v��1H�~��z^K���a��v���Pfmm�Ι��4uȮ�F�� �T>8gy�Q[�?[�?H��]	�Ռ���;9<q�����)�w�l�	���.;Q�Mx ĴE�M�D��G�$�Y�K�����7��k3��Umύ����z���|x>�M:8��U��?m�L9NT�UNh��q$p���'��F�5P�����h�?ю��;+�^吚���t�N A� i��DGhF�ɥ#s�O6DS��$�w����n�X��uAS�[��\���]&�H��%��5��ȃ��IE���鴀6�沲��q˶!J�!jZ5K��(*3a_�Er�e�_C�uT�|'�h��Kx"��Z.w��1Fm������Xv��k΅���yfH�ױ�s�g`�_ �����cga�e�v�G��x�.��g��(��\ppq|$9�Է���\K����7G�Q��{:V���� ���1��A$��E�A���r���l5��q,:��{��r0AoK��i��O�-�}�n��S~B�8\��C��iܲ�:]o����W���Y�������K"�26�����;"���=}��[T7����)l��ma3`^R�5�x*�����~��OL��� �є��|�+��^�5�K[1�k��ݳ�㙖�>��D�p~^j��[�&�������oiMy"�=n7���I3�|3��!�ҝ�}P�����;������'�/�ΥJI8�r�͵JK��(���6X85���C`��5hd���ۢ�x����s�"B�%vX�jV']0 �1E44悁6�ݬ	���U9$i�"K�����$<�}FF����+=|J����ӯ����
���5�=&�Z"ZpowY�Y7�r�5mD��W<��0�W�frF�p����W�G^���=�otє��U��+d��p~�+.vj��<�Q�P���ġ��k�`c2�W��"[ySa ^�Kɯ_P���e����2�8Y��^�p�|0�~9[U��K��s��B�-�nޛ��w����ʵ��
Z� m�_���������8��)V���_wy�2[8�.��،�Q�M�uY�� HJ������m������<=xr�<��4g���3牻����ԽxdS���co�K���{��i4�`�z.��	#�&V��a'�?������-���WP�X��v)�vH��s2���-��ĐS�v�u�%�S�a��nc�>D�\�@��(��}̭	��\AZ�FĊTE|��_��u�(���/��K��k�pD�x���A��L22��^�n8�Җ�P�=�IX�7h�;Oح�|Ի�K���@�w�q�K�oU���5d�ci��0j�B��=�㤪j����]ҫ�﯇������U����V$����|F=ة�Ga�8י>��g�ܗEO%���D�M��v�'k{�����zQ����r�PU�����_������ӫF��<��-�w�zCS;h���OQ�mV.�|8sD>�H�'UJh�v�r��d�6r�_�P�9	+K�=�g�uE��4<x�*��$7�$���R%�:��������Z�F'�&�}���/b�P��
���v:�W.�6���j� ����r��O���#� �B�t�e0(�&Ƴ��um�R`h([�y����yF���:Kv2ԁДn����q3�[���z��s��D6�tEe����'n�y��Oo������$���G!���ӄCp�@���&B��X>Lw2�Z��2���Q�'� �4��F8`�m��-KjwpA�K�x�ۛ��w,�i������nMǣ�B��ۮmQ�X.����K��&HrԙRI�􌁺�,_0jl6�`es�Cـ.�'��&�;%%����!�#]m�J`���'F��w
�P]�љ�䘄�J�{R��q	݁p��t��e��nt��Wx�yl;�`L��:�ӽ��%�M4+�x/�@�D�d�%R��f�9Gn4��N��p�Ә�J�d�"����4K��%��� ޴��8�+���T<�ХO��W=l�����̋�5P���#
�Ez{ūʶ��j|C�t5ft�(����'&�!�X_�*�?m�ܤ$�/�,R��Ch����7����N����$��6�ej/D�%�s���>�<9����C�Ϝ΢�[���G���-4;j%�u���^Ga�S��~�2�S�u���b����w��z�Q
A�@:�G�G�V������"v�� d�'���H�<5�H�J׮��[G����g؊~��@ 7�V��Td����I(�oY2��F��ཐq��`���U�1L�=�-��Mvo<	k�D���|h]q�^j'�1Gj���Bf��Y@���e�_<�~qF�,� �X��4�\`��=���$¯G[�5���g����\�U�g��j%.��w�D��˲fNptJ/yܘ�f�Zs	�c̆Ĭ�n��g�2�.i*ؿ�:r��1�����
��TɃ�;5��u�WN dr�q��&��+A-�Uڵ�c��9�3l'�Ǌrz������(��l�D�IT&e���sY�W�O�'��s�9�$����������4��%ufV��i٠6{��;���;��Wq��kX� ��r���û䇸9v��pR<��E�|��QF�2>Om �$\�LP������(`�";�Gmp�K��w~K3���67B��������鵡
�8�t ��]�S�Ҥ����D��_��I�ӯI��,��{�|~�O�&v�����j�����딘rc�Θ����C�Ž r���LO���I^��mqD���ѪI!G�T���>���/�hX#v��In�}�5�3\�G�14��(����-�|�#�G���
���f�w���c"���<v����]ҰtnD��u?IQ�C�l��W�;t\:�Z0Sf�����s0��'.nQ�"O�ƄJ� >N��?��&������C�&�6V8���Sң�����*�>�Y�+�O�wj%�����Ȧ`T*4#�����ˇ�����U˺��nA��+V�*\�mv��
@�D��.,�\hp�w��ע�������3��?�
pks+���2��@�c�i��$��c{_m���e=��c#�v�������;_��'.!d��ԟGx�AU�g^&(������go���k��{3B��[�җh��n�UKI9�올[������x�o~�_s�5n�#,��Q�V��g���fH�֙��Ф!u�J�p=�W᱖;]0i�.�y1u$�~q"����J��cA���`����C���l`ߪ/_���zUj�v���ڇ�c�	�Fٷz.W�W�
~8�����2�䠛��|+�����|�}Y_�����j$5u��
�F�����!;óB�9������A�ZF���c���%O�Ik�HBf4g�k|Ќ�u�8���^&t{���[3h�+�����P��n@�a2��9/�7�������e�������>��РT!�k#a}X�2k����8���1f#�X��Ɓ�ٖ��)ip���@�79Jrsq8�2�9Jw�B{�<�)Ac7(Ǒ�yA�Gk���v}�������_��������%�������گ� i��7�ߨ}O���r���l�)OE�y/�M��s�8!���]�S��?.D����#��kn�@���YVt�%�1�Kę������b�ʱ5j;�&"��m&�m4W�c,�[g%�Bj͑�'~���MD�N3�4A���I���S� ~(����o
��GX|����$�X	�	cg_��.�r����&�}%�<ΰF6'�x�6-�5n�,�,l8w�@1l<�����BV��|����ݸ�'�9q!�V�}S����)��ˈߖ�����z�VO�S0�F�����WH�]�s�ȅJ��k�-J�2��#i:KR�CI�[�(a��X ��섑b9_4�2E��R�������9;�u���h��9���)��co/�
����j�Ɯ��̨0Hv�?߃P�_��}=�m�o����UF<���w�d�����}��!���T^b���Q�0���\1X6�H��s�����i-�Bs��%HԶ$��y(Er��}	�26%;������elj�G'�Ħ�Pr�����]R�,�+��3v4�	��5@�TBy�;M�O^�<fҫ܍i(Y�M̦n�W�	M=����¤Nl��J�;���C��s�ߕ�$x7S7(��cЩ�3\~��#��fJ��yr��p ��A��k��	7�6�pr>}�v�����{�p�Q	i��R�E _��;n)2�������_��J�,����t�ȏ-���F)HA��G
r��Dl�ݓ�� rO,oYo����f6�ch���fMWco��Q����:���o募9>�Gi?Wn�q`|��y��D���{�OÍ�{��؆y��\�Y^[�)���@Q(��̠#6�9kE��vŕ��A�k+�SP�p��pY��-�X���5z(+Ҫ��#��X<���͒Ik)m
L��)�Ax��*#AEK��F񚻦5���Jy6fuP��/�s��!,�=w���\U[U�Y�Q4^�G�z�2�_��dd�k̈́&�sɢ����"aVN�M�K㾫��)�l.Iz���l���aTi�P�H�$3�'4�Tc��M=c~2�{�8Ȱ����+�9P�Z8q'�g�cF��wLiѺ�}M�P2oo��J�䏩�����G�B��ǹC-�G�&9�sv��#�.����mv����8u���G5r�W�RN̋Y�n����b��͡L3u��=��>��[.���-f1�G.�4M���Q�K~�zǔ��^7k�[�)_���U�'�
��� ٷ��=� =|j��Ӏ���ۘe�ٮxr�0T�	�n�������ш��Oj����Zs���=����*���v�U�OP�j����[x�9�G��.���֝(V�������)ť���q��X �w�<ɥ�aSXgDЬSgU���Q��=��+2n����cT�����e1�[�^�+q����͝`[hX��@��Q���e>^��d�{QQus���#;Y�� |jˎx�0c�����H&)���`ö�:��W��u|* "h9���������bo�������D◃��>��� 
�\�S�C�.)@r/X�SfE�ر����	�&��V���[끊���K! X�N�]PJ�t���m�0�n��_�I��ٺ����m���V֤�Dt��0�7_�5�F�_��R��[ R���C��=�u{�{�����C *boq>DH�ip�,bj0ɒ��^D.X�V�o���d�tS��|���ot�����e�i��#x�龩;��k�l�-�3�N����@k�ht1��h��zq�``��m��o{�w��ZL�@dyoZ�!���	��լmg�d��<��\c���mՂQL� �d4C,�<S䫓bڏ` �Ӹ鑩�b����H-�jis��	�=e���kE����Y#;4�VY�J3������ �2f��uwM���W��?'����O5��!(E���׆xK�'�=KO�@~��H{P|�xO�JT��p��|
D�}M��{�����5��fQ�>4�Ae�����˷z��J�ڌB^B���LM��3<N׭Ñ�՗�SR��pqq\'?���M�q��M���������q�1-(�#vir���ڹ��"�אǂ�����j�<�W
����ֿ�R�w%�b/4��E����vt�p��<�}��R_yH��NZ�K�ɰ���0r��g��#���K��ԕ�b�l4��C��єL23}H���=��lL2�lI��M�T�W˿3v��gnĞ����;�`K6|o/LU߇G���Á����^�HWHY�4������K���<7I[��tj�~�MCTA��)��e��"��F`w���IO�!tM"��)�O0�U`B�8%*b�'6v/f�z|ԝ8�7���!"+
4F'�_.�&�a:�pמd	&�o|�e�\�c.�4��Bt޶~pػH��^��8�^!b�~:��m-ߦkG�"��D9���6rt��4Hb�t��Q�͐�
jr��F���Q$j��X��G��q�+��Zn�w�� ��y��}����ݿE�`l��[z���Y �;�����м��:7��I��Lva)uЛl�
����鈻��Nj
�֡�:�NaD�	
k�����,	{��5��ڣi��_�YT����C�3������^"d�!�l0ЇV���e�3�g܌�(��Y�;�^Q5����0(	jnZ�V Rn�$�æ�������"���AP>y��W_�� 2�289i���<�����0G����$e�x�]x���j�#���=�4Ÿ��vw?q��T��=�����Cr{�d��Mj��W�HL/��5\s@Ci�)���gw�`��1L�ו�N}?�N�j�À��V��Q��0��̊=�� l�!��;��織YT����i֯�5��gj�Z3�)���?��P?��<�ⶄJy��4��*H�����'Lk�G��3�&�gw�;?"�-�S�!�m�p�S��#hbu�*E-ʛ0̶�|f�-�,0�sڴ���v�F.�A��H�4��{]��JN�����f�l�q5l�pI �!���=�8:*1�����c��*�O�	J��t�f(��p-Ct�ўe9)�I�,B��~��<��i]
o*Hg��-�U��"�:!<)P���3R�z#���g��������)�/ۚ��c
��d�-�m���yf�]}���~��-�E�
���od�M�WE6F���R�<D���?P�Y03��.
:����O�Q�̶a�F�b�AL�R)%nԣ��8h�����3�3������ˑ`���0���m&�7�)<�-?ۖgU�@w���g��X�e_�P�/f������vل+i�ikÆ�6V����1�����.��´/����跥��nuΓ1�y��&�Aa3�o@�c�K�a ��{�3iT>��G�����h���^�q�=^�jXk1B�9�c ���ƃ0�LlRg&C�E-@��y��["dX�R��}�8mj�	O�b-gPQ�]���!�d�
��r���1���0���E��묘:�Cğ��h���}V��d�>�Pt>ly¦p�={*���TP��P�JU=�sj�\�|Gh\�d��Iif�P�iIQJ��4����FW���r%�����YTv�mT	!iN$�m�I$�a��c�|�nC�#i�����HM$��/�
[~	}�Y�Q[a+Gz�^�e���;���0�>��6�[PX*��C$�n�alDA�0A�6��d��#A!J;��%;G#j��5�����p�@�mp9%G�'`�,T_�x�Q���E��l�#cA#���zI~���g�ڂ�?x�AN�x�x�	���!9�F����d��rԉ��(�50����I��������s�)uEx�u�)
V��^搩�js?9t{��)��*	C\������ �G����>��)e���Z&B��������c�
�N�億�/��E ��`�'� |N�*jV@�Ww�璧t��(�GL'���+*i��6A�S��*��Ghr��䅬s�«�G̼�	�iO�7'���m8j��4�̗�E������e�F�F�r!�9=�Fi��T�x.���M������j�a�5�X�X��ԩN'rs{�Ҷ��ش���zӎaP10�K ��[;����� ^�d�V�{2�����v��*���� ��<2	=�HG����Cϑ˳�u�`�<z0�ǰl�.�I�ܾ�J�P�Y�������nAiF��\^X���P׿n�@��땧m*�k=�J�,l�r���#�������U���ƾ>�J��s���SsU1��AO����)��E��q�´�b��H0�L#im�O����/gK �k#��p����Ҧs�+͇ͼ�l3�W�zY��L[�sI�~~�^��p��_�����Cbr�W?�(������5�����L�B2V#��c]�}c����%�@����}H�)acȢ�����,O:\Up3�l���?u-�Uz1h�4�rWY���x)��0*6v����H��۹�]������o�i����)l��t%+�j���-*�5���[ۅ~�Lr�(��Y|-C� U�Ȉ�����ho_��M�'a�3�"ӂ{�//�!���1n���i�=kz�	��?�XK�O��	U�򔋟��!91곖O�E$�s�Om�D����v��ħj�џy���7A�w+ǒ�J��LF�9a��9x�I���'��H�çy襙0�rg-H�� "����y׺(ϖjgJ�2��YT�f��U�fB����A��Rz[y��)ţ�p6��9ٍv��ڑI�Dh,���Z{?K�"��s+9�l�bD$3�ّ�uq�7�ty�5����ŉ]�,C��v��7E[
(Z&����7�w_bI�09��>%=.?̙T~<�緛`l?ee��K
��D����o�����nï��_Ο���n�z�
s����~�F�T7�#�P"ɾ�������4���Ҡ��l�`+P�z%5�,�!;��t>�v�]ٿ���`+�����Ȥ}C`7y��4&�~�IHE��C x�!H�����/
t\b�ʾRP<��׳���ɍa�\ )�|��.��B�UM@pC"+�F��4$U�c�hfۺ�1�w+\�ty\�״a&݊���(�����0.fIE���[ᐂ��Z��6�)d�"�ٹT��A8BF�������D��2E���Ls���l�!��``���������l����\-�����(�AsN?��IE���ym@+�!/Q��B����2[�w��ϯ�=�PW����Ǎ\�(���*���FJ�� u)/�>G�A�m�.�e7u��[�޶}c������3|��\4��-<��vI ޶����Crs�_����ۂY��o4Ȕ�q����3����tks�� "YH�rjo唀&�њu�\;���'��u�d������c,Íg�vѐ�s�w@Fx��g����=�����r���¹aO�gl[�ڶ�^e�җ[�u!t�NdA���t`*(��������;����X�s9s���8+_`bL��KrS�,�,-�y�
~d�v1ɶ7����ü ����(�}w�A�j�%Dڛ�N���)'�ϝ��g�E��@v���M%/�5/֡rª�X��>���X���o)��[�B�9�)��q�z9\p�PQ� ���t�D����Ba}X�Aװ|t|p�6d��u]�5��K���u������s;cAo{+���v�v{��:�b
$�@�̙��z/2o16-�{f���:	~q���L��+c�"�h7�?�t�w�#'ͬ4�/�I�B�m��I�f�uۛ���.;��WNV����K���P��5&�`^�ء
~[824��j����D���8z�	����)M���ۮ�7X^E���V;t�eIe��Z�AlWH ��Jf_kD��.a^�Y}Z,��k�5.�����ր��Ȕ��2<O���@[~R�^���}��9{Q
��_����� ���	2�f9q���Z3�'O�{��Z򼢌B���cR���������K[�m�[�S�:^�Kdɤ$�Vľ1?_i,�V3̈Ma9��4��R6�����y3Ǒd����i��
)H#��nN*b��J�d�:b~a��!w8[��V�S�A(BNUk�zW�`690&�����V2�DU���2=�У�#�|�7 �v�&[����w�;h�0�Ւ8{��'a��7��{��H5��M���[*��G���#n�/���~y���x��/cc!/���A��[;�˿󔒔`*j�����.�J���ӻ��9��I5(��	�|���o?\I���Y�^�#,��G��Q�ȼ7�yǪ= ��� AUmo�\Pk�!��ms��2I7�0�-�m��4�0I�l�����\��:į�)�vw(��c��t�<�S(�L��m)�g�5o��k�Z� ^�����98N�c0�������(��Ã��/��nHN���(`(p3[�ǌ��n��ߦ��V#x�<��~��Rȟ�[~�Q�L���Pe�-J~L�w������`8��H�:��>k� ���儜�U��F������I�Þ�&G�,�-�??5O���q�^�NdD��26R�`)�X��y��_.���W�5�:pw��U8Q����~�A��/6���������V&��L|�E������=�b�����1&��Ρ�n����'A���@2�ZP}D�>I6vƾ��G���|`�'��wߥ��ס��*V=E�̾�*jF���1ґ�
���䃹UOC1�vP��� �G�GQ��YC��J&�ÑX�U{�Xg��A�r
Ö)^O�k�$_;ҳ�,Qv�yZ����r�`N�N`�k�"L��z�9Ң�10��<UU �:b
��	I�w\�r�g�
���񼟦�9�۬������6�z({��4�������kJ��R:�����."��0��Y��53:{��0��?k���ڳ�i>h
?���;������ܑƹ�x��>������~�О��A�P:��B���_T��0'������i�M�(���b��{��ebL�*m�8�Eվ��E��dZi��r!�����N�D�`MΗ�2���4}�H�b�����x0�_Z��MV�Z���E�r�`�k��k;�ȕ>��I�����r��;�����sm~0?Bāqb����I���> ��u�p�  .�[30�d9{��s��Dr��%@ڶ���s
R^oa0��Vӟ��e� "�9&���l����)>~��3j���%S[�U���QtS"iY3���Y�`�R������$���n�!�5h��#e�˩�9���T/�f/AbE.�*v��b|��6�n�̏~��]y��Q*�r@��1���*i���b㕺�hQÞp;����h���TkO2��㓷B�É ��髅�'%�(���S�ن��+�+����ə������$�h�Y�
E�	"˨�'k��a�o�t}�z��5�<(��]W��C��{Ѵ����^Y�nШ1��0ȍ[b�ֶ�c����;<�c���4bl�H�����t�e�l������ɼ6�eӀi'��sX�� �r����5�����錪����ی}��p�x��s?w
�Vxf ��i�m�.�t&�����]+���]�щ�]�T1�����k���qM��t��M�L��/5��lBiGd���dR@&ߌ����ج�f����"�-����d�h��4���� �.Ve~�[䴱~j�S�:	�j��%�'S��:V�'�v��X��i�51��@I}WZ8�p5���
~�y��@p�|zQ��D�)�rY�Ֆ3�J=�;G��JQ:?��2�����T�PŁR�¬���+��l�M��U?����Op�-��'�\[��v��z��7?�
uVش�%9R�� (-cӂ?"�K,�R�BX��ˍt��$���襵�_ͮ5#��d�;�/\h�l�����ꀾS��C����Is�M���� �Txn��J>$<b��@��[��`�=Xo��Ӵ�*Aԧ"[]7��
����.أ
0�a�8C�=�lV%�C$t��=�
���K�L�TH�]r�AV$62�>�/x���a����
�X��es�$���<�	�.�$+9ĕ��3�{`~ٻ������ ����J�u�B���U�Ͽ_~�Y���ќ}�`�Ӡ9>�$�=��KX �!2	ᬑú��<<1��8dB3`��M��:3b@s�}}�U%e2�QG���$;�Z�c��A�a�wT�6Z>�'���ReF]��v�}���J���Y��{iۙ�4pǺ�J��::�b�o�H�Q0QLd	�S��|��A�I��r˒�T��(����ʘ���uY�:. � ��G*~�с?3|B������s��x~��a�jJ�kݘn'�b�t'_W����Z���O�Ud����Ao��;�[��l�X��#���r7Br�����W� ��%\��m:H����E�
��9������?�01��+���
���O".��+��7�o��@Л����K;fRV�?�W�1Z3�Y�>oڻ:�B!�?f�fO*h���U�����g`jxfqFo�U$RP}z�Z��P��W^��P�K�Rk�Q&1��mT�T�kQ�x4g<	� 9�F�|O�V�3�s���	SG6� .,����t��
��v>���i;α�UT˼U�
\���`��_6)���s���L�k��9��Qo���?˿�Nl0�0��К���h$-�>��`���|[�A��0MdC�2P�!���[�n�B�{Aͽj3 �k��k��T���ik+*q��i�@�/�Z���u����7`��
���&d��xF��Y���NG��:]�i�vR�q�6���6V���4Yl�$���@�Β��AVV/���P�~�i³���q1.����u�>�Vc�hH�Z��(�|	�T���\�
�[jz���B��}�V/�ѭR}�?	S����H:�C�Y,}�mⳜ��"�	�
j0V��w�����Q��7�m���*L�pC��*xVJ*�wK�F�d��k�����b�{�)���n �υ�䬮֓��k_�	�����_V0��M%��p�{S���R蹖�,��>��HJ�,b|�V��Uwg������0�G9Ż�������+�V�k}�R�7��8��D����H��]�7=<|.��¹x���R��qn��R���BB�s�+{c���iH�v�4R.q&&\���f�B\J��߳���?�\Ʌʰ�ot#�H�eK�wZB�JlQރ���aU픭x�[~^��0��|@`а}���\���Bz�XM�}M��!���n�!N��n&�@�p=>o�F�3�����]Q���r����4^)�a�x�
�!��[�t�߀5R������(��X筭hr>�_�=M�k��Q��t�%�1�Y���(H�(���AL8���H�q���h�p��.Ի�0��]H�⓶����֡�NfE�]iCe>НN��A����˄�D������9� 92?���N���nt�K�ǎ��5���d2?sf������2m�ӿ\�h�{Q6�k����6h*E��<]���~l0e��<�~>0�Q��FYõ�%�[]�W��o�*'��z�Y�I	����]^���"!����,������" ��;���%�V"�q� I
�D����N�(LV��E�C�Ϧ��Hg��|�]���������G#h�����J�M���4�j�7S�jU��v� i��l!Za/c��C�y�Q�p��� �����U�\<�0�S��;��UӬ|R$�wB��n.ê�:�r&����l��˘��6X�b�[�R��S�A�v�a�U�_�bz��L^�O*�p���QuS՟��#��,�5����	��57�C���A7�'��,|W���"�#��	ƣ�&e�<�ݛ��x�L�����~��A����@���B�m9������	**oQ���?Q,�a���#��,��֡�����N�����r<����S��32�խ0�P���5�I�i�6��ƫ� =*�o���!�9�v�I�$�(Ҷ�SR���O�p"��f�/�V7M���M�}󂴨�a�֡�X�@������~����
gT3>Q˭��_��'"=�\r�� �)���X$*j��V�)��&9zq��֬��v�dЛ�uUj�+P��]Q��g��@�"l��Nbˆ��O�o(�׈\�:u��Z_��VW��D��Pb)��j0I5Hު,vه@Bj'�'�YH��~h�P��8�,A����|h^��%�%� ϟ	�N�5j�p"����w�b���8��D$^�!Qpѓ�s��mU!)0	 Ee
�ƪ��ɯ�t��X�K���jj�H ���@e������I|W�X�}�ZN"�.��(�+��9�[t]G���S���2�W���%Q2�F	��3*�,�iX�mS=��$�H����V��lqJ��,�+����a�Xdu����D�Y/@]
Gn�q������J��:_~��Đr����-�7c}��@`�����K���	��9��C���=V�]�k����GyF��n ��֐	U������@�Yۓ|��U�l���9������B��!2�x&�|�D�J���L�8�q2׷z|��Š+9����s P71�U��Iר�S�,�p�dA�#��a��V�/��H3�_���?ŧF:��Ν�vDp��yEk��E�����@M�P�ժ�/��i~y!n���\�pR���T��B�q�,��
go%��hh8�v�zc�սN
$'er�گ�����b��QY�̙\�g62�G���p�T�i�i]�@��5%kM0CD�Y���*��y��!�WT�]de��hE��]��<Lc��r�PC+5�M-}�9�IK�4���p?c�) ٱ�ҜP+�f:n�1e�QWУL�I�̙@g�[ \�GY-�l���,p
c:�g��@��-�K��Х
��k=���U�o�f��f�iO�A���� .��Zg��ܼ�#����L_�w�O�&zְ�pW�W�:�Yx��yz$h�ڵ�9"����@�����נ��-���'j5��hCt����G��C�f�W#d͈��R����M�5�ztR��/�f�A�Rם���#��
V������U�'{5�.hȝ�%�v%�o����[�@8��Ͻp~�p�ҷWz���bw�8p-=����3�8�f��?v�R�c��\����[�
��6O)E΂7���f�;���.E�oyH�E����|`�U��=�.�@���i&Bx��ۀ�G�kRe�����d���.��i�zN妬 �f~�M?+z��3�1S��%�M[�YY�C_0�M9Q�~ʷ���]�eZ�/j��꓏y�mB��m����� �r�E%`�xK����,���S��P 4r����g���S
V=~Kg�������j:�;Ha�Z�+���_3J~dʏƑ���<��\�AS��pA(fƲg��=����s�6�Ɋ�m�/s��U=bRz}�t��`� �K��V �;\�U<��y���EC�f�)1��L?Q*i����:��r�F��!m���Ճ���Sm�,���V���8�Z��~��L�_����|�R����B�zq6yO�~�Mk/��iL��E�h6<�J����nXֆ���%=1���!�6�A�U��Um�3��K�#�.�	�$`7X
�H��悙-�W|�^B��'2\�rRKF��3T7�+���� aH� +���V��@�n�����7q����6��� �a��>9���,�ڈ#�Cm�A7��+��Eq��y�%#}Ö�6�[d���vVFPg #��#���ct���z��J�L��`��s���*\#�n9��7�����І�p��Iȯ%�
X9����`./�Oݞ���<F��@��G8Q��y��7��RN2hP ��1s��K�S@����@Ҕ��!bt�h�$�Y�� ��t)���M=�s��g�nM�T�Ա-����A�_��ՑJ]C�Ԥ�Q� dd튞�g<�֕24:��&��ݍ�����
�	���9�g�Yq�|]�x�Y���/�jP��L=�E�^��m�2]�-�C�h���u�wd�D/�!�� w?��W�.��k�&.��vb^��Fw��f���	T���H�.[nՠSO3D*$Vi��z;M�L�PP�ֳO�g�~��D�/�e��>���i����cu��K|�w��T{�M�w1�r�f�ʬ3�J]��H?��O!"Y�p�w�v�嘜�Sdt�b�Tp��v���X ���<�J�@����E�&>|��	�	��C��Vuvi�s�Ƙ�Z�y??
��7�)�����So6	�y����e�.O�3䭌�e���qf�އ��
��[aK!^�WR/[kt�� ���:�q}3��`��:c	!����	����C�T�>��"N�W�YZA�'<ǵ"�`�J1�H1sbc�=P�!UK<��<p�W$��������۽=kJ��/0>�.��_>I\�؞q
�e=9;*��)?&{k&in�t���g;�*\�g�ي���DzQ�����f�qٸ;���*r(	�n���ڑM�.	M��Jf0I�ԓ]x��L�7-2NF:��'�O���I���d1�ɑ��-���mH�=i+,����OԳ���&�HGTe�۫�������[7�Dˢ���p}!����qjc��h;g-��xc*O�N%���4�H�Xnf>����?ꣾMn��0���8(�r�=n�"yg������4�\��^<ȶ`�������)?�,��u�Y$��F��@s)�&��DW;�f�=b���U\M<��̿������%�b�wt��'2L��7)�A9c��	\='�zLNOg�T����k�q��&��V�0������}E����")�Յ�EO��9�w�6cɁ�H�$�������>��Y�RL���O]D���&&A�H�6� �j�c��J�����I2B?a=�/'�%�UB��ILÔ�5̉3�3v}r��(��9�9jf�;��S悎{��@�b�	�s^����4Xc(�a���p�Ǫ҄���?��hƈ�ƻ��QI��:臇���^I�iQ��$TPC�Q?�Op]6B��gO-R�=t���N��`Z1� :�9fO�u&K{�%r�4
7޲�%X�����'T���k����~�Mb���0W��hQ9e�438��ȸm�IQ�T:����s�������P��[ky�����D�+��y��V‘��$�S�xFL��~X�ŵ�c�,��ͻ�4&�Ub�`�X���d7_:�2>m�S�n��$贻?�l��	���2oa�Q�@U�v���'$��54d3�\JNrTn]5�?y@��z�h�B-�2�U�	ADq#�ğN��E(3.-���V��Wu�����b�R��ŕ��]"�h�� |ڽ>5ރ�}���+����O���Gq�xڍ6���0�Q2*k�\]���7�7�����-�B��81����'(���u3 .�T�����l��0�5e�+��dKޗ��r�I*�����L!�����z�<633�ޔ��T������*ɾ���mW�a����<�a�:�r�|�PX�G���]�p��<�v��u:�����4ޛ�ͦ��n��v�[\�/��ȓu�5[�E�?����`WI�^�x*�7f���w���^�g�������L��Z��m���R:��G؉_�9��a4)U�"L��B"X�qL���D�%שX�Q��E��3Yp>�W�ZJQ�K�)+?w�6�U%0ݘ���d� k��_�;�h���/Q�X�	sc�:Mx��ö�?DUI�������o�K*�F=
FR��_�P+�R�s�d1��~�tH���>uW4�;9ӌ`4
�fӦ���1em'���7Q��(�fQ�"?눹9�I4�ju�@E߉�a��]�|�� {�}�w!}?��}��>mpŭ� ι+��������e&Kb4���r� ��D�)o:��F��c��uY#d��9%�b�"����_o�\�.�I�H���4��u��m��M'�m���%L�\0Y5��e��;��6��,���<�A�5U������f`�&�(�3��g=���^�!�mK ~�{��H�P�BǶ�U�߶zh�����0��qO�N�[���)�� �Ci�Q�H�0�.7ۍ�-pq�/�)b�mY(�I������;��:�B�rx�_�s����[�>9���X����9�v!�����
/�Cs���.^���ƾ�/��e%Nv+'35��䟏�17����'�Gb�;E��ʥ��
��
4�$���sXS��^���de)Ȝ�) ��{�d$�����������d�r0��o	��p��o����~�+W�=S���8%Cb'-�l���C�Ux7q�u�H�cݳ!�>�!�_L �	N���~fQ3�6R4���;����z7����@
ө���q�CW�5\�h� c�7Bw��/��T�̯^rDI�Oq� ����꺳���,�������R%�VI����#�|�D)�]Zo�u�=�$s���ڏ����L��m}|\�[ 6,L��Ͼ��
���@m<5u,y�F0���@�9�hA�������/0�m�<�������#��#� ,����Ȫ^ĭ�|Mv��@#;1:�pdg-�s��;�(1�I��-@����co�)ru���w̹���ĺ�4R�,���~��n~����5�!����G����zL ���䥷�W�M�k)8`�p,�إ�����t��w�4��C�o
9e�;R�1Y3��/JS!�$Eo�R�;3V���k׾q���p�/��믞a��/�/�˒5#(&%Y'��t�jmH�I�{��eщ��8�V����\���
T��qŇ[*T�.�������_죐5k�u�u/6f:/,�م�z)�0��®4	��n��#�Z��^mӃK	N�dV��.�@A���iY�	0b��@�����S�ܜ\�o�*��@�A(6����@Č~�sy�f)%F�xش�M*T�{=�2-l��*%y��]&�-��7z@
�pL)2�Z.����<ʺ%��H��J��C��>��r��i���C�`�hJ��G>Y���#�G���N�f�J� �� ��Kl��*��X��PB�(އ	�p�Eo������J���e�Vd$�`�X��ʎ8��}Kf�����c���O��h�����5��n�� *�tuA3a���˻�ˌ�u]�x��X<�Ӑ�s�&*�U�׋%��
�#�?�j�6��ۑ���aG�UA3�0�M�+q�)%��z�cW�x�pȯ���i��}APO4"&�^�d�l!������~��O�W+�����|�G9��M��)�ބ��� {�]N���i3���'G��S'Xį�(���;L�\tGE�
�j��p�XاM��]*��������|`��V��6�Ѻ�8�"���"��G�'B�2C��q�=9hB]�M�\�HS/�����<������X���DyЯ�M�t���G�z�zl-�B��}{iW���^@�9�#���E����0�Wڻ{��#�q\��=�c�65�tˁ�@㾔�]kMkOwO� �QZ%�j�(nw��Nb��_w�]7�,���<� �`6���Tx�܆��UL��g��$䪜ce�6
��K�ջۂ~>b�S�%_�ʟ/<��m��l�a��V95f�����_�����=S ��.��ў�+�Ma_^��oS�.8��<�~������q
W�r��8�h4$пk8	/���fe�@}x�׿�ߌ0���j�"����)��(g�r��	��{}��H�U���;y��0�x����:O��MQ
�~-"�X�4��i�Yz�M+�z#٧�LO7Fܢ��=��H��=P���٨����F���(`Y��\�f1֭��vP�����e��L�'�媜��"�T�'>D�oEb41@��E��/V��^�G8��Z���4�Y0��ࢗ����ԃp ��� ��[��7Z��$�޶��$�ye�I�qm[i�yY��ʈ�:�CR�����uj*��<��k��{6',��͌�㇀�S������bԗ��[�koS�T��5OG�ѝ�Z�S�T�S��zy�6%b��VY�#�1<	A��捡�1w .7��f�=1� �0���q�c����y�nƸ�aܾ0ap�eS1�Z�mL���6��1_a&+%?���Zz%s-
�ͧb�K�U8����	�{�v���/���=)�zp�w�}IBk�$I�tZ�sllc�Źŧ��H���iT�>��yWϱ~^8��F!v(eBWX�T�*
#�b3IQ�(tۺA$�R��*X��i怣�?��Q����)H8O/���`�!�ZI	��H���{q�������+�\%�i�T�"�<=�yD��h0�%�x.
="ޑG��1���&�~;�z<����e�z��2�ƕ�	�
�n=��W67K�ܑ�d����� 8MH�-A��M�z��@�B"����� ̆�u����5��D�7W�z�#W�G�. &��!�T.s`x��[N�j+��7W/,|i[(E�+��2��L �<�{?�[X
IQ�.S�Ԁ���d8$%��ZT�^���C�`�_)f�K��-�+���K��hM�.�j�~��I�*~j<8r]�����)%����%��G������ȪﻯՌ�P&�&o��N�R�'�A
�>���͜RP�l�vkى�X�LGz�[>h�6�Ty{��p�W�e�g��R����`������)��'�rHR�E~����X"2,gp�8y��O���	ny�ܽ���,>l��gTMv�1���`)�?L�lB\�+�`��������Q#�4"�8+��f
񇀷b�9����Ӣ�\	o�2�D/��Єu��'��HW�� x���i	���e�+�z�Z�>;<��4�\��Mػ7�p�����P�#�%2��q����V�ٮ8f����u��J�@4γ�Er��/�lf�Ur)V�Q��$nؿ�1���H�(��Aì���������ef���>�����nI�1:��O����Rqi�<$�xz��31rAY�F�����/bUnwZ�;��xO��x����꼱���y\{v2֛W3��0����|34��1|
P�,M�]��$��E]��xic�+��I���n_@K%l�9�b�Ku����]��y?$��ŵ�0�9�q�	�E��W�~���QL��kT�Z 8�a���g`�=G����ە��Н�b����W�eIK�/�d�˶'.[e�E	}AbX�6�V�- �2`}K5f�Ƃ�U��hu��_A����8iҋ�yOE�ɍ� ��%+^�Fk�Uf�u< �6��¯ǟ�����@u�r����1P�A_��*��
�]�@�bڍm���*ǐy�g�:Ü����!�Lw��O�:���_c�ܠ��3�u��.j8��y���^Q��vS��U���%#�8��kО�[R���S�]��,�ll���8>x<R˼�����`�O)7{t}\vMݻ��!�<k$s����*cd2����dr(U9n�.2�	8��b�D�W�_LNg�'Q����C�A������J��'dl�~���ͤ���<IX�u�Y�aa�;��;k��fAK��Jf���J<�uYL�OO��p�̐`m:�VC[^i��ZYV�Bt/��<����ص���c��J&�=r�.��^k9������8�3ٍu2W$��,|�-nF�#s�����x���k%�%�4t���3��m�<�Q\Re�'�u���%��tJ6��f>����"� GX���� �e��:"K�dDJ�/��$5h_�Q���<��w��x��
�붳����_󇩚��͜�q�`�X�1����k��Y��h��g̅�xg-a+�=�_㪾��S5Ȫa��"���
X�<�X��̣#fKv"(.tj����{P�MY�v�&C$e��=`8�lLiL5��U����>�G�9�,ؠtG��Mt���ӂ�K��A��)OwRŹ=  �X�ZUl)J�ꢄ.����Ō#;*��,5��\;�=��|i�![�n��lҵ��5T��[7n=W��9��-�:��� �0�i�ZK�����7)��mb��R7�?<ͭ@�i(�N��fK����1���4��o��0�p5@/��ۿ���kU]�`� o��aI��<�df(�[���=@��]Tf#l��)��g�Z����5�qE�T�i�݁��6ђ�����!��y�+�ć�^�jǈ�fb�Ҳ@���C-o�}��SQ\.~XP�ph"�^c�U���i��O�[�*i���l0�-�c�`y�0udA���s�\�a����a4*��|��?<��n^��Z;�F �W���&c%��,����`Yߓ>�lչ������e�Py>�x���,��:���pD�`U����,��W��������[O����,D�����x�>�T�����:%�?���V۳�
�z�\9�Z��}z��iݟ4�Y��k?�B���UIf���x����0*���E�>K|:���-B\��u*n}I�`	8�>�0?����{r`��L��Q<e�E��(\��Gݤ���⦑���w[���f�����M}Dי�!�q�����I��W{�˛��)Cw��������Vs�LŨ���ꩤ-�SΣw0��FQ��A���Ѷv�:3}�=ޱ9!.�*w���${��rv�{j�@廩�����V�UWp���L�_3�m�}���}/�#r�3۸F]sаnݡE&CU�ԪІ�pclU;�p�
�� �?	8�A5bة����;1���J3�9ʖb� �U��R!v�d��7��v�c��ܕUr���m%~���SsW����,\�N
����|���̞�����(×X�e�c�j��x���d���=�Eץ4l�REL�&j���\^<R��ŀ��:H$3��·�Wɱ&l`�!N�K*Ii�E-X������L��́`�A��
��Qk��2�t���7�v,X�|��B8�'���Ȅ\J����	m���uW��)�ߠW��Q6��[D��?����UT�q볈`;���)�v14�H�vh�E�'4��cp�ҧ�g���\|���x�W ����J�o���;uk~�y�AI�����	�H��Mj�L��2`F����D�����3හ����[$ә��W`)�+w%=�� ��\s5�(9*o4�q�M�S����s��y�"�n����S��?U����ɽ�9WxEs>{��}�4��a�lH�v�WЍ�EN ��H|��L�3�'��D�,�E�K[<A�0�qꪰ`�i��hז�y)X,��dH��n�L7�d���*��sǅy�!���ToIqL#K�n@(����������AL���՛�����M�8�%;�^33�.W����x	�	.Ρ�e�{�����i�iֻӕɟ$��e՘�<B6}�l�t�)�D���	�F���r}�z�&�´c���K���	��弤-ۄ���������X����o���C7��4Y��ʢlڠ�q����I��_�`��zs&}�:�f��7�F	��3��*
Ffbv���LPYk.˕W�;�"�rL�*������A;^�c�,���)�R�z}xi�w��"� ���������|���t�ފ��rx�-�F(�к��	&�7A.0&��X�mO��p��:��E��y�d3D��^�`�!{������v�P�����k�:eL�=1gj\��7�� I�&?�bL=�k;��@���Pμ�� U��;�);�V��[���A�y,�B�D�C!<��`�Y��f�T���*��s���3���?zb�iG�߭ $�0sUs*(�� ƄpMG]��3���mhb'��oy�,��Z�̔)S�{9����F�o�-�t�ʃrj�9�]"�Iuҿ}�-��η�l���Ø��?5���%�+^�98O�)nb�şVu�����^8�ID��`�Ŭc�$��Z�_r?���$p�����|&={�~���g��
yh'�t.�\��4�-l���(�����x�|I c�=A.�6,xJ�)�Q�3�[):_1��ch�l�b�b��!�dv+U���x��u��1`�e �N8�~��\�]��1a��Т���{�[���,G���e)�,?J�!��vy=�F�h�N! ��~@���S��QO�����cu_fFw�m�^j�/=��j[��[�\L�FMނSk�Z�in#������ǀ��:�0��8������C�ڛ+[�l�S�o�xv�ר�@��g �b�7���z�OzI�[O�?�tݐ��=o�{�ۉ$��.
&��X*�	�sF�3lkq��^�l-�OV3����_�@%��$ST�8;lZ|2V�)��L1&����j�ž��t��0vk���L�CA#`��RQޝ:�o��������RHj�@�#���n�V�I\��U�a���04?���Ⴅ��Q*S,����:��6�)��(	�� ��㉃�aX���v_��wnBl��[��P�����Ȑ~���P[�����b�1Hk,>�?��!�NCj�c�`���fZ�ڰ�_w�.L�/;�C����d.YW�C�W�����E�B%��~�mO<�|�7 ����(�4��L���?���u���H����l�ja��$f�V�%5��`�m�`B�t���t!/��l�3
���i��(@�u�E�w���1�h��yd��}]�>��W�-�����VOe�M�_�l�JⳃӞ�����m~Q��g�Ĵ����n�Җ���a�'ӫ9	p���e�����In�d��s�`y�ZPH�Q�.%>��$Uh��?��qc��p�Z��H;Bw�Z�4,TIς!#�p�uNQIU$�<�pw~z���,㊋��h&� �̎�k9��Et����YUg�������Ҽ`�?�3����^��T-rw6��ֳ�ֿN�mR��]	�I紑��(����w�Oe� ܔ~|A��%���s�\s�k��W%\2Kń8��=�zB��Jћ�_�����ԋ��&�%5����R��_Z�&+��J�A��"�dO[�Ӧ�US:f�qp��`C�G����hf3��nt���v�'��SR��0���F��/���i�q�Z���fz�M����M�������z��z�y���|�H��O	��b���G��#.:����뢐��}��=J~#7��?̡��s<Z���L��b�)�a	F�� S�M��%�|�FkSo�tr�6�4�!&��g��l��FD���_���V��&9�]Q��_��+�҈8*�|l���<	?H�x���n	q>�Cf���<K-�(����E!7U�7o�g���9��[e4ҜZ�Ɗ4�So����u�B�����ʝMp��M/e�>���T�����Mt� *Y�(��鷧'�iD#ȋ�ŭ���F�G래^,ą~/SIy��he� q��s��(��]�����|�k��0_Go�t�B��`��D�t���"���#��x$_ػ�j�,wC<)Ҵ�ap��k�Z�0NU*d�5�\��	��D��hmۉ�߬�b0i��*��`6%�
�8��)�-�(��K��
5P���YPM��KL-��J(�B����(I����g�����}�W{���)B`�zb�G ���V�q�H�����0N�)�k
��Ԟm�r}���eS�U�+�>)�,�?&�1���)=C[�%R��S¼?g��x����;�C���%q6��~��BT0*�	_i.-��|ũkT�$�o��ȵ�,Qr�%�S����`��]�ƒNrِ��]�o���V��͊E�0e�S�P\h�M�h?!>Md"���o�2���l�R�Ũ�{�d����A�����Q��%i���~���F�w����E6��u�dC�ܖ0��Y�ݓl�N��G�L��C"�bLN?ɹ�\4�k|O� 2+��ɖ��MM���ɦ��/�'��
Í�P�o�!����b}92�2������}�q��I���ݭ��96���p�x��Hs%:���a�d�s���GN�e���C٭�վ��_+E��2�����ݤ��ԣ4f�����w"��'ƛ�	�Z��KS�+G��
a�=RĤ��t�a}l�aB�(�{Ǽ�!��;�����Bo�ֻ�4����[P�	租������,�mFWg�B¨��_y1Jp���ִ=#ʋ�O���X��GJ�~mUx��"�W���P�����׳�UΪ�E|�p|�oi�}7�Q�٢ adyw����G��b�V.��9��x�H&]|<>�lZ���\��P'�����a[�|���!�Q��p���t�����h=6i��u⊺~�����5.i9e��$�EP�����*��c�|��j&m�x�lkɷ!h���e���h�Ӝ�f��^G��5��'����S������Aþ��U���dqgcj��O�I���)i��x3n�-p+G��;N̴f.��ٮ��Zsq L=��]��{��ޙ/��ַ�+`T:c����d����t�o/�.�[aw�G�x��z�g�nMB�2�w�:X#�	��V QG�q�{���2�m��t���M*���rA��������`�ƏpZ��H���=�ޢ��O�7�M��խxlh�D�]�����Ҙ���k����fw��Xgf�a~r~&3�C2�|�M���/>�xj~��"}MȤ)iOeo�}�x�ed�w�Cq�ߺYTe�7���]��ӓ�
�����Ί��H��}�����Ř��r�M)YѭkhâEe���[Rn��~~�1Wa�aA���t��E�̱��l2��5"*�8~H2�����ra5USy�mf�v�ٚy_��"
�ᢁ��
�d(E!�g��&��Y�Q[��\��$�/=�T-���Ǜ��mh��G��uS�)�yk+���X�'�MuqM?_
���]h#wp�4:����15�d��Lz��P4���(����� ���{���������4����1�Af<�m���@���/�\lrf�8��U+=JP��/N�fm9� ��ݒ�V�l�F��?���۷�s����K9b�!��#��+q/<L�ڑ��v��%�o�<R��ޒ�	N����%�ID	�`�k6W0�EH�? �	�����4���8��]'�=tI�6�~B��p����f|���㕻�ȠҦ�Fm��^��"/�@�����T�)��ā�#h����=������?���*�4�M���]aǾ���@rm�K\�z���\�æJ �k�b�y?_�b��'j��5�o�d'� �/5����1�v^�=����{i�#(s0�P�p
z����,)��t��2X܎|�2��~�9{D���2�׺��U�`8�_+Ĕ�����k��"�#>(K2���B/�E���7��l'fO�/c��($:���7���o�r���rHa�:hB)�h�ge/y��|�.��]I���T����o�
�+piX9�ˮpɊн���G��� �l�g�K:gDLxC����'B?�>V����s��e�R"����Y*e��G�d�h9JuCf,@6gk_o5\X��������6����D��SL\��aWٯ���,F}�y�`��<�� !��)�
㘨�ܪj)([b�F-����j��6��â-S�K�w���%��]���4�a������b8;�b��Y!,�wu��y�{�M��̦��
�4�����+��b�b��3a;v+ި�R�X#���%�p��,�S�k5n:h��5IF� ��tV�e-���S}c�V�9ѬwH�?DI�FFk�L�<�lw*my��3z}5�Gݜ�!`#�$k ���ai�qK��TZ��E��#=�O�v�|�!���G�-!��Fd���FKլ���X��h��N���X�Ӗ����ӟ�LK�-=<��3�\�!���H�!�xs�	#�Ԝ�s(�bJܼ[H�)�e�Db͓.*[�kwnI�~Y��>�R�lۃF��&�`�a�+��d��T8P�v�S�y\�|#%c�pa�n^h�9
@&�7~B����uN�������G�BϤu�Cz���&�����,K���1a�?�ck��~w�$քч, �-�(e�U��P ʴ���'劀���nt	��	�F5T�T��xG̳��"��C^�謘vt�� /�$i˛�ye��O�FG�����4~�\J���`�4�g�u|��b��$�ٺ�D�64��uf�)̯��p��̵���d~�Կo3ܳ�~�Uڃ�♈�Ze�N�pF��)���h��w﹌֜S�)��Vh��j�: ��GE�&W���%�f{�c���-�0ꪇ���|���(u��_��Q�M��Fz�iPh�]����yH8����/kaD.��ocN��U�B�Nr+��o/�ҺL+�niʕpC%�u�ǦM��&
�%���p �X���t�bP��3�7��HR|�y�M�aq%e�p"3V׎�|�`9CH#^�ZBE�쇒ص�<�I�|�Qp�K)�)���\����[(m��[e���Q�iO�Y�{���Z,�y�Ra��TG�������܊}�F�1 ?�A�bU���z�@�`2��&��\f�?}�Ey1|�q�<��o�]Ө�T�Kh��j)�02�9N�����q�2�	僊ώ���<S"��@mW�o�^'��y-[�M�P�����?�B��,��l�킨��Z�{N����ш������?"�)����y�-���@�t�G!�*��q����1a |0����e�1���*9�NAom���Q�J�$T�,*,g@�3m�S�3!���+M�c<���Yւ ��Z�n��n���E��t���`�n����[��X!���rw8�$�}�)�)�0����
#Xg X7�0	������'
�o�p3��������G�����`���j�e�<��N
�$���c�8�>;�;��uY���tƑ8�|
���p�dzY���t�f��ߘ�i0t/�:��b�)�HF���x�/�0ٯW� Nf�K���2�
���'������bm �?}�~��vDe�ET;�9.f�Q��*�)�L�lγ�i�7f���,������|���lG��@q�{�u�_���@>��ǅ<�6{0W6v��0^)D���z��c�$�~Q7�ݚ	)����'���Is�����*��	�W~�����r�?[(�h}���=*
�v�u��`����@�`h�~4��5���}�;�,���{���ѫ����FAk��D@S���h�P!^��
76����(t�ڟRs �%^?�����I3§#�M:�,��혿�c:�@	��]q}�N�5��2|v�ެ~ �X�Ѻ��B�F 2�M2#n�{8-7Ɗr+�v/)��f�&�P�1L\��'�H�
ߥ��zQ<f��C�qU��K#B���^�Q�z}`)�{絛��`�~��K���<OE�Ϫz��?�lK-���������Ǣ��F�ůu1�M-Z�����$��tFM��+~\��HHB�j)P�=3��vn�ҿ/ڿ���*n�(����6e�Β�\��B�l�V��r�U���-��$*YV�nܜ7N�K�y�)��tT�Mӂ	"R�;�BAP�2�T���Lg�����	�lp
�CM��m�����^!6+�� "M�gh��˅�A3�օM�bsz�w�="�8��%m��8�b�0��e�E�ʊi
�1Z��Sܫ@��;͑T�\!���I��jǄ$��U�݆�#��a�jYcF�?�
��a2�&��#+��#O�^�i`��jZ��r�h�{#		�t<�g�eA����?Lz���"��|VE��Gh�[�t����a���E��欠	�ҌB��0��3T	���:��]�7��s"��t�����Wo�82g�؏zrye�*���8�����v�Y+�d�q"w�>�Sf��#5����un���VB뻡�EߍЏ�)�"��1�����w�p��%�E��&?[�d�h��V�I�b��wk~擉b���n�h��;�!���B%$=�����e䛬]�E/V�CKj���u%]E��R�v~X';9_׏��}��AI;o6"�IUt\�7V��h	�pfD�A�EGR�h���3��1Ę?����Wx�=^�1[����q�&0�����^����6��[��+}R�\��Y�1��@����	�:גN?6�h���W.1"�.t2fM1vO�XͲ�H�la��b4��=/�TM���g��>�䑵�o��	����=��/��T6,AEl$���xԉ�Vu�_�/b�)0�3`�Sh~�����H���D3�ǿf ]�EOt��l�w�mY�%�s���٦|%B��#���d�:��$|8E��(m���J�W�J9�4���P�<zZiRG�������Q�H���ۮ��~���X6d��43DM���g+&������O�	飮�Ё��a�9�9�x���^e!U�P�Ȣ� E�o�r�]��Q�Z!fr��$�/ɵUc��Z�X�Ə�?���ҹ��.�:��L��3��4�JSD���1�JBO�P��4 ��\���b́��tI H�i���b#�Z��`��A��rr�z�_�^¦�`4�e���$Xɧ�(�0{���#����Z����%��n�i�sn�r�pdқv����*Em*5n)�����~�؂�n��$��αSA:�L�n�>|4�\(6��+p�!�ьeF"��i��Zw��j���ʷ�����5P���K��t�?�N�I��5�vJ����*L�v�p^A���(^#yD�]��8�h��&�v�v̤���w^������v�MUTxhy�	���N���o�R�l�@0KNk��o�J��¢�2��A=�p�h3"������]�3��@r��v�u�B;,t�=�}�����A�˕yw1^O���{�O�� _�ImZbX�4�y�.��[H������b�O����@�рa�[kƝ��Q��N��]��t������#�:�ʨ[.�;�y0�HT�t�lT���#>Ѻ7��&�8һ>:&��|
ȩ<���/i@���x Yf?�QC>I��ޝ�Pg�P@I��q�anI�Q.?��g>�yj�v!����^n�¾�́k咾���u;J���Nk�C'�~8�6��&*A��Ry%!i�����ȟ�����[�Iɝ�*+
�C���D�Gbr��U+�f�R���z�U�g
�_���P%`mM�0�0�K�����U���;HZ��Et'�_£�N'z"��`FS����*�
B���͆���քmpa��UN�8��)袉�m��/YѣڄF?��n��y�~�SJ�
�ܲ��Z̯Xj�-�tJ�R
zY���"}�:
��!⣥yU�X:����j�����3"�Q�7;�E��{Dm�Au��|������#�qOϣ���2= ���R�D	����h���H����A�	p쭠N%��������`}������>8�r�c���V����D�9w]����S�� ^�MGQ�	B@�EA=�o-;�؇K���O\MH��^�{eb�e�܆M2P�Ǚ�e-NzH\���7f���*	�m��Lp[��x|��G6�52�oH탪��f��^}ן����%��8'�$F�]�g,/4�&�4�&�bY~o���؃x2��z��7�|3�|^��UQ��C���|Æ~Oc*�BV�h��'ڸ��!ʊ��Q8Bl�ZT���8w;��� �����cߕ��$�74��b%�N��䞸��s�
r����=�RÇ��Mư͕>�"�]vO ���V����r�zovU{���Va��s|��?���ܒ �wc�\ft��\�bP�7�oCKRbQ�����b��*��,���	f�*�ָʓS�8jO�=�F��Ti�Z�çN���<U�B�#ͨ�
O��Ai�+Au���9�tb-w����D���C^8��*�7ƘvCh���-��𧁶�dGt�ZK= *�߻�,�^��u2����e�j���/����ʞ�Pv���	�T���$�xX��e;��� H�[�y���c %Yܰ��ʹ��o�ݮ8)_<�Q�&+LW^�'��x�s��$�g���rx��V�b�2ݖ���3����e�oG��L��J�;�`I*�k��CP���ȯ�QDQaf��⯩d<�0܇ٍV�R�+�*�Nh�q]a��cB���i�cg�#Q��9��2څ�Fj�z��E�l��@���R3�8p��(�Q+6�<u�R�a����{��Vє�C��*@pѸ������6cݕ7Tz��UR=�	��,���8�l>�~��/��#�@�T�eZoT��(�����}�: .������ 5�����^f�<��䚚E	���5�����Noi�D����nm�
'��M��׀A&�JAY���b";֞�����1P5�����E�9J+�C��2,q�~Uش8V$�ٯ���]�&N)~��X��J�����IH�:n��]35�Z�,X=a�V�f����׋���| 1HS C8���nQ\�4���^kw��£����(�=����O�z�ӠR����0���쑔I)���Z'�Nj�v՟�/��"h]"@���eZ3��WL�	M�#&!�U�id.;�H��m�!�$'��MJi�旬ﵜ��2��B�9;�_}4�cZ���v�^��C�EwY�x�߃�G��}̛'s���ﱉ~���Ƿq���ێ���.�G�R�&��F�j�/Q"nG�ɽV��/3l}�b�1�~�ޑ�]`O�%-h�k�:!�1VݥcVer�2�cofe� =�D}�����RP��J�$�E�*��Q�H�@����j��T�3x���M5H��
ÿ+�.*I^�e9�$`��i\��
�</I�e������]����;�(���: C��ΧU�ٟ�U��m��,��zƯ��oi�#Y�"���ZV5'/j�s�-I!�삶`�����e���ܗ��ŞL�S����nIq�߁h��o�T��<�aH��4��3q�A�� �~��{%\̺Le��~w8{+�l��7P��1fW�rfI9�b}���a���i쫏�";���#Of,����)���8	4O˛�J�g���r���	���j�S�J��f�Z˵s�Uy��4�a֫~20ª;�^0�6��BgM��n[i��	����֢�Lj����B�ݩTW�ך�����<�g�������Rɳ��rO��K�Uu��������oj�����_2�i�a�]7��4u��������/\Bx�n�IE�mE8�;���Vm��'& ��E�v7�ͮT|��� b��t�q7���m$ͫ9no27�0�,K7yG��(��������?���X�����y8N�}�o�8�B�	h���"�vj�8���Duؤ�*�_�F�FG�gt�?��5��a0�m�~g���LaS������M��/�Ӝ %����z�dZ�a"�IO���7���I
������^O���Wٳ�t��ד����k<��k/�ߒ�.�3+[�`91��솄t"*V��D�1z�Ĕ�Q�M[�p�{�"�]�(����<)s)1�\\?��X\�E|0����f9����r�Ae1F�P毂fY�I!��6��T����H0F �Xf��0
�H���֞�	�&{�2�%2O��b �#h�hg�8�(Ei���Z��{k�Y_�����3��1	�=���@�w$q�V&g��Li��XI��#CI��L�,��&�'&[�����m!wȐ���0�}����Z|�@Yh[n������!����� �¶�9�8���cv�Mx���d�����
�ܽp�L�����)�]:�G�z��7&���9�JDWl�7X�'�q�;LL�RRp��/�e���~�o��W3�|���H?�o��Vwٖܿ"�8�qfD��$� ���[+�b,"�y-��6%�*'O�����%Q@+��^-{��fؠ{i޶^X��`����xyO<�7l�X�)�k��ٿ�i@�݆��sʚ##�~h�ϬUI�?+I�F����\\p.�*�|=�
y8a{���r	iC��F�ߔ�}�t�SW|�$q����Yc@}��T�����8f�F�����۴Y��$IP�_"�R�b~h�w�Uϟ4~��)V�
HdW���n]�z�#-޾�:���m/��BV��{V�Q��.Uu6[xo���'aH
�I��U���M��r×����ܨp�`|�\/�E(؆�G\wu��		�N(D^v�Y��`eO��:J����P��܉�Iy[��t�Y���z��OE�}~e��Z�g�/����x��PBn�}f���`q��MvÀ1�Я��Q��@����m~�)#:�@睇�، {M6�p��B�r�b�������W1� n1�� ��mN�4�Rb�	����!�Q��ě��\��������CE0��<	r|�0̺c��Cf�8١���V�-�����k�0/gu�������5���̍��va��sbB��#���~�9��]������9�o#/��ǻ�@���ヺ~�Ӻ:��X"�%YB����K��I$�Q�����fV�/���$�z��h�#�'}b��I�����mN{sQw��U&i�6d�������m�k��eg�b��)S�vqP���V4%�,���)���I� �g &���6^d�a��W�g2F��+`�C��=�l�_YJ��ը�59r���d4z|S���P���ëq:EH�����~����j5N(�Վ�Sht����J.b B�����s8�i��7E��G�~�G}8U�������E���O�q-_^�G~$��Q�l���8�y�5�2�
߾��Q�#&�$����e1���=�E%�iN4A5��CL�qv2HT�8���Ś��%w>OK!
֏-�)M�(��pV;X"����!ѥ�w�k�%�5<�i1�%��M�	��`�?��*���yu�a���ƿr���8ㅿYD����?�/�JB���D��i/{��|"�͍D�4�'b�Sj��5�V��(�x��#)��\�(�GF�}J��'ƹ��jə�v�:�_^��Y�vx���U��ѭ��[8�+ Y��jr��T���WU��ew_4m��=M��qwp'��Pi¯�����=nuE)WGzϔ� �6HG����遬��/_�����h�d�#�v`9旑�hW�X��i=$s)6W�:ZC�qG_3��	�!��D������	@DA+�4)k*sW�s��VVBv�O�����y�L,k.|'f���t�Ol
:5�'�a�m�����g��ʄ�\E�C�c5�m�@I�~/PI1#B�q��%��`�!b��]�s*H>�GU�1�ǄM� �*�:!h����:͍�Tl+w&�L�#����6Iߝ��P�H�k��Q����$!/��>D�R$Xe0_Q�y#IN?����ԯ����ʆ��%�g��m��]�3�d�8��{i[<T�l�`G�$��<�_X��H1^#���MM58v�$="!qkЅ�]+�0:@��Yp��u�M;�i����|Y͕�b�f�xF<w��6�dK�=cD��%)z\��L@�h�[��u�=	�K�W���*��{�T�@Gژ�_Wx���o`JI���=Y�V:�^t�+U�N��%�!�=\l�b<��:�Vu;fSO�25��a-�[זrF�����cC��7C�~\�5�7U�`v}x� v��9���0єR�9v�Ri��:�Y��ʎe�����FZy2��r�" xL�L� r�6q��������J�'�-�8!��]���Xv't}*�"���p�����hl8c2��h�GF�����V�>�%����d�y$,'C���2(���Ԣ�uf�eVJ��Ę�*�g�E���0u�|��'nǕ��QzH�HЛ��B��S����2���'��t�����C�*�OaQ��R?��Hk,��=�z0�?qT��� ?��FW��}w��ém��e�ź�x��i���-��k ���Uu�A4J�5:����(a-c������${n�/:�K���9����R�';шQ�� kR�q����M���_H��'�.Mo))ȣ兘��l�����i="G��e��a�`�����Ya��f�r7�c�����i��U1�mI��<�I�D�'���J &��-��5
��$q��#{�A�{wo	tA�㖈2���a��H����nO�>�zֿ����N���6�k��ηқ�)VI%AnL�%��L�P$YI�{s� �އL�"��=�Sj#�y(h�&�/l�qГ@��,h�4J��[�xa����p���a�j0��0e�tQ ¥$�k�P�C�W>��C����N�J����b���2���U��ʦ+P���K�,9'��;[ޫ��,�!��efv�Τ%D�q�M�:�#
���C�
m���&f2��;GT�U��UzR-�%\؅��¯�T�z�렔���B%A�g�/di�g7O<��N�/,�D��Ds��F���l4�́ɀ��$�,���;����E�yz,%A п(+��$�n�-Խa���%ԁnA��_O���$��+������Ov���#|'��v5x��5y�	c@�9���~�6����
muu��B����BX�&�Ϸ�^�������/�G��{h���F:W��c������B�?0M�Jc�V,�Be��k�v�KY��/�O8*��j����'v�Jp���e��c��~{�`5n��j�&q���oΔ)��pH\� ��G�t���U5�m�$�&G���4��@$���<)��|ftyD��;�hi�R���<ށ�֜���SX1�!�vh���`����A/��'�C�S�SK�|%���41z��Gru)z�A�^�] ft�N�,���1�y���׋/#��w�f���,-7��:r��.��+�r���5|?{
�f�yyuKw��k��� ���D�ؚ�5���'����v����'�}m�w/;��&MM �D�÷,��O�CvW�f��M͂���M5�)SզE�d9Qdg�tN����;�U-1�M�r�g�<ASE~tq��x6h=�W����:�A�s�*VF��W�~]�k���Nlָ�����ԝ��CF�����x���QM��<̟�����ݚ�En��9�ɓ��YJ��U3��J�p�������a�j��X�⧸�Ą���&"Z�9KT��7Zk��G������ �2�AP�N��J��bk{f/�2:��)�y��0�TC� ��X��r��o�L ��=ԫ^q�`tnnp���aH�{�N�,������n���4�F��yV�0�u���K�)�5'�P�GU6N+]��o>v��w��"o��G�.BL^�u���2!b��0z�׾��'�|�={?�.�����w��M����ǡ U�!H��H���bw�mY޸�rm%#er�3�&'k�X�9g8��b��0���Fg�	C�<|	T�w������{V?��O�/hl�!��`��_{��UL�&��S�h�/�#&��$�����^x,���޵ٹ�}�����?@u�;9�q���bڥ11���x�a��B�C��\���z�ǀ�Lq��oC,��C��X_!�$���W":��B�=�hO�){y��{����MKuF�[�YaV�U��[f��P��b�B�,S7[��kT��|Ղ�	7��?N����[|�2+�HP����[����d�f��Hȉ�`��kw�,}c������wY����^�֟Ue=-�#[��MP��#�a���kF��AJ�@�l洜��*��A4F�)����ej5k8�$�e�� �}���[9wp�m��1W�C3�P3d�k\K�5�*5i!t�,�������'y�%Y![��eC�LJh,"50+M�9�����`r��?�ș!F���������,�e�,AJ {(�A����%׋.,9B��S�>crz]��(KE�S(��_�O�����fl��uϥS�8��:���7P����?<�$��l~�\�T"�N+^�f'��L���e����:G�X+l�vy��s�Lo1�,Q���z�
o[54�L6�0=�Si��Ɩ�\m�vFU���$-��zl5+�Z0�g�R{��4?­z���aT5���m~���j��ӡ&.�S�;�Ā�/��.�xUdq��.E�V�-A���n�r�k�������:R4��Z��4��~�R,�%��K@�G�����5��bv.�q頙h(�C](��h��I��Q���5��|l���A)�bT}������8��zё��y��ZmK�"m��ܕO|Ah��xE���2���H��I�����M0L����X�ql�2<�f�zG`[��H�d�e$�}�z��	�"Փ�
�?��L��)Xj����" Y�.d5{�ӏ�lg����C%1�|�����y��MG ӴE���qf_i;Q��W��������לjW����B8��Q���Q6��{ L^8�M;mi���>bx6�w�������q�,ƻI⒓��&:V��ɉ$�V���Ԟ��Tj��(:$ZH����d�wHf͐F�����o\/��rꀲ2Ֆ��J�ϒ�1��	g��L�>/ѵ�{@_�6]_��#����|Xۈ�3��&9���ǔ5�� �(���41��Nbv�4����C�
�%�#H���i��r�y��@�����]A�@P���V��� �^�I�B-(2M�Ph���STSn�5s=�d��e�. HYo�6?i���x:��Q	�s��V$�I�S?�`����oO��P��u�p�����@��B��̆��r�ĚM�;ïj(���7��0%E'΋y���XjH3՚6/�jj�D��Y[�4���^^S6ïa	RjB~���mЭ3b����C��Y��TLVR��=\t��6�!�����u�c�-���4d����lWTp__�C:*h5:f�.�L8�T(���<}������zP�����->�k�6��)#����yz�%q��Fs�֋�i{֚.���Ɣk�(�+�pq�4n��$x+�|�R��ٍ��^�l.�)�������*��p�)UgJJJ���,�+
��D
y����@M��W��f���-�չ�R�
NQ�k�kn�ys^ CE�e�!�1'�E���(Q�K����xfvb���q�;��C �n��R �H"�iH�.����>0UyX�l(�:�!h~���Цa�a�I-�	�nFp|���8
O����N�{�M��Q�	�d�ݞ��fX��YA��趠��`�lْ���i5*�XЯ*�bJt��9��kZ"�6M T��8�ʡ��K
��Us<IrՎXK���%L�\�$�&,�ԥ�$X�+Y����m�=�J��h�E�9�a�03��8--�ӥg��hpI_u>D'�u�3�b0'�c]x;���_�^����i&zC�D�C���&�zT�U��F��w���9꒔��+g���k���^�z�q�|���ݰ$Z�@��gwJ��v��Ҙ���P�>�(��L|� �`���ox/f��BP ����\�g.,T�Z��#�3$�W<�C�b����Cɼ��(1��G%TQ�$��Q��5.u$���T�ҩ'f���Nw;r����d���b��(��t-��x�:�NK�(Pˏ��F'D���)l���ZT'H+i�;�Tꐾk2�F��Ǽv `��{8�0�!}�Bg��-�\�t��������=`1�� �r3�5��k�f��F	�����#�s�Z��� ��dp�-|;Xf�S��/Y�0�*-�e�u΄>*��梴�m��T�{��p��
.��25�{��-�Ԝ粲�7�JOV�ِ���Y�1ѧ�Z�6�OEG@�,p)��c~D�\��,�8�c�T3����yt�Ӥ�za��u�9MQY�2��[mA��~�WL�Zl�'֩?L)�[�K-��QgL3)����xυ#��Ɍ�ל�����(a�fd�c���oa�ż0�yG�U�j��-5S�����L
��^�J�/,!ۿpM�{֊ �^a�:����c�͝��6\�ơ��W�q������,F���n=�Sx�j|�#�&Q:^��s{eA��+Ϟ�~��8��u,����c�j��K�Ƭ��Љm��a�T��n>=f_c ؤ��JS[�$'Q��F<	�ڽLZ^#�_��cw���7�lǺ�3n�/�s}���I|8�Dp͓�3̰�?���8iG;�^P�T�Y�X�-�6ny]V}N���)��Z�b�]o����ފ�f�,��g :����ؼ#)Wk�}қ���z��W�ː��S�2Ԉ�7�����&��n�b�OK�����������SzU8���>&Nc
�Y+��l�����/�I�!Zj#�9�q�!���z�1rd�p8�kfy��!��W�����V�+/<�C%�u�3Â��Eؒ��01��UD1P�pB�����+���A��	I��A�G��������yB��kD�C�rA���w^���1NU�l�'��|�tn��q���l;5��E���ܟ`z�8�ƫ>,�[��x�����U�!�2��|b��jv���[5w�ݔ7��d=�uT�S�3x�k�W#��(v��R����4>�J��'��N�˻���5V�wK1����A��l���
ֈFp���Q7�m?h���*�cw2��+��0�OU��S{��|���}l�X�'�s�𱴳=e�e��'{F9L�q��$����H���n�dx|��\�RPpN�[g����d�<��z�O�R Gح׏^Ƃ`.A�~ԋ�e���x���f�_,�tL���(Ѱ[����h���i)Ku� rP�*�ZBhN����Y��q�8*��8p��/?2����kR���t�6�ꍴ�Ȟ}�~�<`x�<,ڗP%M	[��ha����m�����nH�m���f*���iJ����G$�,��1��x�̀�^(�{���d� W�㚢=�aԳy���xMp�$ɻ~��5$�P�L��j!8_�)�'���5�?����v�R�	���{a|/������~�̅���;�@�X6pT����C(\����i�Z˂�wP�1e�VA���%6�{��Eu �eCW2��JQ?�*��1*v�<����e���D��]�g9ݼa�
���|=��M���.�2�.3A}0�sX�i���A�v����X����^٦Z�z��4��Kԑ�U^����߼v���_��͋�|�!�E`�5�T!x�$�
�p2uPV�J? �N��a�3Uk�E?>�6ė����ʁ�J~�i6�!��ՋT���Tq�k��,و��� ��*��H\X,A,7�����J��o0�R�{�����ᤍ��Z�⵭�&�����ۃi��(G�y�L�#(��70�+ы��׍�^:�i� +!�����ʐw4�v��M���m@�	�h-�������*R�L��4F~̓�J_�M�Ē0��~��g�⥘jO���>��$1���Ap#k����k�%rM1�ǟ<��.�`YF�o�9'G�pC�M|�
x@��@>9����ug~O���R#{H��H��}}<}�� 	"&�!3��F�z{W�b���Z��6r�$����T@�Ւ�!.H�-/�D�d�
�3��BMV���#���� U�(4���b �s��@�[��(`�貆��A�:�w�W��o}<�t�**}*�X3��C˘f���W�s�q6�,r�Z�4��thL�x���j�R�~��ѭ]U�M`�@I�R��<��|�Hv.:�~�cţ�b.�e�+䌬��b`gl��j��!�o�B���T���h�f�p/�����^Z.�8:�!��u���]=10B@��U�|�-�����B�<XU}K�w�S��,�y��V>��z�KϘA� �u��w0��>ҽYtN���8�S��q�������r��Da��tK�0�#h�02�X�3�mȵG��c�J�u6��B^�T���3��C��]ܿ���������-��ÐQB���W�>4�J�k���ևn,�_�=e���p KrCYD�V����b�O�g+���r��z_��#	g���2Rn��P Ն[̆%E�A.	��+��F�Tc�"��^���F�<�Z�l4�?X��Ŧ����3J�������}(K�M��pd}�j'`��f���a�޷��������Ϧr
"H*�ݲyJ�vk�~A�r��V��%a� �2'h��,U&��~c��4Hz���� ������'�/�-)o�|���)�޽	I��chY�^��/��aR@,�?�yx��BA1z��|彦�$����i��+	��4�A#N$x%E�p*(�r_�*���2����B�r
T�����F[�,�Y�1���Xֻݜ��#U����aַ�s|�Sltm^x��{]R~,>Sh;�j���n���:B|��+�`�ș<�>SF@4�&��+Z4 ,��-��.WW���L��?�t��5�*R)c��N��[�v�Yi����2��R@UD����N����Sl��%c/"�yrF+�t.��LB�\�~s7��{�<Z�����ڟe}�f��`�K��SC�&,�ߐ@�l��ٖc�v^�����.tR�,�4��Ѭ��Xq��wΕ��&������(pc��
���~ϐ�,E?`����Ϩ<F>�q�a�
%�*�R�v���{�j��t)(�v����pF=JV�㥳���zOê�Z�D!�������N�L��p�<��?�	۵d�?ӑ1L���7�>%����+[�3��l���!F�xC �)&�m;5�g��rO>�N�ya�tP D���n�}�e��Cang�hyvx״S{i��A�.�#ꀛ��k>����ŀu��o��=��̠��ڈ����g�u����_h��h_JB�q�Ӵ��DلzX��.���%]�}M	�G}q487X>]���Kݷ$yS܀�)`�&˟�R��j�D���p�Y�q �^��8�{,���"���(N�4�qϽ��Z.���ԤMӾ�>�D�X�/��Jn��PȽ�>LF��N�$���ڿ���.!͂�4N�h7�M�P̳�T^F��a���(���hR�c��Z�/W��i��DJR�G���QT|d�,t�_�F��p�
főj����J)Ɖ
$~��	r���M���.O
P�r��
�B�
��Q-�uGp�� 2EU�������v8,��U��D����H��]AT,���ch ef!������ Eۏ�ýjh�!�Ks�	Q��-6C����b��E�����_�ɕC�~��R�;��o���H��HN�'�c��]9$��2�#}+���uU?�Ζ�h��C+.��Ma�(g3���4j��3�^�p&�666&ʄ4�W9@��JO�R���S&����S��U|�r�.q>��D�W�����g���Oc �|S��#��ɼ��e��U��Pƣh���͉e�<8�kH�Y��h|H���4�i�'����Z��'��C�-�������O��`���S��y��i3aBr��8g@�-�n�y#��S�U��y���&r�P@:�����ڽ,]q���͕�7#��kc��La;�]���N��|��X,�o���NT4N�/�&/��ڂ�H����)�tݩf൉˙*��[�l~"���ytŭ�� g�{{`q�`��(�Ĕo�,Aj������1�I�b��G�@��du˦>M�|��p�����M���."e���tiܕ��7zv>��AdeQ�7�e��!� �j��]>��9��#����w����z����ۀ�kAA�Ye���d��6r
�P��[� ��\1l/Q���5/�O;�g�[F!�g�X[ג6�W|P��3mW��3N��;��di���
W�A���&g��K�~%ӓ�3q����,}*������F4OXU|7�5��]�`:VA4"�m�3\&�y�� l����nٻ�P��}�[����ޫ\?�ˣO�Co�~�V�����KO���=?Cf��)�*A��(n"c&
��T��ݜ�".N�M�W���",��zB\(7Y�-�'�W$l����rd�����]�A5��A}]qW�O�Yc�j՛���Aٕ��^[�1qj��eoy)��~������!�X|R�ԽN��	2�W�&tъ���7��W���͐%�nl��V�%QN�eʻ�c����SX�ћ����97T�Z�N ��(��=������r;B��@��E�R������dݍxxr�]0?��IƘ׃\!�My�c��dV�Rt=HA�F�g��܎Cs�G[���sw]��$P�;;٠�i�oJ����&sm��^�T�많���Mg�X uH�E.���,�����IR0�K^Ȳ���(�3=Df�7�G���B<=��Kz��Ϳb��+��XM��qp�z�(�,z�/�����䜨7m��#��_c�E���iH6-MysMy�l�z;�'<Xs޺���X�A�DOR�1/נMxp�w|�[�ˍV_D�m�:`�w+H��=����3��5�dg�kD�x�A!��ґ��ג���0tiIZ#�W�j�lh�j�@��B4�#Ɠ�
!VItE���z��,l�Q^��	1إ��p�>�,�3����Q��&Ύ2ǲC9"'�+P�%gʟDh`�۳̏18Ǽh��QU���6n���ȭd���~HR�uF�W.fք`=�8.JO�D&��s$	�ZdP�B�WiD����8�����)���k#q�U[��g"�Fc���ӈխ���~+P*T�"����_���J�S╰l��R��U�X�'�M ��UƐ�Z6�{�묻"�d5����{8�+t�{4�+�XF�X��-3�c�3��\h�Q�h_^'�Y�N��Ov����D�ߴ�xk�~���j�z)�-+��l;'�\����B�]�[������TǺ+���V���Fw��sr�7�[��)
�3���M�lHa&��?�l