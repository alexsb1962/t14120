��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aЫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��ƀPfƆ�������/�)����ǃc}�Қ����t�Eޑ���@m�37��=��t���F;�Q�Q��G�5����K@[G~��*� �ۭ�Q�6M7^�H~�K<17K�WF5�8-k� ��� ����.rĞ��En+�C�w��e�k)�5�Q�Z)��Qjc������fP�m�����*���c����D��lz�ֲP�:_�"'�X�W���ы��.v�9�����Bq-�� ��erh
�c�����Rյ&��.-��m6��dq��HB�=6�KQ|��pa����r*������.�{*�a�N��������&-SYDоwt/n�;�����.1؉E���F�y3YE!�y���t��].�z��p�D� q�g�Z����p�M�5:�:6P �>.�z�c�s�a�a��`^a,�t�)[$�����n\���*��r��'��Y��@(,�gi��zS�-��z�j��@#˹� ����q�@m=�ٵ��_���::�_~ͺ.��(���|�� v�:�W�ёA��'W�B6��G��:��}��B���v��K}M[�h,6)^[�Mg���E=�E`ɅV���d`��%��)�[$��o�߀�%_��H����,�j�P�vç��d���tW�x�&fR\�lA�RL|�f�q$ޚ�� |L����
R�L���|h�?�ȝx���q����W��s�{��Z�����ayZz|���`�hd�'�)s�s�[�}�I F]R���t�V�Vp�Z����[�,l$�Y���a*�)�:V��Q�C'D+�D�u�������S��h��8�0�=�	�.��;�
k�T�]E���рZ�(s]��/O+�(�LaHk�}Sz��+���QPl۩�?I�g�#V�D��M�s��ʡ�������U��hW1b�W�������G�1�l�V����D:����Z�=�<P<�/��'�����u(N5zq��lSTא���7�����\`R!|�+��i'��?�t�ۃ1�gj��������$΀�~zͶ�ʵ%:Ծ)O/ݐ=����Ԅێ�a��U�V
�2�$߄)dɥOC�T��f��^N�𘕓n�*��Lo�g��,F��:�m���ڢ]>؜�k�eF��J���+�dX�L�>���ED�T�����L<U��̤�X46�AP�A[`�X`���j�������6D�$��I���0�4V#X�`��/�k����&���TaV����]��4!���ؕ!���y|U��A�.�%D|��"��!X>8Ț^�bF��B�}����{�Kj�lN~�l��-����R���m��Wq����(�C<�﬘��в��0$Ĵ-�b�z8n
������!o[l�'��l�s�4��P��f��װyH��!�)˥�+|FN2��`�]l����V�L�E��y�2�R���^t�6��-Ż�+}�+ڦ�֛f�d���ٲQ��O�U5���	p!FEbc"�0������?���'�	֫�S�ى�c��Ŭ�b�ipÝ�q�[xC'v�-�I�F���>Żh�!�@Ŝ�5�=���z94��H	k��bcD�_��K�R��;�0�N���Q����X�[�K�<A���!�FB�+����X&�+m����xL���20��S��깖��#�ۊNLs��y�ؙ���&3q59�צQ�����'z�Қ��LN6m�Y��5�����j�����K��8\\cN�H���\u��I3�%[�-6m4�,(qS~�1Q��{����� x���Tt~��~*
d5h$��~ڹ��箴������[܏)�(�svZ������IW�j?`{o�RB���<$�'N4ڐ|�`+�Kb}b���/�����z�]g��尒(�J�/nGڛf��O}����0�����(������J�wv"[�d���u�)?.~��UF2�B�0�7�g�F��O��Ό�w;�\(����jC�H�λ��u�|`(˺�#&���»FN���UK�6=X����P�Q>R�=?�h^l*��Ju�?�}�-��!9Pl\;?�=�̮_}9"���x�u��c{��Dq��v��Յ�;B\�2�w'EU���V�w6&�/YQ��!��]�9����Cv��@�\��e���ȇO����4�޶?B<D6OY�^/)5֡k-�%�'J���}rV�"�����Ӵ�]�7�O2d��[���$�b�>��Z�:Z�-N�8�xF����f�̷��}N����_���W��mO��{ftܻ���/t�	�IR�?�CUH���UL4>>\�c�R*Kɇ�f��AC�G�k�p�T>Z�p$	�s����4!�Z�m0�6{z�?�D;�������j��dz���)j)�jGX���)��%�
���/�-�������C������t��ُ�`/��s�
�U�0�\���4�3.Z������>�L�Y���t��Cm����6ȏ����)T}�@��W���u�>���<&���|�7â+�;5S�Ր�#�`ݱ�G���"M]�3�8J\�&xA�jj	unp�vfS $B�p�<`#'�O���(���dX�s�ݲhc�gV��վT��̄�@j��L��;c�� ���'V�$� &p=�	!��c�Bd�y[G�/U UOQ�'��O�u߉�_(Y�?W@�&kG��R}����%���X�����ޚ9)D�����t2����_��;�؍�r�&2��o�:,��2�*9��QǮ]�d��PH~���l����t�4l�Zj���-9_��*;,}�j2+�:&��&%��>o'�Z�K��r$ѳ�F����*�/