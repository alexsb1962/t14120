��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����t|'�dWJ=8��A��9~5wukgwuAF���� ������'�$�$rٿ�\C����ӎ��ˁ2�O�-=�\�8�td1�^�������.��>�X�nwݰ�.�k�� Cwj0�c_�<*�iǼ�9	#/�5��}WX8v3Q� ������X���a'؛�,˄GgI�fD�S�6[X�����!�XѫX �&s`��h����;��jdc��������f�X�ذ:xyY��:0{��t48" ��{�bDI):��v�y�u/�l�����zFo�������/�&�h{�9Z�L�Tu��[h^N��ޓ���QDع�v��/ۨ^�����`pЮ���1,$����	c��2Ge��ֵYE?�`B=��ug�,+Q�]Cu��nl�><����+eX�1K����lZ�u1�_�u���a�Ꮄ�%��nظ9 YH��u��Z�9��k=���R����4���ݽ����|&�0Aq������~Σ��R���-��q��v��bH&e#ݓX���s������n�W;��{�m����*J���_c��t���i4���T��)<+\��},�)r�ڡL�����+�J;X�"��y���*�2���X��@mY�+��sI���Ar��7��'���=�s[��ZkL͙����,_ލY��u�wsw�3]��e�q��7�H������<������ľ���@�S�B���ݸ�<�V8J4t`� D@�c�uf��cX92���V�L�&�Ԓ����Y,]ba}xi2*{`��'�-��~�Cww�B�	�.Vf�`�������0SE�I��;>+��j�	�jNBz��Q���� E��ҥ[����29�I��m�7�j�Y}��;r��$��$%.Zm�A�a��r8��ޞ�Ǥ�!wP��5G@ER�@x��3��*@�f9<�����]��'+O�CX`5R�j�vv^Np�0�TY������A(���2�^x�����?���+:j�f(�Ƞ�K���f�z�;�g�풘bƃS�6�:���Gf���c������Ә~���1�ݳu�6��$�d�������4Bē����g����ߕwdtI(�9/�$�l�7^�I����n���mJmK0}�盏�L��tW9�`���*y�U�m2t��{PGS���ڤ�V���Z�w�7�;ZDH?��s���4� )��wG�@�3���u�����Ҡ�Y��3�s!ߨ�y� �#
{��a�Ba%n3OJ����z�zT�Ξ�>�aV�H�C�gU�xD�����z�]���5��	5���u&�'" �y-�4$/S#\�>W�?+I�"�9�v�^��H\]T$���$�_ޞ�,��2�5,r,��́��D�֛�&�����M�`b�[ ������ܴ�9�]�!g��bV��"�]rw�.�� g�6��b���.V�	���9�F��:82��HfkZ[,���
m,�%�a���J�}Õ��x��Q�x=7��݅A�kXczB>��ejи�w��(ٝ��0k���g#����Z�f \B|�qe��J���s=:�F)J��4,�%*Ņج z�3И.t{k�:�3�uKA7����!���E�i��J�����Hi����>��|*c/u�l��SS��*�BEj,��D;x%����t��n>[P�E���e�Ç"*ӣ��\���F�?�%rנ����5
,��"��4�[�{��
�^0�&-��H�>YvHJ�%U������V�j��GH�e��ek�]�t2Hf�y3y�ǡU�1��O��Ӹ��2�B�:ס�AE�X�.��U��t��B��:ר��6�Ď����T-6UŌc��M3!h1h�gɻ�-!J�u�X�9��l�T��H-���A�� ?�r:i�!T���*4`K���I#;}kwy���v��A����=�����v
?�=��E�rCa�qݭXą攇)�r��d+��՚?��Q���
%W�+*n��wi(�����= Mʺgm(:'��uH�ع��=!@�M؎����1�uK	�2��������֣�j���=��J<��G����=N[+`�0s������8��5FJ��.����#PQ[���r�K���kK
�~�y}�=�:a&��wZ�$7��td��C�9q��qDCK~�6��Z@|K���k{g.���T?�;�vu�:�鮀ɽ4��??D��4��V�$������r�h �-��1���~0٢R1�-�3�G���:�]���$%���?!KK�:��šI6P��,�Z�1-Xa:�� �lJ�$&�NMC��	�g\�&yQef�'+�����Ӂr�EgT�(4����k��@�v�hg�E s$��H���{>m׻x�_5��|�FJ���$�\�43���l��<����V��}��r��F���`� �̜��P��hc�T��9#�S����VɎ��
���N�"��1iJ�J��!��Bd��ѳ�<�5��K�E��E� ���
o�w˻Z�Խ����S����)nS`�nr�0�\f��q��1�*���sK�lcI} ,�.�iu���X���r�T���׼�e1�Y�d�y�g�����h.��	P�:}H�H(�k9������ܼ��6�G���N&:�,�J--�Y3�&�����vo���^S�*��-�"�፾i$��%�i@g��Ut�NQ7��! ��F���C�|9��?�q�\4��6��|�85&���((Y���v��G����1"�g�Q΀%�Vb�������(�!%�T��=���,j0���/����Ȇ9G��vF4�L�&^�D���}kX���<1 0�x�����8>����K�g0�ו�Қ�n�oT�6Z�H�-2p�H��<���	�ʌ#�!��?��sR%��K_�c��\�Œ��#w�$��P�h"��Sz�\�:+�xG�����p�NQ4ۍłP����"<>��Oě�ow�һ!_$H�E��l @:�|�`⍞9����c	��g� ���݃k��]n X��	�����fֲ��H�:�����}a�\F<���YAgt�KWNȔ-8#Ř0��Ay_���4���o6��
qUO�al��=P(�<i�Tv�������E'WpX)�y
�.ebj3�r�Y��P�
2A�5tLa���Ab�װ�Ҳ�H��ˏo�7�>��)P������cbzU�b�%��i�ѠԈ���]`Hgq1[(�"�����Mr��f�,�s�:�#"~Հ|�ڕ���� �f&2ҙ-L`���F�%����ࡄ��X@v?d{#�- E./�w���pԽk��
0�;ۀ�ٺ�wZ�y�	�7f��Dg�F��|�h�����>�*.ӸV
��S�:�p�wOH�ۋQܢ^�Ș�F���R�]zo��~�5�w!������J���	Q�yeB{��:`�-S5`����1�A-O}bh�&xY�n[�N�SDt��䨡��2jE��~�������)2\@�x�<�(�
u��ܮu�%��N(��W��/* ���E�ۇ���'�r�j6l�XrD��]���RUJ4:4/&ֱ�;�����1��n���5G)u���i�L�38ǍJ�{���D& �E�X���yԸi��zp^�f<��/��$�ޗ���6�����s��N��'D�܄!!AǗ���ML���Ջ=�;R�p�f�@�����z뻆G�	�>G��ʲ�e��$ǧ����s����Z O(�ɕ&9s���Q�Ya*"fXj��}�@���a�or��ѓ��2mF~���K&G[jר�;ޫ����d�ì�m
ԮQ�p7W߻��RON�$,!��U�P����5��=�<��A�U�DWg?sMip�<�Bڳm�w$����T�܉s�V��T�o�Ph���_�~��Y�������O����߬�Jiu���Ĥ6�1��*Z��/ P�t��+�O���ߡ8ۄEy�0;��-�*�:�3��g�I�%�y8 9��
ttEL|Np�[��2/���GjPs�s��gHp�p`fj�-��v�Ƞ���,�d�Нϩ�̼H[�D���S[� �E2��[DT#�����ח-`��b�*��i�g��� ����Ӏw��EĊ0����$nE�u���D�}��Ow���T$'���ý��T�9!�pW+$���/�W�Z�i:�h�y�+����oO$�{<��4�#і��,#T�H�U^|�cbA��β���5�l�o�� �d���1�ws#��0Ѹ2�%�X�O�U���z�Z����1�Y:��@�꺱���p����L����m��5%��	OO�#�-���u�?��K��A��ͺ�i�u�M>� G�N�$?��'�d}"�J�0��S;���o��O�*�?�g�/���T�f�S�OL!��t/��H���'g
��<�r�����i��r�Vx���:����znX(���T�g�ġ2h���:���Kc��Wh���y��0eԋ��H2���1%�9?��n�p�F=�l�-�u�9Y3}~-aFA5�懨;\?9�����:In7�^��em�r���6���J��]$T�G�1  |����"�ඨ���� K|�L'�T(Qh��O���H;A:a���s�����,;�2��G�j�c7tЎ�2�-�$��x������S�7��P����������b���{�܁Eּn���tE�$�p䷉l����?Z_h1!Am>A46������2�0�C@���۽�b���"�fj��%`��#`����n㤬�x�7�~�b2[,�)�814�#-�,�)��ɋ��G�BB�g14?k��yq�ie�-���x �C��b���ӲS�,�C�����[�{:�ʂYO��
F��)\E~u��A��&�r{^|j9u)y�v�/w��קuH��6��2O�����P���P�b[��EX���7r� ��a�ӿLg��l�>8i�1����n��Y
�H]�Hw;V'A�/�S<��I�L�q��-8��t�2�mW~Z��!;�ݚ��<�lH ��K��I�7g�Z~�~��5��s;=3Z�^� o�-�,,e��ο��y~�Fb�olN"�A�,��8���L̠��
8�q����%C΀(��)fP��#f��_eCq�>��v
�a���pG�̻D]�+�n�&_�����r7�M@��ͦ�t�0j��h��bZ��g��6�P����j.����y�W�7ٌ$8×w�֤��|ٌ�:�T��O{ܶ��õ��yG X?��Z���}��0�nu1�k�r΋�16���Y�Z�Z��&sEh\�ܒd��E�pI���=�&SP�D�PgW�F���Bq�e#ޓ�I�i�l"�tN��ֻ�.>Ok ?����^����o�C0�J[L�I���Ӈ �)�{m�$�B��熋ߧ�=I���jՆ���t���!ב��f�G"��<E���
��j�$Au���� �/���X��R2,�
k�7˟�{�SI<"�_����M�7�ވ�M������t��8�HB\�<Mό�0P����r�'u�#�tr�����*�I�i,�z8��
�:��Pw"+��o�?qP`[���BM+Jv���3��k=<^�m�W������"�k��gʳ�7V�������J{2_�[_�����gsΦ^q~F_�+k�Y�� L����g&6���SQ�H�.���9�mP%��w@U���Ɨ��ac˾Mn�����<���	Gc��h��G{?/� ���#��t|��*I+T��z�X9�9�p�1����P�
·t��ʭʼ��r�s���U2�b�2_TT,�p�>���~���tdFֱw��$�{|�1�Z9LoC�x[�����(�J�	�����,�6�u��!=22�#=��|:�l�QW���tz�I�1HR��j�N��׼��N�e���!HxD���Ԥ&�_�T"�?!m4�m��m,�,��Qj;�c*�DY���-!��uY�Y��p�ۘ�&'a!A�L3�pܧ�,�oo�L����m'ݠ'iN�Wa��Ⱥ�!�����:02�[Xh��s������V��ŗ�^a��vB	
�{��`f�u���}��bWv�m�voj�h�5� +ZS�hk���s0k�T�F^��6bU:^�7�嫪f��DJu[J��Hf��mgDs:�jsB��o�jB/��*_ks;���$�D��^1��'1;�C��$�˴K��e�O!~�3ҵ
\n�8�yt�hw��׺G�h	�An�!�-���4�>�ڋ�g���n��C�7+��u��Wz|?�b�9G��,�PRMH�-�����t����r~/���Ͻ9�S,��h�QxP��s�46*l&��l�l3x��Z{'��T	��5�D��
Cz�y5�pBx��PL�z��� �c�PN�B�qE�:�(��GRW[v^��@lN]qC�=�ƀ�`��{�Z�����5w��<D0�!>��)X1��ؾ��sj؉ԗ�U�b�N4�%�:���S�4'��Qy����S7U����D���ؕ	�W+P��Eq�D�n:ѲnB�6���OI��ZMB�QV{5�i P�+��+<��,�����؃w��ƥ9d�	��ڋ�u��hwcI��1W�!u�.���o/7�~^O�R��q��1+���ư]����j�Rl᳾�\A�F`WV�0�GX���|zU�F��9P�����!�["0V�;�<���	�?
%d�A��U�X�ޝ3SH=K�$x��2��r���#����a
�[|�r���A�gd��D�B�4訳�S4��mo.�B������+*B]���#`���g\��Q\-�T+��N'vPn� �6;��s��3��XlZ����&���i�4��&C��O�Ul��j�셵��g�>p��p�������pͬ�����;�9��s�BYFY�2����\"~e��_<?hx��Ho!}�L�F^�c�F���p#�V�=w���ByB�+a��j�n�{)�<#|�0@[��e��YO���;�w���W��a1�G��"��GE�
�,V��; Ȫ����=t���Mc�m;U{�o��4�D�Cd�d��n�/�g8�y��ҥ��X�'Uwb/F�[�7F�-�n��[�X������Y��3ܨ���Yv�'�kԤL:��`�+�3�{���H&�S	t��kjO����8��8��4@��ݹ&�2�)��0�)���{�:w�2���y�#��Iv�^yzŏ7=}��'	@�v��U��k37	֙D�+�ʍGp#�n��B_w��Rq����A���$x��q�k@6��Zmua��`x;�����WwQ1q���l�g��F7a�jh�͠�+��
e����	x['�S�G��a���Gؔ��
��l^aR$w�h9�$xs]�U�{L���Y먟���b����m�]��&fX��K�����v�O���0�0%���5���}���;��{jn���Gu>7VY� 
���B
@�p+��k x��D�q-zC�t�����@��*�oNRn(���/�Tn�4��K!�L1����*j�@��p'������@�`��m�5�\���=���8���e�|5���+��,�n���I���Rw��uΙ�.�R�@<�7��W�H4ğ?u��N���(i��Q@�t[[����0
�^Mn_k�
�?�`a��Nm)��-8���Ec�!����)��Ӗ�~9���9���%\@�uT�0�'z_]jz��hEt�<�GgSb6l�2��M���p�7۽u�_��FM���9���@/��0�ǖ7��<�P.5��J���ym�?���5{O�f���h��خQ�*��w��#�EO{&�o|�u�=�J�$�XH��i��"��ϛ��r���hw�u Sw@��{PQ�UùA�A��wjg᥂ ��-(�aYP�t��K���d��� r~���η�N�'8�1o���U�7����3B0	�-<�7��p��q�gEiv�?�����p3��D�V^��U����i�<ȯP���-���t��!��KB5�9�lAJ	�:!2c��d�g}���u}�X*����lė�^^�۟:�-��p��vTW�����WX����E��}��U~o��R�9��,������k=����5���ݣ�s��Cv�Eˡ������o�lUIR���	�_;���v���5�U�>S����5�Pi�Ts��� ���v��*������kE��ꉘ&�k4��[j�`;��m\�tER���*l+z�5����_f��s uL?�-2���8z�[����FUն�U�*���S߱6h	��T�� ����Xd�bLS�H���@DH�݌*�E��V"t�N�����C��&�@��m�'���|\�,�7��/S�:�ǉ_^e�� �1��T�y�qW��DRV��~�nN9���8vp��D9>S��7�>��9XP-p(6?u�M�G��Gb�:��FNP!I��)z`*�G��*D���~��u����UX��+PÀ�fN��\]%��i�^:�AK��4�TxM|�bAb�\�I9l)��͎���������_��*a�ـ�X0X�lʶ�/��ù_�����f2��Y<b��e�t�ֻ�	7
\d����u��X�8\G��͊VF@F�ITȧ/1�a��	���܆|ǣ�~���M�h��>��[� 	M�@Z���2��Y
<�T�\'�}��]��\� /EyKUЩVL�!������y��q$�����{$��k�HhY�ѥ`{��8�� zg�����<�)���u��B��D:+ʗl��-��t+-�~��[��S��0S*�2C��ݾ�DI���6��{e��C�>�N^�f?BwF(��B�׏Q�~����!d�
�uV����pF�e��,��L3s�<�CU���=�J\U�>k�.��[�V|�§����('��G��>�<v�+�P��7��o�G�����7���+96��{'�%u$�
�v@�YHx�� %�^��u8�xj���[���*��̔b�֐��#�J��,h�#���ݥ(-�b^���,/���̌Գ�� ����?��Bl�C�@�_�4>�(�G�{���=��жl���b�%|{�a�Y��Jt�6����#�t�~��%���05Q�I<8���l�3������Q�|Խ�9�y���TIZw#T��~����+}M�[�09�K�Z�i���H%:��P�#o��1�ȼ�bk�.})��_|	�Ձ�P���"�	�p��`̌�@���ъW��R�&WGA>��+�u��i��n$XO҃b����_�L�zu)���Qd�*�_d<�R�<�;�{��Q�9P������� �2�Y��)]��t�0�8X�>O�	�.��"�����3 �����{B?S��WF���&�)Θ�`�l&9F?sCk��hZ$C�����J�`a�������f߈@"�RN��(�Of=�yfk��d��j_7�2Q�l(8 �D ����{^}Ǧf]���3�IpU~M )UpVov![$߁C�^ a�kv-��J��>�O��:��0����nzn�E\`�p���q�� �+�O�#Y ;y��
����*�iv���S�H��
H2��V�|�Tw����HZw�:�ekV[��a�6Z���g�p�*:��>˗6�2����zʰ���^����.�nQ$8�
x
D&w`�s��O�F��� �b�!:��ژ�6��ϖ�ڎ�Ju�sh�����mi�&�T�?U,)��C��'���ȇ�S�����Nu�����ku�h\.���/ݛ�C�_ń�9�ݽ�ru1�!0�A�5�^�5�9n�DƁ@хr�c�ĕ�w%���d��>���3QUv.�'���N<��A?����*�oi�Z�14���V���l���V����(!E��?Y@���6�rK�-1a���*q�S]"�@��}[`� N�D�X'T�h����Υ��[�kW�at��Cxä$���ݔ�>��Z�>���V�S7�1o�+l�[B�QBcx��5�X���2���-���,����{g'� ��þm��7��|P�`�#{+Y�[��u-��+#�Ys���:n��Fh~8�xK��[��Zr&ǩ5��V�<l�RK�r�w��N��h�t]2I��N�xΘ/#�y��q�\��'��S�)���3o�f�E�(]K�P�˴ɣ�z3$]�'�߫\�.�uX��0��2���L��!OX�����p:��2�H�U]:��%86�
���d	�5���w("����*����-�B��~�7��������(�ͦ8�i���	��j��P�4�.��y�n"u1Ezb�yVD>Ck)�8�0K�|V��0���U1�Syz8�	�'�K^�e�|�m�ı�|�T�)�޾��39hO���x���|}��q��iD�����?�|��N��v���b�@�~����
�&��#@n�N�*�ޓcn�J]Ҿ����yg�e-�AE�M�������.�>�j����aS�=�
��؉�	��ܕ\��G��ٻ�� �H��᪣JT�M��ko��� V�{���ۋ%���U�@ĉ���1�T;c�~A8ULW�>*ǩ��*/�\���ǆ��F6���r��`����Q@F+T��{VP�����*JluJ�P�*�N� o��n��{�=��©����8��!4E&�G���$���Ym������8L��ccBOj7��ey:���VO����->k-�'��#���$E:��p%�IgT.��1��E�NًK��+6�����>#�[�xP����^�x|M�S���x��2�8L~�T�0�߉{m�@IE:|�3lո1&�\Q#���~-,�a���l��E����_}g�\���ȃʽ����Y��tx\]N)��<uyF��c��5]W��)�K3�`N)|U�a�ϭ"�4��p�����`J��y��B���Y�Jf�t `æ���c_W���Lx6�,����Ģ���@��˓��1��|��!�����\}�����X�/2b��Rb�~u��PRt�EGɭp�wJu��k\�-2+��E�w	�^G;�PՅ�RQ��� �(E�"�3�e�N�/44��s�bW~����4�6gF��ϼ��a4#���w�70�U+� {��[�G~�X�FN��
���7�U�di~&Gu@>�-o�pO���Ƨ���}�W������v���a;�;�4Z�1f���9L�̀z��~;`�1I�#,{��s3c����O����#�Ĵ�R��g ���}Y-������A���K׋�r�?@B�SłCvԠo��IT�������Ӈ��ZI�إO���I��t�sN+��㲣�"�W�,n~�HR���R��E%Ým�K��V+>#��>p[@3������|�_Zb��0�oL�������S�iL�����෸b���Jjκ�J�b�\6w~���t�Xa���PG��W�wj�~�.��P4U9A'��'������IrE B^O��1~�t]��0���wF�����&�d�>��˽���NRD��-Z狶���3ƳZ���$Y�N��Hv&g�w�D�P���vjP_���-��f����P:_w���C��h0c�k\W��4��-�)���*q�@0d��̕�A�
lI`w�kK��dP6'R�X��&p4W���҅��M�]�P�%C�wrT�M �V!a��Z���Q�/���N��X�N�������wc�����I��:Q�:���[�Rޖ�@(�󅡙H��t��<ߞ+Z����j����d*&+e�-�q@��QM���9����Ĝ��&F̊�7�u��;��o?Aݵ��{ T�%I�5"=��R��
��̋���%<��ZLj׎�-���P����;��"l�],�$�]B�`I��8�zH�j7�-���)�b���@�7ף3��ᰢ 9n�������B��1ܗ��N��'�f��� �o|�Sj��aoKw8�F�vg ��S��z	�<h�6Ѿ�{�&��+��-_�}�o�`$: F{W9Z�q��f���y�.�I$'"Eq���Z,��!���N���:M�F�x�$3K�Y&<���U��<&p!��&e�
%��Ũk�i��Tg�h,�N�N�Aa���b~��:�?׈q��R��4CX���p�q�'�zq�3ɣ��R���G��"Ϙ*3B,3m>�%~���ȹT0f�*γ��g����c��>��4t�VL{��>?����Y�?�	��s	��˂���8B���T�fKG���p��b�2��e�]�#;�j�C��8)�2c���=�J�/������YH��b��k���i���S��9D� ��6��9�'�%��PF�$n�yl⟨�Me\��=Hx�5�8?C���u�M��Ri�����������|hI u֑>V}F;���a�hûʊKr������tKq�MG/A>��s̈́�Ȱǀo0����"����pP�H)��T�%3�aғö�<9�D��A˔��ъ���يIcY�Qq��UU�w��I���������0���Sc��{���&Ph�(˜?��z�n�q������'�'\���v玻� �	���慈�ly9�ZO����dJ�;�9�w�;��m��J�/���}������Q�hjZxd�U�x<���x��k�ĭa�P�j��<�Q����W0~iS�vEf,�_m��`E54��(�W(�lT�G�ڶ���mvwޔ+fH��7�P�����^(f�1��,�<�6��1�xÁ�5o���l���2�p'��bWV��5RzȌ���!^l���h�*Vx��uo*�Gʧ��HZ�1OV��b���O^Hļ��%-gҫ'�LF�5S��k
�A9p�[]+���k�X��eP8e���4�CUXv|�Tra��ih�z�����."k�^�%xsk�v�����.2��@ΞAS"�t�@lhH�y�����f�eo�	5���zs�I���#��k��jG'���u-��4��d�wL~���R���ׄ(c�^�<���~sq�5��R>y��6�d7�ȱTB�T P�Kx��hR+U�*������f��ʓ��o��s�PH`fI�_b��Fx�^��W�
=MuU[���6s�0�WnB|;}mF�`Z�;L��7�p�5�A��A����P��)=]��,�l�U�j"^xq�',���F����W��	e�Z��a:���@�����= �������`�_Vrk�f�ٍ
os#��5�4ae�!bي��*���	6`�w���c��Ѷ������������9��ּ�c�#�}`I������࿨74��_@G문�Y}=��B{�=y��t��̿g�[Zؔ����B�A��v���1;vW<���<�x���d�Օ�Ό�G_����W�E�������˦5�[�>�4c�a,G���������)��Ec*�l�ϳ)�ũ��I�1P��R� ��3����#�0Db�Ż����O~��T��* :���H������|���#ɥ\/+�����W�s��((f 6����8�Єݛ�f�7���'r3`�lo�]���Cx����ܟ��"�&�GaY��rS/&�@�"/g+��a�Ĭ��;�����&O2J}��B�	|=�T�愕��l�t��&ׯ<�M_����mv����V.�\:�|H�n=�}ES龭�G�����#�uޙ�u_������>F^fU{<���\$��fU��C"rq�D�=��}�JT	Ud{%P~���i�v=����Y��ǔ�K4��K�)7������#��謯E����卑GJ?����,Dq3x��g�VPJR�>6-�  �Gt�Lo�D���~� ��&Q,�Ђ�,mؽ��Ɣs*J����V1�#�8 @b�:ۂn./dQ6�qi_�N|�+�߻�_I,m�s6d�MnE691-:����%���4����u�Ŋ�9�}h�����\cm�w�[Ή�qԐܮ�%���C��ڱ~�7r^�OアYm\w~���H���JH"0�&����9�=�A��8�����/zf�k��'9�׀̞�tk	��'�`G2-�?I�$_�X��w7s*��J_�Z��Du��P�p:$�ߴ�;4Y��Q�5��x����|�s3�Y䮸�~yU5�p��ބzK�&wޝ)�NR
9K� 2��@N���C�rC�R����jK8&�&kt9ށ���P���[�*֋Z��i�ŭ�f���Q!�n��=�bҹ����3e������������1��G����zh�{����A0*��@�6k�����eG��xQ'(�뛛OE�_�6Z(��GR�d�����T]g��w��Os�g9]]`z�_���ª{�I �@��>!�8��V%��K���*{���8��Ց��)�L��n�e����ٌDH5$�d��L߭#�jx]����;r�1��N�0���8�GlS{/��PU�Ap���8�� �9f�I䱈�:-x'�#�k�S�r$������E0��%�gM�������N%�o{ARz��M5�wEE�yF� .�ZQJ�z~r������ǡ��4�L!s�"}���zA�:��ɊN�ک2F����p��m��p��Hsgh�Uc��sń�At^+\+�m�,��gb���o�O��d�{s<<��-�m��q��*�	��-!"�FL� ϱ�j�⩌������BI�2:s�An+Tz�{���K�.�N6�&/�o��?�+�������_4�%�g�ԧ�fwH0&%���M2��c7x6�[𩜺��1 ��m��2�\~�ߪc�7�|-3�9T�Օ�GM��_�:�{�閗oL�b&F�]͇���3S���'�h����W��*�W
W�7�('�������`@��EO�:�.�ֲ��[ĎUT�����9H&��-(���n�$�ť���� ��ӊ�X?�EU64|��(��E=q�9\ʹ'�S��(
o�J%$s
��ǿ�n��뷻��h��'q�*��+Ӓ�]�������M5�֘G���TѽO�&4vfS�G����?S�-�7���E��I{�Ј�����i�5�8֙)�����ӼW�*P��L�FX�J�T�ƺr}���U��P�)dx>�jRVR�[(>�᪈��mG��$JR��d�y�Z!-���t��@"qx���.�y�r�NG �f���O����L��&G�`>@^^�u��>1d)�Hn���P�X��o7����r�y^,���{�I�X�����RgDS��F�|0��C�~%�R�a����BTL��@�������$��*�0��U�"�
�Ύ�7�㥬Ó �@,�h�(�B�塣�厧x�a�A����qqY��J��l��/=E\�_nHx��<��q����v�i�#�9sſk�dز����:�l?7Jak�)��D3������36O� ɭ.���@���[���
��%��f�BO��}�`M��/y*ư�I��;ⅈ҃�L���������g!�H՝�T`n�"�"4��2�rgk�Qb�m:pO�
0�G1M!�:����庵=���еu�'�w��8���ģJ@v{K�-��˄ q$�p��S��XM�:�ţ��К��{��5�;�@Q��`�F��&�߸6�W���'~O�>S ���X��[�7�1�u�F_yE��U�[�hb�L����+�\����� 1�=馉�}�+s��M
��-	����)6Ѽ������T5����GT%$΅*bf��(��A䙍�m6y*A����d��`g�K�l�y�����?���z�����X���Ä$��)8Jޱ�9�>�~ΰ�3t�&��kڜ�{���m>�F����ЯH�t�خ��� ���l���j������~a�;;�XG��#�H�[��:[��P�T8`_o���pև�04���$#o���~v��t�� �6��Ǥ���I{z�������;ȹ4{bؖ���G=�+�a>�Lm�	���r�ˌM@�CD����}��U;g�Ā�oS�a?���_�X��rD؝��f��o=��PV��J|�@
����|��y���
x�<t�z�j��Y���@hgΨ|�
���������~�wh���MN�M�����B��;TDF�j�aQ�1@s\���8����@J`N�X N�
<7چ��-�r|0�YO���/n��mup���&y[�����r\2��M��֐e�㗨|��0�r}_�U�3^�O��!�g��%��tJe�e����?�L< ��̳�B�Ɖ�*�#N4��v������/B�7��u2�v+���Ф��A����u�L��&껶0��������V�l�(J������`p�knGbR�PXl�!�>9�aB�}CJg N���b��t�K4�e�u� �_?��~~�����W��u��':r�Iz�g�j>z�R/n5�w�ez�3Tʱ*������S�;�M�q�06Hӡ�~���Q~�P�Cf�Wٖ��Ͻy��Q�'����y%��gXX>ʥ�l͂1��
Ӻ��ΐ�G+=�+xu
�R@i�ɖ����Ɍ��t�E�.G���t�p�*�\�jG[D5�uJm���̈́�=��P��� E�@���E[������mC�3�:el�%mٌ���ۊ?����w�I�q��qϩϝ��כw"T=A-gP�� tƈ�_
� D� �8(�֖��z�GHQ��-��-)f�Bvs5�A�Z���	C`Ӄ��[�M�mZ�Ֆ�,N�{5��k!�@H���X.������~Ń�
ڇ���-�3��֩%�^��QE1�k+i�0}�o� (��騏g����t(6���L��Ɨ��[��P���8��g�=5�6��6�٠�JT|���l*H�R
��c�-�`�{��&�4cv<�-��VR(�
�Z�J���� SHRjlV����V�!jKq=�VZ�Ϻ�*A�nN��?��yzm*ݚ����[������h�8��5K��a��pF����%?�>��a���`��#s\��h�Oߠoj|�uz��Ҍ�=a|�H���.�DAY̳@vզ��w�c�$3�P���՚������H�D��6,C�;ψU���'D��?�=#�����}�	������UV��on�����a�J*�k&=d�����a��K�-�Hu��Y�]ӝ�q�g������J4�u���!Ŷ��Zg�� �,/�to+͇�Ϫ& ���J���!��H��q�zx�X���l�J·���|d�ZFOɎ����0XcRf7���W<��eo��Y�d�:10���Gwg�|����7-�U�ً��3�_HmM)�J��H�|�Y���A�V��mQ�'�'�]$��\�q��D>!Ǎ�"a��[?����ҟ�������,B����iQahR����;�h�ZY���D�O-5��(�e�m?[���>�[���q��U?�(`��_�a�D (��z��Nhʖ,����%=aV;�00�����#'�@^�l�u:���豳5��ܲ�^zK�gh�B��Wh1k��H����/pӉj��1�sC���d�y���B�]6�%r���/S"^{�}*��!i-��1�#$��>b} �a޽�TD\C[�&xB���`@8u(� ���d3j���+�8):�t���\#�9>��o�����E"�a<8u��w��E���#�$"��@;�q�+kB��z�A���>���c��:;�k5�bd���&5�"�Y�V�d9��!Sj�C�ؑ��~o9A�X���$��d�r��'��=�aT�
8B=)�.�����b1^<1�35�Ӷ.vl�+�S&Ѫr�G����8_y�="�V�ŮF�h�;X5�@�M�����0�������Nͫ����=���s@,�,���g�vU����4�LW]eS�Y��)+⍳�Dl-+���4%q��hgL��V�,���,]��* a�ǌ�V����B��>��z͐v$@�[�^0�"!и�P�P�*���"]>2G����pC�g|�T'�.7=�.-���@���� /?4�9:s5�K[^V�
Z�^v>�g#���p�X�������@��j�$��C�OS헛r�,h���a%m��;=����E��8��V@� ;��t~�Zh3�.�ʺ��&uh���J������_��t�Z���`l����