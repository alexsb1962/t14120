��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:��������uA��@��y���<����xDET>��W�����C%�=U����3v���hj��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ��o��}��
�;Q��Z\�"}b���tgQ��V]-�`X�L��ڨ�)OKe�%�V<%���C"I��!�X�n��m��N�g�8���Ґ�m�}=h����a�Ӡuj�� �эat�>V�Bw}�3p�d�ATռ�~xr�U�i���nP�� ��U�h"��U[W"9�?����p��1Ԇ�%�1�'�?^��Yfj<��ǐp9~s�d@t2*�{E��롌A{�皼i��*x����n��Aal�<s��I�F$&�lc?d��(��sV#,l�ց	�PGB2Y6��^V~#����o(D��Ei?y��n�l>)��S@*���3���Y�X��D����0��C􁭷�k�~>m[8�jT�;�܁����΂)�=��T��.���P>��3���N�W�?9$��*|�)�ս>-��x�\�i~=I9�g��m7�O�z�p�1�v�M��݃�����+���"�pvd�""�4t��jV������d'���/*�Kp�U�ݱfEf"��|�F΢��_
!\���Ag��M�\>@4�VR~h���L3���^�@	�����g�]�y����ketɭ�l�dR�� &y��'M��B�l B��F�����U��/|��ͭ�Qu���i���T�P�J��7��ܴ���v� 7�Ӯ�F1^n�&��=�ژ��oCj�t��}V���"��{��*E����l@2��G�7����ś�TQ]П�Kf����\�z��9��C+�@�y���ր�}NS�x�KPK%�c�l��᳕q�7���~~��eɣ��/�m�0����R��@��.͜�i����a��+mB�C��� ˇ6d�����S9z�bn'�r��}���͋W��)���F&�=���8���0R�&c���I���7P�p֓��R�6����m��%H �������k�s�*D#^Gs�La�$������2��fc_�be"���l1�7`
�9�g`��P��ȟ�KXUΆl��Pג�{�$��}��YD���(}� ��Qye��,p#���IJ��V�MinF�&SJ7�h��wͥ�c�⪱��2�?^ ̔�٫�p�E�F>g�;���71H�[*�	0HCu�\)��X�4�GR��2��WU��_�E�>5�o�	�#���#�ڻ����� �?Q;����X̳~S���:;�{
D��7���A"cm'V���[�����&����{��;�=�������ڸIR_	r�v:��XBU��/���A��%`�*w��VZZtZ� 9ʆV�>���5��=���������ą♵
i~i?����������	�F�s~��	��59,Y��Q��a�|^{M^������Q\�!�[��<�W:�*�d��2x֓[2�H�Aoez����~c8m@�#��DL�o�?�7�
cXۅ�ϳniML������(R��<��۔��+���	��]�ǁ��<�U��;�eTV�!i������ː�s��ߴ�a͗bG��� Sb8;�$J*��$	?���m�7�uk���1����[s�a�**jߣ>5Q���
B��'���b�
n�e�k�����m>����B2c%l�϶�v�_���YF�(e��D����ny�2����dPcX�^P�}e�H�[����Tp�L<�Т���p���r������ ��Z�K���Ǟ �؃�%��Ƃ���'p����=4N���`��j�+S���,���9[?O^��)��צ�}��VC�Ag�!�}�6�A��
|�1�a�zD�Ha�⻫�͚�"R��O�iw	d=:$^�b3����p�hk��t�Í&-�|,̈́i�C+d�Tc�WHLR�R��pA��P����\SN����5�5,}�"����,���p�œO���F�25w=3af�*i�@������0"��U+O�ͺA�H�I\��[�HAe��bE��f�8�����S��o�9�Sq���g�c�k�C/��.�M������c�[z�k%#x,�4��V��),�k�7�� :UfC�/�O���H�yk\��{aB�[_�KhB��E��C-p(�"��՝Ҏ�fY+Mm�QP�s�H�^���[���E�/2�q'<�MDk���>�a�P�.3�����;u�S�H��G*4c��y����f����K	��}I�+��لI�cW�V����h��1e`�S��NC
�i�e����f���O~�7�4Ʋ^�����������޻���0�G3R��-u���¦�KFZv���YZ``6��ځ�0����(,2������]��N�8~��H�,-�d��j`�݌D������>?<jX!�@1��у���*�%g5*
r��8�+��&8�~Ow��!ͮ��bi���\���N3���Eh���GC�5�p��I�l4\BM����CN�A��ٟ��)��7��1���	�ϜQ$�%�{w��WW��Ԏ*�{N80�30eu�c��d҂���Y�~��L����E�>A���G2�ex{]���/XcϢ� �(������ҵi�&���'�΀�3;mj}%Y&׸t縲�$����Fx!3�;	S�yf���,�b�+/P�S��.����,�e{rg��v��I��I�Te:h$�n:�fƱ�q�Dg�K`X�T�x{5��S�3��	9bc95�S[�/^%|�:�$��^[���|K�����c48�aQ8p�J�(���(�'��`d��o_�/�Z({�bV�{��JYrB�<�+(�(�}S�����t �\Pe�'�ɖ-Ң~<L:7ʍޢm4�O'��ry���a�����fP�fU�Z�/�~;U�����M�?Vj}��G]~⣓%��Q��5O��i(�k�%�ip%�"���W�����]��ʟvD&!��鍈��8�N��*	�-oA~ NW@�S�r!�����~�ƿ<�ݫ6�|�ǲ����m�zN@��3�3f��G���/�CI߈K��}��r���PGCu��*���o"&B?��Ǐ�X�͢�%u|Ď�N��<ᣒ�2��$9��%��$��O2&"�>Պ��[u�a��o�(�Tse�|��`[���F{}�0?_Χ�C�X�"�.'�}#X}d�q�N���_'�E�W����:�+
�����`�V��ދA�6P3y"5y�|�����Xm#tP�3m�.�3��1i������8�����d�PO-]q�p��*�f�1{��Q���m�w�n0.�i��}y�"5*�F��1���M���!n-���DR���3�fQ��Vz=��^N�2����
dP�bu|
!ڧZŖ|�p�s<�¿A��룑���ڋ���z5Z��oL;�|24��1���BQ��aR@ԘC�=/`����1�#���'T��ݾ��|9��*b
u����3����y��nަ �����5�gAh�!�&P��6�}�.�Q����E,ڳĪ�k��<c�P�_
�i�̜\@��Aqb��-E$�����c���@b���@������5��^��ww��}���J���Uf�y�,���Q�/-/��y<%ZPZ�MdB�o'&n��L��sVwo&bI��������?&RCg�M���Ì���r'\ <��4| ['�>>�����x��ZQ�	pi3�Zzi,k��my9��Ub��"�7�f	��>��!����DȄ^,_�$(S��F ���h�Ԡ�Sد�
,2������հ�0����(�4�!���tс�eL�L���bγMl���3԰�NbԻ(#.0݅����� ���w`CKJlS�?�PHMK�^m,f &|@�K�V�'�%!i�jz���7b����p�G���Ó����y��8�Z�q�>�7��t���l��i3�R�>Zq���U��69���uT�'�Q+�_���<`����&��:�>5�6\���BQw{�*Rn��qgvq&�_;y�]�>�7�i���y�]����:����
hHG���5��^BO/�tQ���%Y�=�� I�Z�����I�L,#INf���+@�v��r�hp��F�3t,�P(E�[��N3������0����s4P�c��+�����B忯�X�Jm�;���'#� ��ŇA�4~����Y����s��'7�uez:r'�H[��j�_� �iQ	�)۝c���j��V���qX><�(���&��2��ʩ�����$��y�S��R��o�0��� �=՗���N�	â@�� ��gy�q�*/�Ҋ�~���Z�In;{���\�bj���]$?�=��<&�F���>�%l��I`��V͒~IXC�;:>0�,�!J�ye�C��N�ku�٢#�����)��ֳ�������D�ޤ[\I�d�z.�9��|ۧU�q�:O�y�Ӕ�n���I�Ĵ�T�b�j�L�� 3�kY"|�Kf�_Fa���:��
��V]x<�q��G�i�{��@i��M��@Go[����3H �z��M�!�rdC�k�fk�,Xk�������9D�hpf��Z��`�b�m�����5���h~���
� �Pi���ۻb/#���?�;�2�3��$9�&K
x��ᘑ�W~�������V%>O'w	6�^#p�$�6��u|�|���_*e�3�_�m^Ce���e�-�#^F�U!�i�w�(��8�3x��ik���`{��)Q���hXKŦ�Џ�us�c�f���n��҃�v�o]6*�\�vRE����!�-Hj��U+�M���s(њ���L#\v�Qr���#h�U�S�m�yE
�{ΉHC��)���������ޘ����`�.�-C�"���?�t��>)�7���)����I�8���"�r)���v���Y�<X� X4��L^4�r��+e���=�Hk��-U�+k�0c'W/�h�8 ��(�K׸�������� e��RϨDz�0J��ܕwUm���gpM/3�,eU<T��ѧ�8M�k�Q�/s;�!?xuQ��#�(�m�&t�I��p�'z�:I�VR.���O��闐��(Uv]�Y;iO=u��-I^�?��]����d����-��(R=�^�UwD�i�������(��zP�(lĉr#�J�p����E0a����=qX^��]��۟X��L�"����wd�Brm�q;��l��Ђ���g�bw����W�,�(O-�hU�� (
���Z��yZ�{�N�v%}�3Ja1?a��1�����r���R��R(Ǖ'�Gm�W+%��`�tIA���O!�a��/U6 �<�%-L�����!�J$�RX���T���G�Ng֘]�(���dq�q�g�i�zU����/���][n~�`�����Z�Q�C�qN�,��贅?=0�ޅ9(���^���1�wJ5R�NE�p%p2b���P��g��"ۺ�ś&Jkz�z�.[� �V������U�����*)���md��q�JN|P�X0�t�P
���ᵢA�#��`�4���'��=�\������=��ǧz"kjnW�bne���5�ۻ���!�P���X�bn�Pc|	��ċ0����A3>b�������J�H��m<0��ᕚ�>�:�d��lX�*՛�G��8dU|���PWn����%����~+4��}=s�ė�yx�l���q�W�+_cO[+OZU��]�O!E-�B.�WxI��֨?	�~�Rr�-{�����l�g= 0sh0l�t�)��܇�`�rk A7�&�&}��u�nː�ƣe��Q�1B�P�n��F�pa������������Օ����c��0�>0���hf�Sv7��А��ߗ`v	u,��3��Zv~Nq`N_8o�f;�B=uj��
��;8'gs.�Nx�xmx�h�'?!����|o���H{tp�u�vbF�������O�,6��Y�`v����ɢe8�����cTX���BY�5����?����1Y�O6�	V�g���,gq�z .Q�fZ� �� >-�q�A2�T���ڻ�{�_@�%���W7#��l�^�S61F<��8�ה�~��S0��rQ�6���	#����C$����+��i7r�t�5wI��$�l7��M#js$0���� ��XY�ɧ������K�*��м��|?���;łK�����v��P�12�\�T�q��G�^InX�Bo�i���	����T���!/�́:4@{1,=�L@ȟ��R��Pw�gU�9�7�u�^���S0�!��⋐�(���7���c.���w�]���*n����0Y�*_[�g` .�4r��C�b�y4;,g�t74��4��y��Zl
a��+�X.x�2�Ł�*{�`�([�V�C$��x���N�%����~;l(C���ak"Qӛ��c�ǑE���mW������>5(����{��X��������t`�&�}Z���&
<}����e�GR~�N���
fg��U�:n��֢H�"-d��ͷ%�����EƩ�`Y��t9�a*�@�
��gK�s��Y�<P"�+>��c�;��=|��vz�)h�jId( ���������7ޘh���S��0�>߈ڄ�$�-]񪽲A�̒��tX�Ƹ��|���}��QS�D��u�&$�|s��ߎڹ�� Bd�&[GN\��"�C�W��Z�S��x����+C�ɳC�S��$�P3����*�<���Dj��tmFg��o��bѨ��^�s�mqdz�<���~���I�����Le/�60�NlV�@���%�0'�t<��Ye���O��n&�M���9���zS���>iyI���X�	c6*�(�tV�s��n縧���p�)�8~�/���QAR�X��=M���2�Ӌ�6h�U����vA3f��،��i��t���8����ԉ� �7�E�=��<��@�aS��}6�m�;xr��Y.g(�\�3c)o���)z��?��"]r��'u֛/��؃��*�"̆6��>׎�8�w�8��S@�Ɨ��@�Մ>��n�[l�r�*��׌� �u���5�(9_�啞9I���n6������5���%;W��Ak�?-��ͩZV�'�����Ծ�淭m�P-J0ybf|��!/<�,t�� G�Ό2&F�@�۲�]�w�`�krX���̒��/5��E-@�R{���}�wE��l�w��C�&�R,�E�Oi��� *�Oq�V��8FU,)�BH��d�q��[N]#�=��SY3�?�f6]�X4�I�e��|��۳흅D�����Iޛ�[��೗���$��š����%��x���sH��AO)NR��F�5��y{���m�dn<�f3O�6��u拱U{&y�$����\������$.;<f�2��$��k���t��a������'�_Aݏ�ir����1���r�A��� ���ȩ������o�ML���)�6Y�P�<Z��$X����0;a�O��&�?���,ޥ�^$�S��#�K�x�^�G0�_�6�p�;���Q�Q�Ӆ����M�w�ꗒ&/;4<�B�yb���Y�f�z�̠�G��E���ϯQ+�p��{�I�:�u���Hn��A@E���7�fS�r��U�Ӵ*k`x�\x�K��)e|D�����G{C�)�q�]]�0�V#�NTH�foF����Kĕ>D+�4��DX�?�ux�&O.��oa��`��,S]�ޗ�1��6~4`Ju��Հ����B:�~��a!��	D׷=�H��2�Gu/��V��Ϡ��>c��^dT�.�$��!��Z��q�S����>���Z�L�b�3?'Ҫ��='�M�!����h!UG�i�K�S����Nd�
s,���%s�k򚚦��C&����%-~8~S+�*� ��a�r�e
�@�
ӭl�,Y�~��7������
Cp�|�W-� �*0̠����ؠo���r���Me�ݺa#��{�֠dΗ�X�[\%5"K�=���:����?_��_�����v�m�It����}R�QOV��a�z����]s�*�ٓ�p�A��~�����`�hq�y��f4�'S��תtD�-�i��2�g"K'%��Ԥ��$#b0��6$\���8�	�����Fj�b� �H�"B�+���R�*�n�8�V}	8���2���a'#ADv����T���d���ϋ���.��ᾞ��:���4cB���ؽQM���1)2�����U�K�^��������	vJ�l~�s�<$I	v�%��$��ݺ�{ ��E��hF�=@<�ѐ��M�t�(�J-�O��et�X��$y1\�i��*�tZ9���&M���y��ɝ�� U��pm�	�.~6l'i����cs�ߗV����T�����f��#?����V��<io"]�t��j�i�}P	R>
�%I�oMz�����9u�$���?��L3_f���o��)�: Ј��vzv�@0[m�0V[�d�&�~�Ҵ����O�[7c���)���K��I�p���ſ�GЃf*�Ys��u�n�E�_P�6���?�4[�9�eٵwR�9B�>1{�(�.��1.6���v:�z��4�#Z��;�$�	n	��<u0_SVzq۫��q����1/u��M��7(��N/���ᦨ��Йǆdi�#c~�X�t���5	��h5~�Y�'�F������"9���i�d8��D�P�ꇮ1 wG�gd��}�bH`+�0��l��3|���J���x�4x���B�p�9��&��$��e�x�?��Mx	?�P�.5���)k|�
��~4i+�e��]*^D�< ����_=>��犍笊�ޙr�N����mu�� F3�>p�E�(zTc����j:Х�����:�lL��c�4�68��{>��?��,X�v�8Bՠ<F`�6;�����<�Ί:f�:�y�eN�QIV6��[)x�F�ZR�	�Uნ� c���t4rR�~��
����C�,E�S3Ę��h?��&��"�o��f�AX��d�?�.��-�b�x6`�B�h�����`P�/�PV�m6Ru���8��G`4���,f������Uӄ7{�{Je	M�m���K�ֲ��̒�WY�����f�$s��r:����YKy�Cw/������3&[�@�;4��?���o��R?�z+�IG!�|5P�ZiT�:"��b���A���KV���f� OKlĮ+c��_�t}��y4BDt<�qa#u�����2~Q��Ö��81��{X��������Kh �''��`Ӱ�Un��R�}�h���~MS277�"	����)h2h������Ȥu,Z��������wK�}��]�}J�7���yq��ny�œ����fFQ�$�F�Q�q2р�Ǌt�sM�p:Q�ӉM���6��,i�\��$m��4��BB��+�����v�n��.E��3���V���9�6���s.�L�ܳ�nO�'t��+�k�q�A���q^��Z������0!m��8��v1�dl������ـ���6�&2�/�l��� �Oh��qZfo+��>����(vO��'�D�<�3?e��nv�kgE�f�r�it�2Ã�A"�Pٸ���1�������U�Q=���D��<n��_��q�Ϧo*��P�Ga�\�(\�l	��"z+�x���im�.�JҐk�AP8�6����E�S*ڧ=;ԕj��͙d�-mItw��"�kI�����$����U[zo&�Y��5h��%:A,gi��
t}��n0c�6�>��֖%�]�fb:���?�U��vZ'�U\��p_��}�����d����1�)/�Y8�+�o�d��0Im�D8����i*��"��� ��BH��~�2�(u�'����V�!�X�D��ܹ� �e�r��؎�=���0�h�o�%c�ǋU�yR����!�0�X��z��Pw�<�̕�I�V�aޔh�tP��2�	����˦�v.��vV��(�(my����.O8�#R��	 P��o���cy&�����,�j�V�=��:����?B�Xw&$�������W$�&P1@%>l�˓�_u��ˎ|���2P~-^���w�k�O
fm�'v���(�`r��
Ԫ��v��|����*�����c�Z�����`�U�"N>�ҫw�s,qѝ�8Ʉ���C .lT���Eo������qt�;1���.w�_��VZ�����7��J����&p��it�/.U���(���\�h��E'���E����4��B�����O��Sj�]G`��͢���?$�d1t UO��Ү>7]�˒�e��r��N��;j#�$�����Vzٲ����1s�0]4pSA�5N �玧j+�]nC&�ߌAQ��c�#k(�3+����բ^[~�KMB�I���{�7P���Yқ� ���ZMdD�UX>=|�]>���t�e�je�\��,%�0�_�
����n�k��^��,��5捸(��(aDLđ��`i凛i���;��*�G�	���óFU��S��핦|�Y��D�Ї�p�g2�3�|�	��4VǶ�z7q$�'������(&����OQ�}Jq�#��4�a���½W�T�7�pQ#5�5W3��L�׿�?���rq��j�d��y�נ� %I[��X.���ۙ�E|��-py�2/P�����3ځ���e�
�ح$	��<��0%�����v��~�d��P2�ċ/}0`�{UDm��l�G/Ѱ��J�0�IO) n05��l|�����@�B��M_Ґ5��Y�k�7���e�-K�N��;�+>s�k��_}o�������QY��