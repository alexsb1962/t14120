��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖ{� q:4�ZH�]A�u[�����[v����hM��F1���&��؀���C��@�F�zuT��';N���c͹��3&�� W�S��oE�d�ƺ��y�ݣ.&}sn�Q�		{�4�ZuR���QsD�/�b�P!3�j3�3@,OW��7A�嚐������f*2���ȳ���-��"ݞ�������>R$�h"�IRMB���7�{?>fB��fE�Hi,���[K�
�ޫM{�j�y����9��L�x�.5g��A;\��<����=��P�`Pւؠ�u}<_� �E�*p ^
:W�$h�V��y��h��F#�u�jQ���wU.��NR^�t�#[rO���3u��"�c�N���l��vȻ ��ˋ�#3��3�J���m�F(�r`�,�S�o���oG����a��3�`�j"!��2"�Y�H^�_C�����<���{X� �����a{��J�Z�~s���uL65/��'��O���%^��U�P�~��t��P-���`�i�|��K�cEs�g<(E� �����v3k�j��?�z��0����+o��-R�1�;��?mL�_��GMI�s��Bp�5,�OB�
���%�Ѐ���.�H9WxYҲ�>�Z�3K��`N���l�IT)�q���R���Iʡ���[��]�Ɏ�����3ܠ؏t�L��w�\�O϶�`�-�����s�^���P��\����*\x1�Q��֜]o��8|6����͓�*j�A�L��c�*,`fw��Pc�!���R9��(Z(��i�7{��c�yhb�A.%\��}�����Qi��5� �Z�e�9n"�����,��h�qs$M���%$oB~㋭��S�R<�W��|�o��}r
��X ��v燻�Ρ�&3�!Y�]����wl�<�r�y��� ���9'؀��i�� � �^Kz�:��h���\xX/��>�o�����{��+YJ˕��!�Z�N�\"|^�-2�Pk�A�<|�l~�p�4�0^�%(��Ay�x�{gN�Rj[pZ����Θ-��06aŲ�X�>~c)�Q��{B��-��cU��
Hz$"sJ	, z�e �������	��n�8�<B6͸-�bqP3��?n ���S�a�[e�g����� �^i�[҈�in �+��[YL��`be�=��t��9-�0lêք�͗�P�3�>I��z�ȡ�^$<Y!�\aە,n���Bc�ė�\�I!ǆYv��ba��r)1'�Ј�����$��y��������>QR���\���~���q��(�I��� I=��~抢����q(N��{�37��I>>���
c,�~��*����N��el��8!%��lr�&����[М{�Ӵ���ٸ��s�:����{y��,����= 3�h�B/I��#��w���+C�Ԝ�e}�3S���g� ���S�a����D6OH��뢤ʟX3�~�l���\�D�����S�o�$+��c�V+��1�O����ee^���-�ӊsv�����pM{L��	�����z��n�<,i�H��2�U�eIC���%�JLo�E/�D���7Y�X����]}��-�vl���c(7��|uutSc
��r|�I|aa��r�Y�re�%4�	�
W��6����z�(B��%���0�����o�7Б�Eo�m�s�?L��t5�g�	��[e��d���/�l15J4!j_��U�����<����s��*$Ԓdt�Y�f�U�b�TKf�����@�K��US�l�d`�,���
i3��P��duppR�����4g	��W4FNd��WݤM�Y �;�v��8�������e�.^v�J���uh7�b��=���{���G�3��T�����8��%��#���rB�����N�p��iS���8�at!@Z��z�s��!��{���`��c�]AMz�9c����V+��ٲ,�:����U�es����O$Y��!�lLQ��v�c���Bz3z�/���(��Sj��� �BӤ>t^��c�}m�J$7�G�Q��{>�c>��1m��}�%lB'"��&�]�̂�]-"eܯ�G/Ck�ebU��go�ҿ`q�J�&X�[�ZbkPo���d�}��3���7J��K�s���]�E�)�a�`��\��<NRW��I�m����5�Z����6)�L�M����ߠ�"^�kۢ�D��<~AyM�����څ�$/-��-eWŒ~��_�|Z�T�cC~/�%�zKFjֶq@��� ����W� ����2��eȘydCd�2͑��SO�o��_���'W�T��d6�ln�ܸ���gc�L�YM ����-��K��[�o�q�8C�# )Ջ	�d��� ,i��Y��T���q�(��r�h��;o�ej�Oȍ�FZ
��M"O����W���~����m�<�ɂ�V�vv]�/d^�r$V��j�����v�Z�*g0a�N�[Eys��ъ���x;\�BF�5쒂�e�B��:�V�&�B;!n]��Ə�W𩃽 ^	�I�釁ӂ�9H+b�����#��x]`�u9��R��*S�^��s��ʍmJG���9�8a�������O�D#ŵ�SwP�g�av���ԍg���5,���Q񮪙����Ց%^���m �],�1B���f.?�Y��3<�X�@�B�����̏Cnw2��λ�����l8td̸��w>��}�5���������'I��jC?C�)n)j��B�I���o�DX�ר�� �87N���?�v���!���:߼�����d�MhX�N:�Fm�D�K�L�֙��el�����?a�<E0W+��K2bc��r�o�VL`*�z�L�4f�{ň�ԏm�����{�S���6�����2m@���'��NFߖ}�@��_���"��l�w�zVd�4��9$BHhʄ-4l[�� �!�&*]d�ч���e��k�j�u�t�ln���)8'^�l��\`��F�w����K����ݹ�q��K�N=�fP�� �.�路nh�� ךkH�
�-4��	�h����3s0���7�%���&�"�����N�wӒ\�L�H��p��A�UV����{�S�"�o�����Yn7D��Oc�� O-4�`h:cFi66j��NŎ��r�~y˫(]�wa:�����zy��L� ��5�%1�3�Ѧz� {�A]f�~q�)�3Ճ���p�wf#[�$"(ϛ����EO���fL��Ap�ib��0̙�0@�jVI����;����o�%?6�
�	��y��9�G�����{/���	OY�� �'TRg4�3����9����ҫ���ฌO_�]������
5�6��g_n6�F���|��6�����lA5�n?&��[?��.�UA˴5�݄��Xi'gY�����T������Q��#V��o�"��s����7}-t�^z�E��%Gi�Ѕ"��U�6 �B�EǑMCc����\E�ܥ���R�	�zN�gI������z/SO��1a�A�\Xص���(�����ޠWћ�~=K��ڭ!E��ῠ9�\�	����ֻ�m��������Ĉ*�ԏp����?�l!�+���-cv�$;)��X�y�]AE�Z,��Y��A��:���"������{���`LAl�؏)��U�9��Q͊���Y����`�gU�'�A֭���y;0mI��
?z�ـY%�V���>�?&uE,5���2?#�&��r������_h��Py��V+&