��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u���/�m��,_�v��kH&��bwH�p�ZC�P��ٙ}�.�J�@��*Eu*Uc~�ߏд���Kږ�����H�X�d���U�����f�Y�f��ts�Q 1�<p�
�Q�����n=��7�+;P���l=<v;�ߣ�:GD:+����_>j��V��o#�K�7�u��Ե��*3�iUUb�ɛ�0��?��WM��S�࿅0J��al��Z�"yl�hjtm|S#��M�oe�����Y�X�5�t�ӛ�n�W���8?����v�k-1����f+��*+�P�))��Uh^r:�l�S���TI{��3,��殂j�f�(g�j%�4\6i��Y��x��h�O�% ��>o�^ÅSÏ/�?1{=��(b�zϔ�� *k>��yd��Kn2�
�P��|YԽ������r'a%c�y�W�UQ��ԟ7� ��s#�Q��2Z�5}�v����[������_\SO��R=���],���,k��p&���F+D��l��u��ngc�N�����;�e)}Q�u������r��K˔�Ih��g��A��@�꽄P����E��iL�牫g�Ȫ�DF4bOS*�d�����J�Q��ʴ�K�KԘ6W�Cf���I�YY8�Pe�Gs����XA��ى���\��tY���i~��|YZ��r��!�����m7�bƙ{ItĠ�;b %��0�Zx�FJ%Y�
)�&)�qS���<{x��0PVی� ��)��"���6
�I2K>i�$8�<�+fF�_��Ϸ8�sm�T [HKt�#Dy�ʷ�?޽����6*2'��e�޺��y���8W��Ǹ�[� =��Jjzײ�F̔�$� c+�׫����Tw�]�cX��U0���G���zm�l�]�J�p�DХ�<a�����\�_
���gڵ�(��2h�e�i򁇉)�td{R]���l��Pa��4�@�����f ]�I��~�>�J�vf�=p�	�3K<NP���Q�JyE��^7�0}lc�v�{��)�� j�F���"h}��{���e��<�=Ns7��vF'���
��J��k1�B�,U��q�&�+�t?�aW�"����4ð������亱ZS��/�aљҜeC�嘜����PpQ-j�Wt_��2�XG�d&b�`!����V��"e
��B�2�B�����G,��񌠣⋟z�+Tb.I��ĸ�b6�2ry�23�R�A*�'���?�����	���6��2<!�0��f���hΒz^	ؤ��@d�B�il��X�!(��/�K�?�� �_/v�9����^�^��t����.��-�?p<��9u���H�
��9h���c��	�$�(p�@���|L��l����0�}��%5�B��S�����*����-���X��Ģ�F\�@ԝ����0����cmg�ڬ�(3`臆�,K�"X�>�Rw�[���Ɲ0��L^T�� ���'~�Q�*�%Ex `;�plϥt��LK��Oc;f�9�Y��	'�|j�#�W��� 7uv���W�ҰJ�+�b���4 <Os�+/� 6��6vO|f���t�^]�!����E�q��.�
`n�0Q�~��E�>��d�K)�	�%����
U��̓P��q�a�\���9@%��7�W��N���b�z�<��YVv������'�$/���m�����>�X�۸����I�	�- ���4g$$`x��\5yytzƒ��CAlB,�&��q��1�Pt���0�tX�w��>�b�K
��♜h���\�|��*�qT�?9Q�s���@���C��)H��B���1��x�T<��&�y�Tl#�� ��ϖ�H��Ԟ��{B<�S�*E��u�7H��e��V3"�lJ�щ5�@��9V��c�
E}4������T��㵣S���Њ�IZ�M���v�I:2`W)'�o8�3/��U��
Ȍa����
�O&.�Ѥt#�Rq6��Fl�#B��/#�Lg�s؏��Bp�D]W���E��$qR1]�S�u����'a�A�O����>|٢��ЂEb�j�g#d'���PB�ͭ���&́���D7��0�&c2bxA��)
�z+k�Ns�/#��b���N�W*��L��O��@�2�����U����>$��,:U��],�	�Hj���ߐhI�Nr��@FF �y�G��(��/��HH�9|]�:`�Wp���!�YZ`�ƽQ��ZsJ�ڥ��/��p3�Ͽ��e7�����NQ/����S�.�Љ����������t ��p����E�{)����]H�Dn6�t�T�T���4�&��U��3��'�u����#����8L�[�p�f�}s�{U/�T�0?^��.���c�B����M�HGL������Ia�zSj��]U�Y��V��]�AjSâ�ׅ!�dK��c�|a5��m�1i?M߸���u9Qg����@�vl�^�vjl}Gh��D�-���*�XG:8&*]���\{=�{.kT�@ֈ�[�H�b�@{�,]HH"����� n�e��'��aOQ}J_�z�Mʞ���gʼ�����#S��
��$��PkЊj>�;@�H�K"(�Z����!kFۊ���(�P�;/۝��V���=���bZ�.
4Q�5<g�?1 ��T3jV �K�@��}��X_�t�|ۖ��\O�j=:�h� ��Y-���]U?�Bv��d�!�Xv�s�鐐�	�O�
��\�M��$CJ��W!��}&�'�a��(�^�g�'�	de��n0Y,b���IR��;�G2Գ~���DΘ���f�Na0�J�l���I_�\�y������W ��{�Ɏ��y��H����94��Wk�5=z���x�g��6�8P�=���[�`��b�E̓0�$K��<���:��S�ʩ~�����%i7�TƥRW�����*xU�E�Ґ���Z�w�ދMC=�P�Pҝ�3������[8��%��ڐ����G�R�Ts�+y��{�*"�-�y�0�o4M��4�]��0Γj�9cLʕ<�L[�aU*�d�U�p���fNT1-}������ϊ��;?$����NE�n��/����z5��n��(�*Iw0����*�~�C�iҶږpv����H�����MT, �ݞ}�ڌW�]�d�n��ib�t�*φ3����ߝN��
##^/����O��-�0�@�\@�l��?���D~P��O�;B���;j0R�{��4>�>�ϘI	���XȦZ�.���c�g-�!�D����5T)Vx2�[rql7["NLkܭ��H�"�=�PS�J�,��gwU%L&�k e<i�,�i��(J