��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^��������i
��W�[� jؼ`��;�,�:X�:N'Q��������-�X6�ـ��)�p�~u���:?���f�e���/!��!�����Ƀ��l�\��N<(P�i���3��T]P~�Nަ����?�9���7�]%���^��у��tb��j�u���(�,�]�e���ީ�4*��<��9��I�[o�4�	i�����~�sjr�~���)[B �>��[m��z��w:&�o���#�p��������}ө�y���؞����:-9����ŝ��C�f��}~J_<�a��JQ>X�F�h ��$�Q��oW�n�+0��Jg�?/=HӱCi$I#	��d��>]9f ;w��n9�8�Λ*�H�Yv!��r	�t
��#�4�v'1U2�� ��Af�|�H�[A譴�fS�w��i�{a%�m�v�;#�^����xW\	ɤ%�#d���>z����d�7 ��j�1Q�g��UN㤝KU%���H,%�4$��h�X;xp�	2����5�n6A��;�u������2�(�^�˂�k�)���ڂa��i���?��+5c"��u���)��2[\h�^��Z�B�n���4��{E6���TOvV�X(����/�|��ή�~.�lJ�n����*����*�C�'&�IG։B��t�6;S�h?8��NX�V\:$O��?�����g/ePe�AZ��u�Ʈ��؏BN�t�\	0�6"�-�V�.੺	�p8<%��53�������S�!Q��_8�wOm9�TS�O73ʷ�v�|��DQ^�q���Oܔ��N�W�ֿŘ�6�,���5��p��Ye�����
�]��L2����0�Q|@������:���"=FCI�r�x'f���x�7���D�)gq��+����?p�����,���P1���r�7���NR,��:1�3���R�>>×6Z)Ɔ��;-Q���l��*���t�!����Z��3��a� K'��T��W��D���wd��!)cn)HT !��<.}�������?�X�Ι6\�/�L�Q�֤!�>_�h ޏB�]���~7X^L]7��}�	��x\�*_�F�� f��Wsdٷ
��Vi�X���T�ٲ~�s"U�����R�x�+�tCf~p��Oj��N���\�~�~:#\;"M�q��1�S������?�E)���{X�y�l���5p�n��z�ڇ��fO$�q����	ZY�YikXdqF �P<_��0j^%��2����e�Cb3p�PW�E&�O#���a�N"�1�@�(Um��	�A	�b�o��IA�<l�z�
�I�����*2� YV��߸sG��d\�g4���V灎�7=�ʦ)��o/q�jA} �-Wf���	�	�p#�Є3E�� �ضC��x�2��`�mfd>��8 �����ͩ�e�L���P+�n�^�y�L�נf� V�#d=��D0���xF���]��R��(K�Z�iKC��x(����QqW�2xZ`x�K���l��ڵ{2t+#�	`y��2鴬���H0�>�V)�h���n���׊�{,Q
�]g��L��Өqð��=��������a��*��s�B��w��1-"/� �qe�XD�te3�9e�d��34/�.Y5p�%���a$�u�53��46$��S	s�����͎�E��!�D����ҪB�r��_�ǿIE7j�c���[��b�/��������zdk�ٲ�\��W�Z��Gܬ_`������uBPs���Y�h�kXu�3��8A.�,�,��P�,�Q��4���.{^��>��<~��qA�������I�O��|�\�2&�8��;�8��~���<�*����$��Ԧ���S��z�m�N��!�A��7[.�n/�\i�q6��$0}�=
lzr�r��d�g�U��w����D���mh�=�v��3��k�/����vB�)S���v*g�+�p���D�@SM��ݷ��)G��.)�#�y�($�O����6I�v�`?���y"�ĩ��4��zFT��Sx4��Y���t�"n>�����*ݟ���Í�s���'I��\�3�b���m����������m� ˇ2��9�7�;-ᐙ��֍��#��i�Q�ǰ�"C���J���#�N����0|E���I�PC)���8#��!�A�� �y�ez���~6c���x���V�9�O(U�0{w�uw�H�fU)5��oת�3`�*��A��B�w��r�B��!�P_�˓�H��6(X���d�y3���n	��%�D]�`I�sT��o�\G?��U���*�H���W9Pn���N��{ٚt�#N�w���������4=�,��%���cOa�*���P�%a��� �8�3-��҆C%���6�S\?�k���C�f�h�Gt��ۊ7:����i�l�{��������|�s�aL���c�h^�!%)۫DA�e����.�ۿO���^�a�M?+U��Z,0IQ�D�@j��k�n-��i�J�d�� ~��s~��.Z��fF>�J��3��o���*�W�RVa�=a�v�4�7��{է4W!
a5r���\�M��S�ky���i��YU�B��ZMLf;VqR�[9���%�`a��Q�&��v�K.�&�D���\�;�4���F��V�/,1���YzM�� � 2g`l��{��GCo�AA��P�ȗC7���c�|�u���w���/k5���� R�``L������LB���"1����IHk�E��fPC$5�Ql���g��߶�D���~Ӓ�:�����1�r&�U$�au@`�� X�|�a�qH
��^��!��t���1D���ZK��k��v�	���P���P�F�i��}\��Z��p�MU��	�52� �#ꤋ^ll��Y���*��"�}�&pzn���J���rNx��i?��L>ίJ�[�d��T���ŕ��@3?�Z��o+��T��>���֪U��)x�B� aJ����=u[)�)��EF?���곦N�#�A�����������|�(�4'0th���c��%XLȹ�#��Y�c|ZT�������Jh颧��c�}�vFYϥ:GN�����UV;Pnh0�n͡'g�D[�5S�,7���K�R�1T����u�i7�Z6��v�H$c���+�p�55V�X#��[�S@���퉾��g����(�J͢S{��t�.o�}�E�����k	e�Q��@�-������ym'�P�%\KG<�t�l�H��<��`@N8:�
ėI;�N���H�������0|��Ov��aϥ��G�3>��M������V$��r�Q*���Z���0;�s���&�|y�����,�0&��ج@[^�e`�P'�����]<��֩!���^�[�Q�h=��'�Ƀ��BeRY[�'��"JJ����L�����
�<��)~�¿�؟�ۺl��0�R�۲"�^���q���8 z�p���+���'G�=�l��zf9�K��~��z���l�7z�d�Z��caɸG�!O�>����tf�w���PA
ʍS�_�m=�>��+'
v	�~������-(J?��b�9ʏ�K�ƉŸ���?��0���&�N��hG�0�e�����x�g�q��j�������~�F;���̸���QĄj�N��>�v3!��h�(FgD�ה���?��7HL��uC?܍碍�<x판"WҟY�?�v��|��$�kN��e=)�#����뙮��۱����\t�Ҷy�����t�I�)3x��E�8�-�ϴ+x���P�d�?Z]��⧔*����z֚��+brۍ*�f$0��L؟{���ب�l�:}�����5E�|  ��X��~Bm�ί�\��c�Ӳ���Z`��p�����2*#@�Ţ@}h��z�w�B��A�U�Hqt�|��TG�?1ӆ.N�_��7��m�Ό��$J9Bim�'|o"'�J&S��U�W�l"A#���n3�!�0�-5�f�#i n���#�g$�w$0�E��{ΌE4d��99� ����lF-��_7�`��a"��Xѱ�Oؓ�������Ұ��3�_�����Cq/X0Tj�.�b��QC�+0�~{́w�9=���\���̒:	Ɗ:|L���|=���Y��+c��h�:����z4�j�ʈ����j�!xB�h�?H��t� � �����cjt�1tK5���@͏f\��h3��g"��?7:AY_�]8 ���W�5�"��W�!tTuZ�y�� �|� ���ʼ*��wҶ��ae�:vdILkɨ�����Z������r�:o���:�-R�|$c�]���M�$�O�Q����oW�����|�M��-��>�Q�;���ϲ?��O��T���uLՄ~XA���&�"�W5�
Z M�v�N�\�m�?�"�� M0��_���� ?;���]#!��6$V��TA��f����»~��6`m�����?�>^�/g)���a���T��p0���Go(�M<Y!{|HP �|Gtc���6v��O+�P[}���E�(�;b�vi��Y��W�����������{�7u3R�"����Azya���Ιؘ�m<�K@s��m��r��A�C[Y�ʽ�(Y&m߆e�."��%m{
B@���=Bս�Q�ܼh޾-�0��Mpx`@�ә������o���+������h��ޡj2����+]�UB�� X�J��Z/:�I=�?2}�jql
����)z�-'���@�"㋮���}�$m����1�0���.]-(��۫I��pu��?�!�O�IZ��?ص�6
.���W�f�*Y&  ��M���$��Y!��@���ޒ�'�b��ֆ��_�Ar��B3�~"���p0�_�<���#��}@e>�άe����$�*�e�ο8�&3�:J.B�[�ky��{!�#��p��t���[�8������� �D!���)��)kD���Яb�^�f�9׀[U�	����(_���/;e jp�~��wҍ�	g� ]zXZ��%�㩧��>�}_���q��7���V����g��mW��L�bq`�����}���|e���JT�(`$���{��V(���C�,� �n�PIʹ#�"���TAѢ�	�ӚS���*F�&�mfn��Ry3�(�/h!���B?�\X��	ȸO!pp�Do�W��_T&�|������@����1�3�u!�-N��v�����~�*6&U�%$�c�5�3ѐC�$wq���S�V�nS9���NH|�[c��Y�pQ(�C䙈(2�kx1Lש�#Ք>"A`Π�1R��/5�ۭ!��[@#
m��2@���7����l�iaN�t�a�_��b��2ʝeRc��;U*����t��q �Vm��d\��Uz��6ͷ��������r��&��FH�D�-�fH�ak.��M�l0�p �#�㭖��M��NK��aOqɧ����2g�6�.-�iדOZb*�L�R1���kh`C�;]HF �p�e*�e1��b�b��S��������ߠ�t"
�Lh��4���bl�	��,�IG�n��&O�w���*V{��"�ӡ��Qgk�( �d=&z�u�J�.^\d�tJ�y'0��ú#��M�I�_UE�R��>�1��򪾶���nRvs�]S��|�7�A1��̐�uw���ܠZ�~��<��"�k�ZOt8&8�AD����ĤWu���@�YO��#YY��J�FJ� ��W//�x{fo8���&���W_^�����A_��а������'�g/OO D���(�}%l�n�vb鷕��H:L�I�����%�]��	S� ����'�"���l�r[" ��e�nu�TeW��§�����]������!g�W�k1�(,�U��ly\;���0�Y �10<Ջ�.鵑\Ɖۺ�μf�ԇٙx����s[���<	K.�� �]�d��s�Ju���\ݭ�u"_�+g�� �F	N|a�@������f���j%L��}#�l��-��6"���M��2/���Zb��M8ZR�j�Ȗ&���ю�-�J�?<RQ(�R�4`:�4JՑ=�[[
����n�ώ��t��.��dE�Mܴd4����np�:n��P������7�5c�q�W������'!�z$!���.�ѯ��g�{���"7�7�G~huO	 FŃw��${O�ăO|*vN��s�f��؇F���^	�Еj����Kۢs��Ձx��X���'ψ�tE��@��*��><�@B|:n��0�����rl�hi�9���<�+c�o��n-�<�X9�+YD�#�����z�Hվ�rc�h�m2�L]����L5Q������qQ)##���eZ�X��[<5tC�M�M	@;CJ
O��w��6�M� R/������ׂ�AP��>��"fYc�8G�.	L�[˸��<;�b��/%�SР�:�{���^�s'����*ۉM>.��uF3`/ �|�W�,��xf�y���|]����1�L0�f� ��M laSOӷ�I9%ˡb�-t�բIjV+����O�k����^��ZG��4&]���2��B9��%���^�;�?�ܽ�;��!9�ql�Eq�@��z%��k4�t���/��� X��k��c���v��i�V�w��!�Yoz3/a��}��G�e����gM������,�
D+2
`Y1i
�J�b������#��� I+/�\��VO�w~��dڢ����S�[cZ.�T����6R��%x�K̂�����$�
��|�"!|ÙPFI�{��Z~x��蹈���y�f�Vv��	D��e���76�3ɲ��s��)r�7��������e"C�j�ƣǿ��IR5���^Wn?C%�}��ؙ`efq�*�Q�����ΙkmG�~^�*�(@$W	�A��lj�F��M�.E��	H�+uG'�Cϩc�?�b~'hy.eh��YU��s0�h9H�V;<@M�x:&�b��0I�h��L�P���
��?3^�e��\gq�Nd*��U��aN芾���$5���!~{�{q:3?�.=�(OOX��V��ߣ����;���DY��
t�d�U��6:�\c���w�U��gB�e�=Y?�c��v>�:�t����:��k��:�'����v;�ԋ��ap�+�/�����Q�em&F���q��Z���� D�����t�t�5aL������*�m�M��NW�+g�_�Fw�	��'�d�&�O��}Ӧ�/@��FɽZ���Vku� �����`�2x��J@�&�{E
�R���ad؇��~`�蜢��|ǫ9�\�`����df�:T�_؞_�h���[C���V���#���	؊j�I��/:����eR���|��J���~���Z�'�L�c@0]lA#�c��/�*�Fн�oC��F�Z}5X�7����W�XDϤZ�D�ʼ`Z�h����,�f�,�"Sx*��~Pꉵ�dD�0�����o�i�F�e3��fD�l�V�-eq�k\�H=�c1�at
wNzEk��h�i�L������'��KN���I2Ia;�����W݌wY�_���%��$���'�ӎ0oWX�2�|]O@s#?+aV`��W*@{�7�~�R�/p�%Ö�s�@4��
M�5��\g�fX�VWy�EN]f���ugD�q��'ԣ�c?���_u��l��)~�
^.o1^^��bː��M�q����^6���km];����x~a�\z1��,��wWh���}�F�ь��Յ�ND�U�;Y�z�ڼ��H���8��T�7�u��R2'd�12��9�p=F�[J�����L=��r�z�?�V�t�0;I;?��~�j��r)02��