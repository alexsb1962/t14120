��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2�EH7n�[pOY@������n*���/�%Y���y��:Q
m�=�iy�W��_�!_�� �@������u9s�V��M��ˠ �4|��0�f�~o����}����z�������
�學�'�A~��.��h**��n���\#�*ɋ����;�C��U��U��f\c\m6"�m�s%;�ҋ+]>T����5��>��8L�2"��L
 �l=��
�7-؊��L&ɲ0$<��x+~\$Ϯd�t�����85����O��X0��g0M�� �m�6�ޓ�ScOS_���k�ٯ�"���4�����.NJ�6x���擱�W��Κ�9���IUn�
��Ld��4}���,�7Z^ù� �\vcW��r�C��j֕fV���d�P�B63g���L�b[���H�ۥ��I@�5���/$�%�Fߖ���L7�g���c~eh�C��73i�(���?Ŭ �<�/��Z"�!@�h�7Q&�x2VL�\��o�zxC�N��H{�;}�H�X�G�yv���N��O�����@oG"j�mr�����%g"�o ���ڸx�C�'�-���[Z�XjY/Dw/��Yt��QN�ƣ��*>:�4"No��8�����x8Wq�̹h�Ǌv��\d���.�bc���5��� �ƌĶj}_��u����t]Rt41݋�Җ:�A�,=���}=���4�����!�!zf�{T�k|J'� !>m��ә��`b�d��8ޮ�Eל%äL�\9�M;�D�db��w>���8�r#�5$<�qV]�Ƚ�7�uma���H��z�A�d��ت�� i���L y�\�WQ� ".hA�eH���Z�}�����W���*��1o�^ҷz�H
��u>�#���L�[T�9W�����!�IN|������,"�}��i3r;־��<�.�5 "M(򦺮p�8�	�<�B}�Ơ����G����P���$_^ñp�`�#,��Qu��f�<g`8�6�Q�ۦ�=MB!��DP`S�\`λz����[������* ���CX�17�*<Z�$R��\�o6]rf�ܹ6���oI��!�74U��Y�4%1��>������LL2�.�0��lO�B�C�P�&��������`<x|�d��FpU��F��C}0^�z��"\�1l��pְ�;ޞ�-�s�"d�n�	����E��H��l�x��r���^ABt�@`�X(U�Δ� %���@�j�J�D��ك�O�3B3q�+}źQ�Jz籌#��E$k_��ٍ���eu	�lm]�owF�s��]'��2+��Œ�j��N,����>0�{%:��Y��<�Nܙ@a/;:�ɣ�u�p1`�D��CeO��/?U"���9qh4R�y�������%I��a����,4K���w=9���o����Ty[pU\M�0�4(#��^��H���Os�'9�U4��<�ପ7Ȇ��85�]��ׇ�g`�BJcj�T�/��2��-,�"дC}��"��g�h/c�eE���k�vW}�"��d>� ^�f8,]�����]��-gC4ӣ�Z���u`̀|������s�FX��SacV�W� C!��YI��n&׿��k�2j�R��e��t��ϩZ�H^m��JK̃3ט+�7�Sd��Ds�8�G~�s�qR/�BU���@���k6K�������� j�Oͱ���ǡ@�s����($s1���jy�$_�QQ���<�x�LX�5�G�N(�f��r�I���0��壍�YB�_�� ld���ʘ�+�$��1ݤT#o����4�ht��lKw���ˮY�0�ʔA/IU��HZ�(�T^Dy��ꄛ��۩*���YU���~w��V!�������N�Pm�����lFbָ~��IK����c��+���?{��?θ.� �j@}K�����/���X�Wm��ќ�y��%B�m{��E�������פz���W !Bgv"��\~�G�"��H���@�59y���qHh�T�K�8�~4��zua�8:z@xތ:|�`څ�f�}�ڱd�g��o�ŝ�b�BO��+�k��Z�d���Ɋ�_a��-<�p� ����4���9/_��3�>5�r��ֈn����R��p��O�R�$�է7����mX�6%�5t���8Ht?�z��Ϣ����`�GJ��?E�c���tL׎x����=Gr^���)�v��r�ņ���n7'���5�3�1������>�jC��w���X,g�.l�]Gj���YaR&Ż�$�rO/2�ޢ�j�	�[���	p�lZ�7x,�(6OF���Va���9V��+#r{^��={1�:�Ph�LX5<��U���#fz=�2�˰�bk�x �3fҕ��b��I��ث�[��W876*Z����yA�h���*�'�<��/v{sw=QR9�/â���'�LP��KX��+̹I����u����X����N >M�w�ss�$Mږ���
����Ѹ<o�gn�����;6��C��';�V�g�C�"6�9��D˵\�#RXƹ�S�вu�����3v�x�w؇oA(w���tjS�jS�g�xt��f�`�hd�Ƿ`PO�$#V  '�I�!�#EQ@����l/��K��c���^ݛܙܛ8�J��X&TğT-��e��e����/�p[W(9����������qjb�()����/�B6X4Fb��92�n�۲L�m�b�Ef�y���s����x�o��p��,��ư�����J��$����:D���jΐ���^	r�(cVv�@�v��~�J4R�O�!
?�B�(Å�V��>��	YU ��q4?�Se~�~�yڕa�k��U�M=g�ݕ4q� <��CyVv�T!�G�W7��C�SZ�S��M�ّ��3����������o�� �9*����N� �0�o�`-�٦@���f��.��ΧQB���7o�����2�+����x1��I¡ێN��V<V���P�x��4�^�x>"a������p���N
4 &q'>K.���&��*�i؁�j���5���`Y7��d2X���\����������k�Ӡ�kW���"y��%�u^_p���l�K�N>z~�u)�e"T�ۚ�9��Я���L�Er����I��`���"�UaN����A�[�<Г0���(W_��K٨�%�Ɋ��܈Hʥ�{���,g���A��1t؎yU�n/��65�N��=j�����Dq1e�]�F�<�7��t�ﯷM��qN<�u�j;7n TA�є��G�bNΌ uVF�;�~>��]Ɛ��̫�6�X���͕F���p�����
�3k�v�Lx�����{PH�C]%�23T�q�Ɋ�R�M�$]#��Eϥ�`'j�[L���	�c_z���-�^�1�m��sިѣ�q~q(?1���I��MT��B�L|������%��D��6�K�����u�s(3�ԊlR�Z��΅oK��g�es��x��������@�}#��A�~���ܑ4�^��e��7偒Yk4ߗ0M�}#B�ur�E��_:z�>�l� �n`+�_��
�Y���(|Ij8i.�Iھ@�G�Cq�$�� ��G�"Q ��ACO$�M�W���rZ���F|��֜;�?�xB
7�r��� ���.{������U����z�'�������w�й�����4wV7��V2f2��rje��Ņ|Wc�;W��8���cOG��4�ף��n��m��;7J���Ӭ� ]��˨@(5{޶ �]����h5�C��}��
0g5�����D�H&�F~e��v��;�p`�8�u�/������q���U�y�ϫǤΡ-Lz���e�%700I�VF��_�ړ
ĸM%5 �W/������]�<W"m3{G�����Ig��88/�#�83ƃ)�д� ��+IJYh��m� �J�u��!���_7F�=ǽN$d{i$�uo�H/���i�����0�^���сDA�{��-�D�<�^1�EV�`�9鎄�}�2tf>'S���
!e�;����9Tp$I	I+XQ��|ѶfHp~}aE�#�#	J�j,&�<z&5>��Gc�>��.�^���ee��hT[���ώ'xo��u��7�A���%8�/���=�:��7򄰦�F����� E�[#�Ӡ���6�0��.#cZ�z���k��� ����s��tQq��!����n�x�ƁC�V���y�°��i��������x�X�;8��B�P*�
��tNqPy3]78���^����1:V��h;$X��-m^�a�ߐ{ڪ%&V�8�)��ԩꎴ��~x�4axd�#5�U5X 1je�Sa��C��ڛ(��)��4*G��&Z%��_UϬ�f��g���=uu�U,�\U��+9���_�c�[P>[���B����&�j�9`��o�^���O+�&hDK�!��M�MY?�ưf�qg�CGQl4j�8�(�XE&�Ȍ��>��s䷛�n�<,Я�n��H����� ���'�`Ľ�V4+jC�� ��"�?)P�I�:�q�D�<����B,9�z�9"ܲ���z%�y��<��ܲ�wB}���7�9���p���xFp�;QQ�ze����4���#��x��8���5��Υ��	NO3�ߛ���z������f���q��V�H�p|��}���V���[#	��'�Ѽ�6Tn��;�CG��g�ǂm��{+� .�\�%�S�^cX��@�?�6�ۚ�Mz]�PǾ����2Y�Jq6�k����ބ�D���^L��9{gu4}/��x�~M��D`%�������2��`�haN@���Ft"Á��M���0�MS��'��?�L��{�ǻQ�d�_�6d����t`�١�`H�1��
�N$-wCϵ��=yW�|�(�l-��=ơ��s�A���vNB/u�v��e@o���|�DB�$	Mr5Œv��s#�n/!ŕOEu�v�� ݕ��T&�h��%�(�mן��{n����O��I~z��
2�a����S7*%.�����.� �:���2D�Wt�Ut��<C���LW��@5'I������/��;�������H`=�b��uu���(�����՝��JsCl��G��緔�l�}z@�9�Ȣ5���`��~����Q9I_bW�bh��l���j�ŞF,���y��]ֹw�ѥ�	�Zyю"T~u����-�%'5��Ѧ���8�8T�~��eW;��/�����yo�|��jD�q(��p����0���-��9R�����%�s�0�Y0�Z�_`�|2j�L:7�s�5��ٻE7E&�������Ou�����QNm�y(K�����.�]a�X|R*%*Ë2U�։��on(O_"���TQ��<������n4�/u
gzg}GG�C@�c�#�ĩ�(DxϪ�QXC�ϻ�g�R�{�ȣ�'�Wg��	dWL��P�*��H�!oa���Ļ^*D/�RC�7s�єqL�!�Q1"��	���F]�Ρ�������9�i�ܹ�J�дjp��µS>���.|t����0��k~,���x�o	�F���"]kz^����/��p:����qI6���\[C�n�wq;}�)��Bó���D�
Y�O��h`�l��
���5�o'+tFu�{ ����TLZ$�`��r���5�o׵��T*�ܶw�mV�[bW-H(�F�]��W����8M����1�F��NVRR$�:M-r��MM�,�;��X�e�H��a*�aĤ�	��<�/fCghs�T�0�Z[�(^ӚT��Qсܼ���0��Ǵ�+y�ʕ��X��<�+�����ÿ́]�l��nѣ+�V����,l��e�xvgP�"���HM�t�Ē ��$n�Řu��K+z�?t%�t��Q�ȟ�Yy��_����x�
�(@��?oL����`�N�ER��6����x�+�*���J���Z�;�x�L�Ew��Ґ?�{b�hZ�UåF�;�V���\ߘϗ8��X�QhvG�81�?Hx�	�z�n�i�Xp�1�@uʍ�ͣK��2�<�N�]�j�׍{��s�q I�i�>}:�p�l"n^2�'V�Ә�M�j�1}Y�O1�I/)q�9(簄��v���=�A�� ��<i�D�$��