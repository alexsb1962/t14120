��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ��N������N���^������A�&�et����tχ�Ј����	i�ʍ�pN���-*�4Pn�M�7��m_���gG��R����(��m���O�E���=t�)l�������Tb���Uw����<�]ųy���>呕X�<7�6^��11�a�
���ȣ
���Y8�?��3m�)3l�V�f�2.��H�J�)��{^1MX U�3�Ϡ�R���o�ǛH��R��@��)+Y[�	�\������+A��Y>[HD��i_�\�Wf�g_�΁{�д�9���5g�P�q�j��쾓���P�ysb��S�B�C���)о���cr��.$�
]E���O&�6N��q�x-�׸���a�	���S��!,�o�1����[��YNH {������34���n5<�|��Ӫ*�������0��eŹ��Y�0�]�Y �-Њ�ZR���t`����V�p�s�_����ڲq�ش5��h�CN[Ri�Yӓ�t8�N�E�G��Shz1�&r���#���w��&-IJ����53�����ϭ)Ψ��c+DՊ�x�����a�B�TTȑ��8�Y�ghmr1Ekv�$!������>�^��Q�	H�n#w��S�ܷ�õ������+�,�p�c*��0(��qlK;OYc���q���"-+��]x$�@��jR�_��7܄�ӝ#I�k򅈮1E_�w^H��jx+�4�����_�/S����4���N�0���[�V8r���Iq%&D�����t]ŽJB�j�+`۹�̅ᤄ VT��.���n�:��?E�Y��H��C�'&S�K�tK`l���o9E.!o1o;8Y����
���z"1bh]������z�Y94�ǧHO9�?�C�]�
D
�1@�XIk�h��d6Ԏ�.̩��Q�8E��x.]���o=v���ZC���W�s�:Bg�[.�$l]j�Ѹ�I��,G��r�rA˭�6��.��@�4�g"srz�/yTڰכ�W���`Y�I[׈�4��~a��~+�U)�<�������ʘ� p��(X}k�5X�2�H���TR���y(�O}⒆�:ɍ��J�Sd� �Q�ƇKd���B�	��R��U�çC9��:������J�́\ �f��S����
�6�i���"�ˣ�"�����L��*9�I��px�Dh_��z�o���68���3������S��(d]L��O@���D�+�~�����B	�-ov���|��M	K�W�$�|t_g�&���A1�kl�ܝ��ʭM����$� ��\��[�N�&\�2�]=MLEV��8�^BD("�ٶ�������f�F
��]ˤ���U�)�Z_ה���O�ߣ��(Ҝtm�ki�)v��Z����������H���\�@�@��R�wX֗5X�������k�F`#��s�,�h)6�F�s�id��%^��1�f3N�7�zO-��)n��N��B0�8Ց�n7�]pݱ뙇A>ی^R��٨:����Ǜ>�5us����K,EY%r��wZc_���݊T �|��G�Dl� �tL���^�k�(��I�̄��+wQJ��BeX��,�p�Q[d�5VԻ�#�p��g��]S�K��4����N&��[�``��f7����T�Pg���O�P��h�*rQgε� O�N0��؃'�޸���(�i��?�؅m��n� Go�\���0�B7�;�t-�oֶU���*�!],_��u��U�fUF��3�wQ���*�G�@��dl��j<R����J�Fމ�-��^�&G�]Fs�����ï&'��
��������Z� ����霩��p���+r6�� �K����de5�:���Ԣ�!�u|�n��}�X������n6�[�Yγ�ޑW����H?��8Gj�
Ҧn��1��m�����&�g�\qra�q5c����}�
���lھ�x�{�9�I\��{Q�±�����`�J����v%I�@�p�n
1`C�
��n�I��~Of[�����{P�]��,t)&�,�Y�ko���7w@�l�R�y4u�U��i��`-�$�:���]|J��pC!��wǈ���x���}��$,�T}��yj�J�72^�_��Z��%�P�zҊ���(�i�f�-.��˘��7��'�Ɲ�n�Y��Ov5K�R�@B���G?�f;��LX  �0��^����+B�Xv�O��?d�ܵ�V�/�na��sEk������e�U]nWZJA��4$�d�p/�<�����ƍI	�5�
i� Ȣ�;gv�D�l�ڔGW�"|�lWz���v��`�����g�`e�+Xf.7�m,�|{�4@p
��`��Z�$C�a�L82�4Q≝n����Ž1�i�͐X
�/+�Dge�l�@7�i�"��uu���p��̥�O����^�`�Q�l8X"&�'3�-����'<�0�)Y�Oi6�%�?}m.�^��#�$�8�������x}�K�6��)tI�<�_�c97b��sQ��܁���۾�ݲ��&x���CV��,j�h2Z�d��������)O�}���$�z]*�H똋�O�P�8�d�`��Y<>���7�iQ�R�ܲ�>���ȝ� 8�"���-�0��Wʉ����U�t�+��
�V��C����DW{���Ώ�l/ԕw��pTk�\%�7��f�y	��䷋���T��)$��B�!1���T ']4.s�(��Z$�7��*�c�@��%f�[[����²����C�D=`	������ְ�^l���k������_cvHoҘ�\mi�ȑ��;O�iҊ�EB�ٝ�@�-Pv���qwLʍ�G�$h���e�6R~$|Dr��[��7��S*�[u6�k��p�y^G�ʩ=������m􊈪�пa��>� ��а�c~q��i������uyg��D���� bȗҭ�TB�1r�j:T, G�UH�?=8��hƤWh�������G�)(&�ef��⨃J�I��aឝHn�sx��`��L~sK]� ?X��-l�O��c"����QDr�(�纂(��z1c��E���8��:�֛V�`C��������{v�H�Ǣ�����pݤ鼧��a{�HW���/���ёhz"R�|��I"*3G�����X����B&���a��͞����� �F�8e����#Oul�b�T�$D�T����\�]p��:.���,�VGP�߈7uV��`+G�oǼDS�>v�hm���6o���S�T��n���K���r�f����Q'Ɉ�uJG��|��`+��Ӕ��x��\x��jt���g�[C�_H��� �w6q�>޵Vh�f=�^�������!�~y���B�VJ2ڊ)���r�� �N�\���D�?vf�ȫn�>p�}�i2�)�
�<�ɣ�nu��;�v�w�a9u�2D&�~�� Z,�=[�>�	��&u��&�r+`a�������Q@S/k��!�r��M�u+�+n����%�n�GN
T�  ���%'�R<q��&r��B�C�F��[�Ӯ�*�$�!9�iVS�M�ñ2��S�'|��^�i�
�Ȅ5�_����7F��f���I��a��UI(�:�t� �HČq�95�i'�-��d��r�U!����P�Ϯ/{Ẓ{�4,�'P�^
�Q�8�*����z�:��w҉��)156n���|��Wr�t���X���Vt�x��fHWYc5�s�"�0�-!���T5���a��$s�Q���(����`�Z�2%T����zi��;��Ś�)�A�.�k��a�*{�X,�i��������>��(���Zǫ���c�x�T�;$�PY>���M>=�y��Λ#��ãF�%�7W��� ����-JS��<<�
�s�ݙ�䂳pڜ��-WJ#~	�.j�!	���?~�(b�j�N�;����Y0!e:��ڦ�{�o��f�v�G�����j�fr!G��ś��K?Y@��sd��>��pʴ�J"�9��hU%�~tv�F�I����;E{څ�>c>�>m����u�'�Еb=\Wl���_o}��ƃ�b����L=��$7��U��~�p^�>�bw���r��\'�,�
�}�n�s�?y�FG�G��WV�I���&���F%ǻ�NS]���.(�M�:shC�����^VfS���� �b��؎�ic�q������
f�{,�n�B�PBt ��vO|�hKTi�$�v�Y�ɹ�}Fh�5J�d&�v�荘�!ƈ!��6?bC=����UT��\�J���ȍz-�}PZ�z��7d�|HXkv��w�Lmo3���~-���֝|T�X���xl}ڼ�ˋ�&Q�P��Yoܚ/��\��J;�P�pF������x����^�������Szĳ@8T]vq�C(_�ʾ%�燙Y
�Y���׆z&G:�+Fkմ��\1A<�i�7ضWO̕?�y.h7�~wl��ⳇ����H�6!�Y�����N�����^L��*P��aʪ��� 1��P68��|=�I�w�iS}��;Ul�ACb-��)���u3�@�H+Mڗ,�����f�����O_$�{m1�w�[������tN�(�A���HR��;-�9 ���Ӣ�j댓K��6��"�P�m._I �����t��;Ic$R��R�V�V~a�|5�t��w�t�=���`ILN�\�$4Im��I�2o��yh�3�+���y��- 䇟-#���������L3N]��)��"��K� �� L�z8�}(�c;Jc��"��e.��.��2��4&;wR�C{竣�R�g�:�
&bl�҈K��X�ϨSfF�-�΅���5�>���b7�>9?Ն5���{�"fD�O�9�ŝH��LIfUi�}��F4ii��=v�0��YIY#��'��~��D*)���T�k��s{�BH:X[���e\�'�]1E,�S��z��i�?��[��jlZ��b��k'���? �q�=��P���)ބ卖\�c)/��p�"eX�Mƺh��3wy��+;ɳ��h|�mM�����=$,���BQd���a�1��S'������%��� ۟$�}l�[�b�w��<��T^�xQ�Vn��u u{�rjw�:�R_F��#d�\�YDR�$dc��4þN�5�E�ډ�Le�y �W��f.._q]�$_xL�1�nQ�o�7�F2����׊&�AS{�7�(l{�L�҅�tH�e���;V�W#-ݳ�)Q�+y�I���<�kl��ڤ�������^��Y> J�V�O�cI~��-]�4G��܆b�;�޿�m��$���`� le����A�IܸS��� ����yy�����V������R�E&Iޞe�8O��VyFZ��@^��
��	�NQ`ş ��\�Ĭx_�w�#Q&�fl�r1�S�i���Z���c�U�]�6$C&ܖ�k/	�8�1d�&�v/W�u_���Bx���q��,@�[5K��lj]$�ZZb׈Ns���?�������֓e�=/�����c�2r�b����D��2�9�(�����{�n|¯�E��n}���煏������-��qj��Ӓ������ì�]���&������EX�7�W���ks�͟M�9|�:���]�T�b�m�_
ߋ��ĥ���D_/`o�D%�m]G׻�԰0�f�ٖ?ƞ0�#�ª��bWm��57 �ԾҰ����N�UB5{��Si��6a��?��R�¢�[�c]X;�QA��Ysu(lq֌*U}P\�ml"9�q�G��K���ȑ�� ��2�$�)�B��� X!�fgȜ`v`���q�dr��۲�`3|�tw�l4�����$��F��>?������&f����c8ͺH�J��X�^zkLm�t��М׬���{�j�?ڣ0d��Lh����`W2|i�Ӵ��A��Th�ە��� �1�e .倠Ylhhn�0ᐙ��G�^� ��M�1DSҚa;�����mq���'��}��8������Qtg�����=����ZːWb���w�iK�pGK֩��Zi�=L1� (#({6��:!=�Ŏ�~��w���îv6E@�^�ٴI��^���\jh����5�Ƞ (��Ι���Vw^�.H��a�`�:�GF��ƀfΙs�&,�MJA�>��e���_�o6n���:�b�Bt���Ӎٍ�
�W]l[*�� ���� ����j���ŧ�ah���sj)��?�@ �?�g/4H�Bvy��u���A�X���d�i,Wc�"��+W7gMq��e"�?��I�BY"O�1�?�q�P�/��$ʝ���ӦBCۆe[��(����[��%6ɨ���6+����	}��+���S4+��O�m����$��P�s)�dX������<Dh;��Ay=��=^��ҧ;��R���sm��/����NO�=p�Sc'�R|�:j�w¹��,�ף�S߸�Y�M��V|=�ogd��<ƴ�λ���w1|e��y�_b�(�;��=��&���x'��x۬�>5�#{j��<���ځ��ǘ.=��+�4����@:1'j�9؃ZVE�nƋ�K~ȗZ'�o5�*��G��]�5�~
�#���V�R* >���2�d��e��m�r�Q��F�ޚ=��s�݃�DnX[��HR� ��Ν㡟��4L���T�6������ﮜ[R͗?�*yM����)$E�@j��7�~-���hg�O��kd���F���"��"@oF�\����W2�C����"�
���#C���Eyנ�Z+]?�9�N��z����䝔��Ӝ��N�;BT�0�"NW�'ʮb	�
�U��jB
ݦ+��a�t�R_���Ir%�P��o��|xl�%��9���#Wyˑ�4hbi��4@?��ΗC�#�p�c/N�'D��eWh60y��G��D���k��+����Uk�B��0�X�q<�iL[㯯���h�x.�Kw���+D��B���c��4��m1z�6����.~�/�nm�3��a�Ja���ϗW���ڢҌ_�R=���Yic���h2�[���K�'Y�T>�������X{��%��+����[��C�T��Y���gDJ�K�zt�k]��B���=�o������Q��q2&���wY�x3z�-�p�GC5&K��Oϳ����C��e���N�j;�p��^��{�j��ƅ�U����e`5s���X
ߓR��Qvd�P�����)&�l�yX��=fY2���KC�k�'����g�?AQ9NAQ[����8ok�ɕ�N`�9>uR^����B!> )�2�(sl���S٪�{T���m����G�C�@��7�C%`�9����y�50xua���@Ʈ7�8����W�#/�"p3�;B����h�8��R��-�<�N��2T��R%r΅��8_�{���xx�.]f 2��4���OQ�FIe���p�qvXm���?�;翁��m1a?2���Qm�0���G҆���!X��5xẔ�<���U	���s��!)p�� ��4xdW|V�k�W����i�}�A"��Y�:_uf��\��2!�CW 5 w��7�l����	-���\
S$ �}q�*��ӗ4��h>\~��UC��&����C�2���5H3f�4�]��ߢcUα�֭V��^��x�k