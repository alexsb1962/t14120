��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:��������uA��@��y���<����xDET>��W�����C%�=U����3v���hj��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`I{*���:�S8����m�InLK�q.O��Mv�I�Z�*��Yi4v{C��%q�=�bL�Aoze:��
�0��`ƅ���<.�W:ay���U�&Q��F��,U�.LZeW���Ut�:�t9X�����x�{ �*����ڲv�S�����&�]�=��cڎ�(ژ8I�I.����$�K����{n��~�Uoyp]d_%��:���憐'��KPx�����f+��p� }#:�燇�@Z�h�4h�v����������h챁�������Ib��� ��g��ZvՠBksVrڧB��l�,5ܶ��h��Q'2�0�Zh�G���� ��r�}��a�y�� ����)?&-RH��Z)\������#L�F�F���N�F��b�k8����N�Ŕ�ö��Db�ÇJ9@P��PC3���kЈ���XۿS\���%ɴ���`+���E�$�	Q��5��2��G�[`�[ۺ��D!ݫ��?0.[��J"'�Rl#W�Sv?~h��ז*a�5�%t2�/�*��$��s@Ĭ����-&�M&�|q��pw��-���
�ya�/�;�<9hDS��Vg�Y�X2_Q7s���֡NhYп
��ٛ��4F�1-���f1����_�I�I�)�2�����٪��BwU���`�!A�Et�dy���ҹ�e����y)|�����DB��q��e����L'��Wĸ*�6��-�����/4�J�t�=��dH��b�d�_U����	�L:���[����q���O� ~m���x�Q�+E������{+T'g�(�6�x���Ki1��T�L�����7s�,u�G*=�M��܌7���L���n�� l1�۶�!�z�)�c��dF�ұɮJ�g���@��n�f �4�K/��JZ���y�%E����ś� Ғ+p3Zx�$�7RxL#�����H�m;�����X/������ ��uu���U ����J:#�I�������Sˉ;��w���7��!�@>ͥ�/� 1����*�?JWOoR��Wґ$���{/��D8RT����� ���֨��: ���������݂D �����)������iO��2jG�'���6����H�-ٱ��2�7�3�jw����n�	R��̍����}\k	�r*�� +��7��ѺFE�V4d�U��T.+�T��v#�%բ�m
w=���/i ��X�Z�����`�x�@�[Ԩ�sS���� ����{�//�\��_wD�S���K��ʮ
|5&|�ܝ˒���tLؒFo�D���EU�������s����INb��:R�L	�f������RC}7��յ�r�{j58�ʹ����J�mr������,�˷Oh�i��c����W��؂0�#[F=���B��t�ۇ� ad��}�ad�Ŧ�x���{3r�P{r� �6r��j�帰SQ?�>|Ȱ��h!�D�L< F��>od_�!��	_x�闓s8�٩�Ev�gw=��!���B���GEk��Z��D��)}6�q�����A��l��2�S;^�����X�Cq�@���78]3H�r�|����Y���_�������*N;_aEf�����_f��$oN1�;�S�L���H��j�$ӛu���KU��O�C_����lʘj��=<47%����>T}���:�|*x�$���.õT�c#:H;�w�,��;b6�,yٜ?P��|��.���$ �VN�F�,�&���[�s���~�\��"�/� j3A3�M5��Rw�/$Ħ�W�D��EO�6��D����gÐ��J�����*��y(�wj4K2��kN���K���XEl'�$�+F�����;(Z��Z0��=n)ޔ�l�3Ǡ�*�h���b@]H��>�:V|	��OA��)n
fK����[�N�� ���#~N�9>�dx��Yu��&��J$�yW�rOm=���elb��� 
�S�L�Lw��ir9�M��$(�����p~����������#YKhr���>�"�-���a�s�@��{�9�2�8d���T���;��1���i1򻬱�7�[�K�J�
��<>��г��_��/!yst��h�=���X{�p���3� v��X�֗����j�N�c��n��#я����>K�WS�j����Z�����I/��N%�o�H��wk]��Aj^y���^�z�JR0�<��c&*�;�Kd�nOb>�(,���3͌-+����u�(�w���(,/	~�e�0ػ�<s��a��#(�_'�'���u����K�!<��J�a�m��Y�յ�B��-�G�0��!q���1��&�DF�X��	"�0���G�nN��Ӕ��ű��o����W�m 
��~�z����9	�_bU9?��w��]\���'6�
l����؆��m���k�.������-�+�X�~7@�O��ѤI!�@�,�a}�Э>����!⋼�,�K~�̩v��;`�ie#0q����b�3I�8�zBTR�]vI��I�Ĭ$�<�z~e<.��&�	�V�Q ����G.����/[�����Ժ���ζ�>N��c�g�39`���·;g�/#��P2Q�;4������[/i/�ޮa�ķk,�jd��9{/��J+�j\�΍�8����$l�!����͜�J��j��ݪݷ�a������?#P�c[ s�t~�k���9�	��#�B��n���|^�]�瑉w>�!}m[>d��s�܈�9���9�v�*��1���z�%����a����^n� ���h����H�-\��4/����ɚ��Szu�y�a�#6�O׃� `F�5�>&�Y{�1~�^c�T�-�w\C��P���U]�r}�>r�z��ѯ��$�W�1+ܟ
��쌳'�x����I�mϣ��J��ׄ��G��J�$t/���>�R�`�/DXX��>��:�t�Pk��F8�D>�Zۯ�ۻ~i`�$�s^[	�ŇUn��^���<z�.M;��1��������j�g�����!n��.5���+�U޺f���7�l�Y���t��*�i<�-�=��w-��Ǌ�>A)
���%���}�8Z��nz��^��;m��Ӈ9��xlJ��&P��'�7���Q�d�Z��v:K�����x��6kxE��$ٱk£��wpv�us��`������"N��2����l�[�l44Phb��N�E�a�K�>�s��FQ�\ʘ3]9�OV�{�8G��v��6����V��M�磪�z����I�g�x���dz������-ZF~�b�6�7v�{`�+�<�FNH�E/&��v���Y@�:���x��[9q���py�̈́XV�T͉�E���^�`Iq�G�PڧY]�x�3���Ҭ!+�cn+Ɣ鱧��E�^ፚ��u����Ho�sa�ZTJ��6�`��(����݉������ɑ��p�p�! @�4P��r`�uu���w�I�L�C}�,k����TZpY�?]�1���~�!�8C9��J�`'wd6��ȏ;�b!���Uh��z�Q��A����U<Q���f�����8Nͻ���\�D/[��!��&v�TxFl�F��'����l~7~�9��7��I�Kd���ȿ61SO�s����=�)|"@��(a]����}�*񷚀�6���7�1�X�]���:
��AmmY�/���#����@��ٛnr%ȘP26��0桾4|]Ԯ1�I3�ZbNi!0����4��M~~U�-��*H���5<������eD?.Ej��c��r���y��ǁK?M֕dw�-���v�{�ŉq�@����&�<`�Zd85PW��]:������J<�����S�����2�
m�a2%�i�\��yY���n��gZ'*�曱|�coĢ�ѭ��s�w�J�WҒ�hX~�=�-�{AI.��E���Q׹���C,�m��N���Ω�~��k8�5�����o��_1+�q�#��5I���b�)[9���f��[�����d���*DI�����`���4~c&����~L݂�$���p�B!�h#���L�v;T��O�O	8��"v��r��0�ho���[�dV��9l�`RJQު��,�� ���#Wgf���-@��Z?O���*�)T��~�D��	R +��$�]�Bv#�Ϻ7���K8Sĵ�Ki�<4��V"�A�6�%�^hMY�xG�a~$� �;Z�q�P�f��[Z3.Z{d����+- ���{��N�v��m听����z2>�r�h٘g��auL�_Vת=��$d�o�8�T�j�i�Q��_i�*�Ǐ૜&���KG���8r�����"�~��M+b�"lT�--�Q$�%�2n@�3Mb�|��{�꽵1�#o]jcI�*��ꮝp�_� fӖwn��T��`?�}������@5�~`�6D�{E'�P��گ.Ĝ}��wr͝��!�/��YZ��p�s��/i�E^v/��\�p�C�+A��|/�1��й���.� "��fRLZCVI\c�K%���tF�ҽ��������'�f�뮢�����LwTf��F� @tMZH��k���|\sC+E�骝^�t@�À�3�����+�7`�?��A�G鵀< �� �z"�K�P�b�Wc
p�I�X�BS*���M-��H�h��9ϱp�J-�95�]�:4�
ž���~��=im�f�p�_#-t�_�%y���Ό�>耈�C_�Bɻ��>D��/��S��q�Q\�;֚�5�d@Le�����m��i�R:�PZ��;�޾><��&�L)X�����/ �f��H5ڢ�
v�yO|�O���&�;v�K���DG��<��p	�ݎDW��s�)D�ˍ�4�
sAU9�3F�~���@�?��?̙Je�Y�Z��M� ���5�Q�5Ǐ(1f��������a��44�)�8��ѮqS-֬�,	�ȴ����k�V���q��P��u�W	)�6�$��ޮ�vl��g�q�=%�Z~M=��u��J���o�r����X�=sί������f����s��
�c؁&��&�Ӵ���x�i�ݢG~��3�=��+q����!�m5�$;b��i�%[(�iU9�'?��n6K�Սq�y�����"x.|>0��E������,��Z���ױ����+j�a� pF�K[70'���#�I@|;� ����U�r<z
~01^��)Mj/L��ៃȣ��ߵ,6��&h���Eٺ���CT�W�7�k�%^s�5;��^ʙ}�}��U`� ��dMԄ�r��o�{�RmY4Q�װ�Q���s�)=����ٰ�B�<�2\�6����k�Z͈��9YP'�t���U�9��g/���<��3d����G�2��EWz�%�z��{���m
E�������$S��བྷc�9�;���4~�V���rq�e|(��ȫ���23+� `ǼHۭ��= �%L�{yk���3(�^��}3�����6o�`xD̯�o��Cb���ϥӓ�z��I$>�l�Yѿ�� ;�/�m(�H�w���O)z?Zo!t� �4o�`���X1��z b`v�Ϭ�ݖ1O�T��6N%ķ���-jo5F���'G���#>����,5W����x�1%_#���\�j����D�-���Xҷ=��J�������K2�ζ1w�9��ө8�9K�>�ߪt5Ѧ?�H?���ffg�-a�W��+�a�ׄ�)*U%�r���J6wv��H�Q�������D��%�Ec�޲���Y �ѷ����$��tp�?�x�OX�3a�ȧ8�p"N�*��k=��$³�aEz�E�� v����z��H	n��s=|�H�H,�lȇFl�m��A�O��� ���D�<ݻE���1[ku��0揘n���w�b�w#���\��nΛ��	xD��֬��=�T�m�މ5+�6���
���3�ĥCՊ�R��0 ���A��
�����[9$9Y���z��^��/7��f+��%��K�|���8D��ģ�����Y�Lcd��\>J�ti�&T��t��۫J0D5U�I3���Zp�B�l8#��P$�xm�����I��O�� �
ݸ�!��EP�D��D�f:�	
�?&?���]���y�x��.���ljbҚ�y%4�I��Q�$=�5VJf��6̚=��Qб��h(T��k
Lbۣ	�!�Q$�ܠ@�Q؃"X�!5C��㩻���>}�Q�ʝ�O��3�w�j�*W�AMuH�Hw"6o��z���¾�����L�_^L@����~'r�Ҏq�T�ߛu�bt6�����Y5i�g�����Oo.���m#��|�v���ҁ�� ��U�s�;]�L��Y})Z��nY���:8�+j�]���Fi�%y�P&#��@�l�R�h��ܷ�Ӭ�dɛ9O�-d�"�hE�t��'��-�v��2}��Y�g��|��*������U0�H�%�P�Ħ��4TA���y��XW����{�8i��rE[�V��&r�4�W�?�EM�0�_�갞�3'R�r�ei�j�e����?p�UԖtġ�:��}	�>v���qvH2�;������^:,�Zr
-�@X�_�7��y��9�(޽!�r	е�T�@n�v7n�w)m6͐5�g1�a����Z�w.���[O�/�j#O��*50��m�0ņ��Ȳ�ں-��y!o��܎��z�O���I`�~�(�t�^ �*��I��pD�#b�Wb�q4X��Y��l�����C$k���s�ن�S�Ļ&.�m�2h���9j��q}���z�9E�� +t�`�g�G��h��ҧ+�^����GvL/�ZV���]�*�uI�������+e�9��zZ1�ͅ��p�E�b�^
i�Q�`��v��O�yT�9��_]x
ėd�/N�ʪRZ&�GJw;�>�<��&����bf�%c0�!��M���*�Ş���v�u�:����=0�	ϸ$n���i�nõ�w�s�JK?`K�-ݴ���Hՙ��`�d���aG�����KZuQ�$��a�<(�������'�H���풅'e	�H\�R���ހ�Wf_k��=��[>n��ϳZ9݂U�a�hΛ�q�4�,Z�"Uy�Y�8��Y����Ķ�e����˸�T\FG�"Sd+HH�-���Sô)��5)W������D@?�w��#4�C�	j4q�[�0��>8�X��1�*4߂�����t����2�}~ڋ����ԓӓ��{����d||r �e'���b�J9s�|�W`ya%�W�%cA��9�aǽ�	S��r�����|6���qka�8���~�3vo"{j.$���Ob]qP}�˲�[�\9dM��/��s^�v�q>}я���u�2YOc�K�#�����o��:ޕ����mB+[��Y�W�؎\Ƶj�F�x����℠8�՗�zԼ�����9N^�#w�k{��!Z���8�����Ǒ}lKS�>�j�=96]^и��a�'����Q��5��ܡ �PP0`�T���aL++�#�ö��Ҧߚ�$5y̐a�wA�p�%i�1�a��������h����o�$Pq�p�PI1����t	��={'��cH��6�WH�;X�rA]�D��vX���a�!��1�}OY*�j:J�����ȿ<�!�[���YC��[2i�ΙS�&��n�mA|k}eM�K.�����	{��V�0�1�V~
a��}̄H �=S'��א:�`T���cF����8V��e�!4CqՍ��=�f��t
�������Vty���5�?u�v@j��G"+3�<oI����a{f���]А�9����\$���f�P��=�a=.2h�^��2��yk�|ZK��LsFW�N�u��X��� h�5����Dj���S�����޽����72�C�x�e5��Z.E��1p�C�"R��:b8�۩A��atqo�SQ;�D^�y�,�B�&�	�)q3��Y)Q��uf+gp�W����uNӬ� ��IQ[A&M�p�K_��j����QO�'�_
������C�%�a(�x2�JL��W%��8�����5�C�A�K�)��nwj��u�|���VM%"�j ߸L&�;2I�_g�<��c8c���T�)�>&��������!yUh� �ƹY����z^yFM!����n^f3�{�^�C�B���?��!V��A�r�Ծ��sc��q�a}e��H[Tx�ǖ��.���Iin����ņ�Gj[�">w�x(��q��J�ݼ��w�|o©��[��ޫ&���(B2��f��W�S絪(YR]��	���T/�n�^iO�y��w�ŀ���ޡ�)C�b�ƹ�JR�QY���Z���Tb���}��π^y�O��oۺ��9/z��?T����v����,/^�C6F_Ki�4*4J���3�9���8��1�o���+Tc�N������cS���=+�JnS��.�-=�2|�2�� ���^J �W����o�hTǔ��6P��^\)�Ϟ�.s��ڎđ��(u��q�v�}]�WR8��i�P�V�ض� �M�yN&���i��|�U*;q�\bϝ�kF>)����ͶW�hf'�L*��a�z�����!zϏNP�2xx~6C�������0B.�(�G�yq���L1��zj�{��Om�Fsc= �f�Ch|{`�Σ��r0ƒ��٠S�g�S��,�v�^%��GJ�1���J�����$3�Y�U�����r���4��'�7�	Ϭ����z#���N��/��A���J$,���l���	��M�\����[m���k3j����!ܽ�G�������쉄݀�|]�@�(4�̍P�BR��x�����?��F��Bhd�,"�����x��C.����Ll���JB��j���)�u>ҩ	W�yӯ���6�!i1%��M�����zE�˻����r1>e�qZ�Y)O�y)}V��_�V� ����i��[j5M��no��$AHgf��D/u.�2��r#���b�Wf3���n�e���������'��o%�4�S@����"򯬟���g���ʒ\�B�%�Z� �ƈ�΁���ۀ�@��S��@=��h��/k'7lz�׮�P��w�b\��Nk{2)���-�-E��̽_A�F�X#���`�c8��O ���G��é6�_���!�^^#��v_��t9�}v4�)ܝ�HG������	Eq�P�mh���נE����C&r�C6C6�&��"�`�4�����U��v�jK�۩�)�e.�t/RG?3��~�|�o�>�/�Ǵ֧�e͟YU�O5�xs�JH�Y��A�O��uZi�^�>�J?C[�e�/�D>�:L2�d��,��cN0ɩ��,�)������7,'�Z���Pֱ��)Qlm�l/��")`f����q���2N+,q�0�r ����
n@�P�LUI���^���N� V�(���xE���Nb�b2�U ^�i��	�n��w�m�J�ì��yp��.n�<t`�Q2������v��@�������q��7�T"��0��B�N.�i�Z=&\B��M������]Q{_^����L��p�ZW@W�	e;}׷���Ͼ���@"��,n���jO�^`��{�EJ'�������<�cN�d�ʗ�GL.vh�tk�$��A��������?@��fج�Ѩ bc�	C};�� �n�(%�?q#G��(i��F^3 V�AR ��[��0�NkW�@�ny뷘���y^�.�k�����{�\/���9�ɥ��h��@\�׊���[*�[�[HK���ϽN�P*@\��7��>���Cc�\�{���8i�/|�v���g$�E$�'���S�UGL������e�b�eOc�H4$��Dָ���8�j�}�e'o�G�/��_˩Ŵ@�B���r��+��.�a'���OSi�Q8��c �UŘQe���L����4���:�*���zWt#��;	��
��sC�fm��m�6�0�'_Cwc��f����DB�BG�0ޙ��!s�B��� ΐ�B�M=���ŏ��+{��g߀��3�D�@���̐�M�� �~�M��LJ�������p��̻%{�+�����R���&���=#��` j4-�o�k��~e��b/�6��I���k ��L�J��̗E���M[����z�A3*c��5��;*��9�6%x�\q=V���z�Ďd~l�ы�Y4�K�hV�:��.�@<z���j�� ��By�|Ih��nvmH�"�rU@�Zq�*�#2�6���|�yG�8��x��l����=o��x�/������Ŗ�R��A���'���4�@>ޏcW�}鵚I�lJ"��ėw̡���0�S�"��:�Kjڧ���X���l"���m� lW4�W���2�&>K��Gv8x&_��K/�,`o���>a:��6��Ƌ�c>���zӺ�Y���i��k:��0��K�Zޞ=�}�y1���_���7__��wX�3N�HP���������,1T�T#�yu2��Tw&w~=�i�����s|�0d	[�K��Uu:񖁽F
{u����<�{yu�M��p)��i���fI[��G�"]��j��+'oSPOi�s�uGoG��BL�T�m����0sU�:��O#Ć�d�(1_��a�I_<�ЧM?n?P�꫸��Z�,����~]� j$�K!�I����h������d D��3G��ᥗ�H�{E���SQ��G@Y�G�{߯��I|�x�̲�8���s$�K���SB1�VM�i-�@�CE<%�����S��{�iu��fG����\�M��5�@�:�P����1�fC<A�-SH~����x�wסk��I��ep�w%����]���ۢ)3ZL>{|4��"��V��2���������
iX�"�#چp����j�