��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����+��f���-��i3-	`�D�����t�N#mh/M[Cr�l��c��kX��$?5��<~�������y7��GK�Y:xX����Y��*�0���0�D��ǙK�ͣ����?��ۅ��?����{ʿ����r֛��&Uۿ��Y���yv�=��b�b=����)���Q��缭 V[
�/�
��x���1(�����q�% 2�*2Zq�'��/,[�U�J��uX��t�aи$%�G�8����Ì}L�+L2}�����`0�J1��[%�Z���F ��N'ĝ��"X?�[��H���DS~	s9���>Y���o>BU�'��W�v�I�-�Z*@j5�g���anD$���C3IF��#f�Q�8���S%�Y��G�Fm��RrF�����%a�-��2#a��J۔���"�gظ�>�?E"aN�_���O�H�hw�Ƒ$劉��}7L����8+�<|�z�g%��n��.��#}�'���u��f{����8��f��z�sh�j D1�Du$R�+�ڿ?ֳ��v��\�+Gӳ��O�\+5��+5�	�����{��Iӊ���5���Y�*S#N$�e뉫}�rF+F/�s����dB5�R�t�� �;���6Y@e�脆�kC�%zq'{2]sZIs�J�pZx�,	S$�����,�ד����]B�~��±qi��"6��X#�@T^i��
�߻gH[��I%J*�Jq�AK]�R�$�����R�e���X�$�X$`.�'�?E�YY=�+��$M,�g�瘠? ��3aH�>��/���u�_�������Sm�+����w@ږ��PUi��Rp�<�b޽��0�|!@%��=y��":Û�g�+Qg)&�i^8h�7/�c�nc>�@������Lrv���ܱ�D�X�4<�/-ݿ�`� V=^�w"�hh������+��^����̬�up����������G%��|ww��R\Qr+��	4�RB���g+�����T����>L:�Z0���9�3K�h���$�������Ri�ζ?�ę���<.�Fz�E�����(��A �+��_��T/�f�B�㮅�*��O�uY<��Am��+���;%�E#���#�_�}�sJ#=��YC�A8�D�<�~N*�E�8a���7B�_!$�bN�`�O�]д�}�P	�5�YrOm򫵫�$eŽk}E�{Bo7�����9]MR���#�h�3��"CY	Yٛ�g�c;o�1��B�m8�7�Q$z ��+�:{�{+�\��AL&Z���*�4Y�?�U�o������q��x�ڝ��Q�# Ӂ�L���&)a�d�7�͗B�W@p򽏀��i�[+���Q�۝�#`�o�yfǼX�e�+G�˔|��O��vvRx&�<h�aڈ*}�M�Ӈ!����|���0䮦>zd��_��i_`ǚ�qB���5C���'�F�#�	S��'��Dp,���j2<q�����E�N�)3$��v�tW���#�AE#sʂ���0ԯa���{ �[y��oZ+A��T����ޠuƒ��)�^��x���C�L~�c't:�m��gI�q��!W������I� �l9<cU���MY46�P�Q��ە��8�����BVq�����D`�0�;�6Ayߟ(��H�w�M��:4L����871�#k�������=v�Z݄�ol.ePڔ!�����ߦ�6����rjJ�$�3r�:�����[�&ȑI:!A�
%m*������1͘�{f�r1`�s��2�� 2�-�@ uPQ�1�Ǘk�:Gw%t�QEM^ $�X������=�x�JP���ϫ�I7�9�CѬ�浢�/<RZ����R �Y7� ��ܞYS��E�=�[��gT���-���L:�{�&ј����ƺ�_4��>�k���n����H4����`�����Ԩ���G�.��}�.�4���,n=}�`���Xb�:���Q�����!��?ȼ�l�CDo�H�=��LbT���oք夒0*�����/�T����51φ��6��A��Ы�]�r�b�@��/��}x� >�U@��Q�;~z�*��t�[$E��+���y${KʸʥrX�F��jΪ�j�r��	U9}}S��l�w^R��$����x��,7� `�X��<�9\�%w@#��ՠ�Al�ѳ�R�0֘<��d�H��9�.�Tסt���8�0���o�рZ�\��3������8�t~am)uA�1��
��3��]*D�Z@�h�)���	3z�s�!	��5��)��&�?����\[w(���=����e��Y�K�~(��\�Z��vlo�����"~��Y-u��E������!؁����
S�	2{��o%�
�\��OY�rD&Py���	эX/F�t�F�pe��g~P+�(�-x��hEUE��!����#]F��9� �q�0�(�WUe<�.`�T��7����o[��  z&@+͛��N��q��x-��Rȡ=�GE|�+(D�.s�Zr�f�`��ux���Y����y�����ޒ!#�=9?��Z�f(�עHE���U�k�+���͉�]�m3^Zq�9�sg"gV�B���E҅$�"�"��@oE J;A-����}ݒ3�y�4<�Ң�/Den�Ş�@4c�1����{ѝ�͏�\I��w��8�~>��ڙV���n!�d:]�/�����g,z����4oi��~���REIH�t�j��:*�4!H\��;�7�l'U�P� pDG�`��RnB������9��uJ0�HF<�;�}�p���c�o����w�B�,�b �V-����\
��ɡ*�=�̈́ͨw���.L�#`jV0��0�cR�Q<$4;v�SH�14Sk}��:st���t��_�R����SB�5��ӟp�۫~,`���@�.�8+� z��n����m	�ڽ��n�AbPW��-��uo�U.(	�]���jC��EY�eL�.:��ge���������ȱR�~��*ׁ�����!m(|��f4.
s�Ƞ��XJx��I���v�K��87egJ�M=��ַ�&���MI�٠	lC�x[q�E����+3Kw�ъ��w�I`;a�H���N�-�ʑ� ����}j0�o?*�]��&Q�J���kj�1�rJ���a\�D�@��a*B�c�<�	\+E)�d6��(W����{�	{�ϰ�3�D�(�f����1�_mnI�7���%Rm��p�Hv��i�1K��8�K�����f����Zx*�[��d�fM:�LN�)XѬ1d�nU�:+�6���^0��U#s�S(���Z��˲��k|HR4b�ե����ԫ�A&籛sx�*��_u���37f8+?r+�5ˬ]�x�ة���f�6�:�-\�yꍀ9�ʖQ#���f}���L\k�}��K���Zf��/p4ZF�Ĝ�������E��AbE2�U|5f:����c��$�*����\���uO}�7
����K����ǖ�oS���jN�xR��<(�c]�50�a��?��w��yV�8`�P8��$���^(h��ٴ�Npk��N\�!�����W�(���I�B��G��=yI+�h�,�΃���=�NǟU]��KXB}İB�|Q�cǄű5A`�w�&����>�m)�FY��Z:�A�F� �	Ӎ�Kl�֫�(��4[�D�v�Vb�#>m`-�u�/~�+��ݨ����n"=��W
Do��xUp���nL��q�b���6#&n�e�#N ���{��c��t:�����"����1z��_G�F&,�(�Λ�^���XI� K��i�v�E���I����ؕ�����g�8`t��*
��N4�ú~f��"���@�+�(�Z�D8b��0�b�&�	�!]�w�̈�ow�n{r����1_�+w�ɔ]�vm�(���Z+3��~qo.f5��a��/�2��`��G�I��>K��p�:Me��:A�=�'�׵}|���7�n�rAY9���&��`r6���@|���-����陏�3C �H���2O)Ď������9�iU���� ��?L�)�����Z�D��=T
���Y&3�+��C�}!Il���XW�ך��� jlh�G��G�񣞀@ׂ@K������K�_v]r.i9�H_!V��t/�h��uY*M44#�D�87�(���}����M#�bd��d^C��+�����Ì�W�c8����Lwi�A�5����n��=��_#1w{�_eT�I"di����y��"}��i7}H�X�����Ո�l������*����K�j�B֏Xv;!��4����r�o�.�{����-��8�yD�y��ѹ7�q�Od,�R���.��y�ʼh�vRc�/�)&~q��髝�v/���w��܆-�f]�(��-2��&�~��L���P�ܔ7L�ދ����JR�P<�49IE>�҄�ھ�7Vf)������U�Lk�;!Bg綴��
Cl'�Q�Hi�.�~��n��Ғяꉽ�^�0�F��S�J{��ie�գ�I�g<��Th|���E�#�XPIE!P����2\7�TiA�ԥf �DԺt�}h�q#W���O������W6���WV���.��D����B�	��'��~=�g�/��xM+>���F)���j��.��,�5wT�(A�\޹繲#Xi����a��BK�	&������7��Y;i��V����zT)�U����e�_��B�3�H�|%;pX(GS��?U5d]�Ŏ�{Ó����<�ֵ�Q�&��	$ѕ�]W�sS�Jux�X_�R>���r��S� >+��9�j"�rѺ������"b9�}�g�I��ۑ���N��%�y�CT�DIKK?һlg�}�.
�7�=; 
�x��"|�]Y�� �o�����G�	 �/�G������Y�[����1<"�%�+��r��$>D��(zu|Y�\:�b�1^�׺R.�Em�y@T+�q�]��L=�F�D,7v ���mrq�K6�'Dr�� �� T-�"T�M�6|M�g��T��Wz�5j�"A*��1&~۴"�.y�ܛ$GIr8����nv�����4����]�#藽ġ�=��O,�g����#�K��*�$�-��'��ύP��8��+�b:3;�j��� ~w�	-�!ΤA/H{��E�zH%��w�ڥ"_��w�|���-�N�Hvbs