��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������f(�7�u3ڄ�Ɂ�M�Y���-4�v��!�<�@�
�|���w� ��Ƴɉ��/,O/l�\�Tgwk�6'CUK�TOq7�[��~Ȣf�~0���Ì�j$Ӹ�P=���K�����O4I��Q��O-�y��q��*��&5(�h���j3+�-�X�0C�Q%���Z]�cW�7Ո,��7��GoQ ����m7=���^�mit�Y M�S���wO�L���ĉ�}����a,���饓�/�{l˛[YA��2�`�x�\X���`�I����G�������%R��F�i��cL��Q�I_������1YDÅ��������6�x��<A��z��S����A�#�+��(�Q��{}�f�Z�ِ\��8.��\Z+��nxU�c��k�ҩR��7&�<=�{zD���G���u-�A�S����S�D_/;d�����������Ѓ������m�A�{�_�?�x��;h�0U���s?Sx=������8�Fj�4W�D�qGVB*���_-_Ȱ#��v�`��ҵvL��u;�e��/�v����<QC���MoH�$�U}��su�oc D1	v��ڽ,�4���,�^�ь��Ln.����P2O���3�ºs"*�*?y��QJ�<nyN���l[|�	�3qD(����vZ������[���@�>�m�"�q�a�+��$�{\��8Z6/-��t�T��`%v��D7���Z@����!80a����"�DX�|թ�N�>Q&^xX{\��nU�L���u<�Ԍ5��Qగ�'���ϓP]+^��(�[��A1��n�]����g����оϲ�p*�A����� Xy��&j�Nvw�r�S��E��"����	� �\�ڄ�-T��0
} b���g�8���Š=U�e�A������Ŀ��˖�D@֞@�u������5�$k�l�b�jE��*�|�7��0�����I*�e�#��AB���7:���B9��l�W�bJ_a%� 1�Y�ӓ��ڂtѥ�3~��ԨC�� ��\dɎ���p�m�5�cЛ�b#Zj����5HaI�'�̅~������ȍ	�^���*�XT�g&+oܢ��V>�ű�M�C���C�w�@��5�Z,+�J��W����I��n�t.�2a�$÷
�^��hD�ogZ���Ӌ=i��ŉr�k�6��J�4X��9r_�v�{d��W�`�u۰ �
�d�Ҍ�Q�UE7GP�</��h{�m�N��>H �T�:�b}����lc:h��Х��=Q�&�S�t�W�*ݬ�.�#+05aP'I�C'^�N����;���-��Y��QE���겓���zI�e��Q}�5��u�%��5�&����;9�}$+��L�ž�z��Е���#�%7
�����=���8
8QR��q,��8D����	��s\�b�*�lؑC���b�X/�����;�s����N;;��2.���׈3$�.��8��/9�y��R�n��,����4.6Ո'�o��Q�w�I�^��@����Vrg��u'��ժC�@J裆f*]�3��h��Х�w�z���l��ی/��A��ghu��K�܉9�Qg�Z"m�P�?����0�8��[gܛu���J�oӀ;{?&ĝ�7S#Vl�7�hQ�ռ�i��SM��=�f���k�ߙe-H��X@�!Tq���U����qF�O�r8��J�з���F� ��Վ�m��1ׅ�=���"�1�jt��YF.��W��Z��s݁�m��)-���V��<)O+=��6�{���	�������"Q���͏"DW~EН��9����(2z�I��u%㠺d�v
�_�gkm��/���y��+)g�g�8�4��3�D`2��▎���M���N���p�o�rLY{ eRp�H)��q�G]��?�?�����d��!�/&�
��%����7*v�:1�gL��Q���
t���U��s�ӿ����q�_�=�^r B�_b�4�,P�aK$������j�[���ope��
@UĽ�~�u�p>'geܧ zR`ٳS�N�e��x"����K��?II�}/ۀ�~D��&���~m��?�|�lN&��Á�e	*C�l� #����=�Q�O�ď�+���嗘(�&�S����<�(���"���T�g2	1��`�̃�\^����Cޫ�ȶA�-�\;/����>)� ��":��?���D�u����٨{�Q���o�Ŭ9:Y|���tHe�U9X����7z:��'�������g�qW��}+y^4Uy7�ju�	�|N1���}��**ޫ�դ����V�.0�Tvm��pշ�Rߚ9����[�Ŭ�ńvyG"�F��߃�_�̞;�r+�����_�\k���5:�($��r�m�nr=� �a�q�+��W�N���!*S�ڻS2�"J\���T���"�[�J�$*��#��A���TbKT�Yk[<Ύ���u��ź���� �vSq�������^6n`d"���nL̰��D��](+iʡ��,k�@)$���>e#�ь�|��d���(;�
p.��~�B%"W/��S��	��{��0tȻ�'����(��Z�5/khU�#�K�t#����Y�K
l�[º��o��?�����H��K���BK�q�t�eȺ�0�)���k��Ϋ?S�9��پ��U�>�|���J	�[��"�ڃlG��Cx���L�p�?�+�=ydZ��ڄ]�ۡ�UmK�>;�Yٚ���{����b*"}�YF�?�ӓ���EO�4&M�:-#���"3�
�I%^#�.�fr��Ñj�iSm�B�&�!ф��%�u�0�C��zw�aDrt���X���Y���j���D ����ЮP�;��vD~ښ���^J���d���fz_�7�c1DSU���fk(�U�#��L
��L���d Б�Ä�>n���S�T<r[�*�8rĦ��r��I5�nJ�ǋk�a����
����8OQ*�q��zF/����R���Wa���[_^�
���A��Y�aQ�����%�����#Īk@�N�s��B�	�|X�5W7�"��Z���ͺ�]!a*֘T.��A֧w�@����BS�6E��؝���K_�Je�y X�F�@�r<����U֮�Vաŏu���Րf�?(
[�����`���>��~&�0�R>	�z�\&�؀6�� V�ł��A��TG0�!­��� �z�"�H4��Е�	Wv�n^G�0��l	��r��x>!w�qLY��gKs�W���&����`�`����g�gΧ��:�	�)d�s�G�����M��������1���/��B��ۓ��DH`b��n�}]�zY�`�hiJ���f.��\U��pȠ�7}h
*�:)�cd���@W����|������o���P� =d�&�znuS�7�/��c1���TxA�0^\�JG�/Yj��6�ZT%�AM��}��$$��M1�i��۷�x^�J3�	!R�vz�/K�H�Imz�b\����FM��Ds�E���Ov��0�F�Z%����cl���RNz�K7�3O���-r���W�@z���7�4^�5� ;�մ*�tK�WTs�|bm� A���&����9?��wD-����W��m�ei�=NY �M,���~e~�G�*i5.W$���^}h��R4��$�~+���{��sͷ;�%�\TU&���3����3��[�TB��1�+��v�I�l�^��=�u���ˇ0��x�J�;�}!`>�_2�r�d��6�/�#	s�,v�Z���u>��|�8[�+�
���S�^�¸�҃�}7]�,b"��&U��7��%�q�x�(��C�� ��	{���L��)V�b?��t�Lˉ�o�n�"}c��>I���nQ�����s�����8k�J���!<C�����5�� ��b���MҚJÔ�ƶ�=q}1�@�1��guG��iv������ъ�H+�8��s
�o�gQ�RE����m�X�J���}�q�u����Y�/Y��]���+��^�#�D�\��#L�DaO���B�����é����`at�]¢L�*�d�ؔF6xv](����̣:
#%"ݻiA�m�5q8>� ��;|���[�:�T���Bٲ�.<��0�0z��I�o���l^
��,u�>mĚ�>��Or���f.^�ú�������I<_"wh��%�0�H�ŪӥQ�*2P�����<.�����k�v^���k��5��ѷ1�*�ڎ��g��"Qm��/��{��V�l��߹1�%M�A&0G��~K^5��������A�j������ɩ�zb�6����d<p�ZS�ݧ��g��M�G��>��m%���a�I�m���^����Z�
��a�/���D��Od�8�7��C�4���	�}�����:aU��T|5-�WUT-�.a���1����dQ1�a1#��ʙu����s[_y���߈�V�c_c>����7��U��-�b���;F�\�7�,�g�JR���_R��oclʥ�'n�:�b�c�6��Σg��9� �2��w�s�/K�?v�h�i}���T���g��z�&Pקn��� �p����gfQ
��v���`��*��,ə�v�I��<��