��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~%���4��Ҍ�r!�4K�����|ű��p䤒.��:B��d�y�Pw��v�7�=#�U�c#��TJ����wj��h!�m�Vt��h*����H��cyDߐ�v'Yg3-��:7��h�����$�����?hN�ae¯�UR��J���sB�`z�R�"��бAd�o��=9��D<��g~�f=10�����Ӳ�/Dx�w#g��U��`�V2>&0q�t�ح�pD��BOh�̉V���3�g��#��z4�o$欿(�$�0�;�B�w������ڍC���h]�5E�=Sw]jw���?��`��2O�ԧ��+�*ذ��Q�x*�+�|R|�iLGd��Kܯ1[��@��o.�^��r>^Ew����2/�k�Ǿ�wܯ��Ùk���q(�n}�~�P��j��B��S��b��{�7�lQ����_�K3�{`�,�K�\&&T�ҁ$,}��Չ����6/�ͯ!p��S�r���RRo��x���Q�-A{�#�/;M�׺�hV�������),���Y<ֺ�(Uc/����BM�^��o��vZ��[��Wq��}�{�+�?�ۼD\'������\IhܐeU��?�4�Ni�C۷�ܔQa*"	K�;�^+`!4AF�0�\e*���M��QƱ��>=��.j�	��3�]�O���� �9Q��F)��8�i�P� �tS� U[���
3�v��a: 5TM������e�{��Σ�W� mMv�$h�=#EJj�=4J���J��c���7�<��=����܇���3�VJX��8	�������#�Y�,ߣ��T緍�R�a/��I�R���XYE��⍉xN����;��S�2���X�Vڍ��Q����⻊����f�$޺$|�����d�L�-�$x<�9��H�hg���@��M "��8l������~{���}����5�hO��@h_�|q�����|3�"�\`��<�K�K�TZ�yP��d�!��p1�y1�E�ϴ�w��O���0T����G�r��� ��c�6˓n�OޚP��#ħz��i�l��^�MJ�ղOD>\+�x�����L��Qy׶�y�
6Xg�'"�E���C�C�*��^!��-!`�"\��-<���E��SB��w;��K5S��! :��S��������N����׊>墳�;�<E@႕�t^���f�gZŇZ��f$�)6NO���*�.rU�Ca�e�kC�=V��:�^|@?jbO�A�u�P9����(7��y:������z��>{�ZQ��&���^��9	�Y�Q�.�<y����Y����=!��8��/]˕��4͂s���0D�V	����()���;�a@�������EÊSt����Q���~'�0��͂.��m��9W�f�����L�v��g�u��xj~����'�*X�yӭev�\"����#uqm��83|X�?g�M��\>N�q����-�"ዣ4G�0�Ϋ��
U�X�Ev�e�4ELƊ�Cxk>p�mI�s�3��)lz�S双��_�K��������B�%x8����0N���!�k:c���q�.x�zjB�h�����<���z�U�w�.(�|����[8���'HF�ĖI���|n<�*�����@
���Ǹ\s���Xc6f��:�S5~\�� ��4�@�&�;\-��4�rO��/w��ęt�C��
mL�eoPj��fu�J3�e���кKgzR�}X巴���9<9
�F�u1�/ $ @ۦ��F��Wҍ�D!��.ZI�U�C�)��+�C���}��I����VM����k�DSg6�xAꨥ���7f(��";zO���w��p�g�)z�Ifɐ�8�̥�yr�!az;,S�^��w �+c�;��hlZ�Y��q�ے��?w7.Χ炸&i�[ˁC�N�>ȉ�k�%�%� �I������clBߩ���Ҏ�sCF�i-��.9������&h��4��fw}u���?�Z�"n�]�eQ���*T3g��~N�̾E_	����A����K9K�|�1�"�Sĝ̰w�T��;�I�?��'�X�3��l�'6j�B٘n7�D�������QWFJ�?k��v�v._�����>�9�p
�
7x.�17f���QF	�$DW+�t>��Ze�G�����k�!찑eZ7;��B�J�C�)��^�|�SiB[#�3���:�璠�=�k�J��ڦ)�i,��椵{����6�vpF���C�.�>��݊j��h�Z�"w*;�v(=o�K̝WҎ��	0M��oG>K���y5�+{ݓ��@j�8-dn��
7� =�q����}Cz�Zs|���և���/�7��~�/iaOd7�����AH�L����\�+��RPxJt��)M�Tv����dH��t��}����,�H��Noٯo���~B=�������ߜ)��A��a\�Ŋ�t�F:�s9���ַ�F��ſγ�yʾb��8���"t~O� �b�*'��[H�d� VN���6�+�������V-����4��b�xxl7�J�m�N��P����85@��T�>��h���L��T�)v�Wup{���߫�KU��d�c��@W�l���B���&F�m�\�0rO�����=�i��H0�~�Re�I��)6?��/6�]7[�U�8�f�=��z Z�t��T�v1Q�u��x�Bm�B���2X#ݩ9m������^}u�h�~j�3{��@�����F���I�,�w�c���oF>Mc�ٽ����S&r��@�I:�����ds����\��D �Lԭ{0���Q�~�~��H<��o�K~o��6�ڡ��;��2ά��{��G� �-B���c�l ��K�R�C��$s������C��?�~,�Yل1Ʋ�qIL��rInVr�������NH��cM���0D�Wۻ^�B%��+
��{.{ڌ:��;�+��y�@��k){@����"�̮,�/����`8͘i�i��e_9�D]��y�k;��/�Y&���o��"�D�|p3�Kg�uZ�~Uۍ=��+j&�Փ��A-��G*�E�m����c�@�_4@z\#:�_E� f�%b��/,&)=G����A4O"$E��Hx�d���C��j@R��_�(y��=͞��m�?q/��g�`�I����2M�L�G������
\w|o���#�g Vz.Z�
�K�������j6�Ďߋ*Z����	w���42w��*�Rn����g~��A����&
�B��7��\nNУ���O3i+"�����|�8�Ȃ��|M��r�k6K���.��0��vu8#+����t�ᆅ�¤���\�w�6
wϰ��ނ^���QDU�*?BL�J^���K9�-����.�V�7�xA�ԑ`/]G���uN5�C!Ta��BY�u��B�B�=�-~�!DބcւFD�,��_!�C��1���9��F���@�F31q�_
�+' ��^���x$h�WD��g���9;�b^�A���'�<]���n�h���M�� $sEBd��Q�آ�(���E���u�z3����z�p���~!oǃ� nB���� n�_(�����;���J�C����)7�F��ˁ��Dz��uȺ�<�uo������r��]��N�.Q��A�"+_�����z_k��OL�T��CqhLKO��2��b�p�V�#Ķ���c~�/�3������,���Ǣ����y��BZ�U^2h��Ϸ�ÿjl*�����<.^�v���@Y�"�S�*���SSHT��*������,r����{�{)����{�R5��?q�gS��l3:<�,���3��yMq9�Y[m:�?_�^���J�7ʎ�m��*��������k��d�c�d�����C�O�	Ђ5X�z� vA�.�O��/}��Y��IK��=��6c���G�� #-��t�{��͡�}�,�����T��Y	�3�&�^�*5�
�PSo@3L��a3u��`# VE!
1��_3�*%=�pp�r���l�	|�:��'�H��k������Y�b�Z��P`^}C2\2�-���A=a����Ɇ����5�b&K?�+b�yi�35�[���$��s���HdߦCjmg���O�У�&c�����m���8N0y�PN�����E�F!�l���<U�l0/]-��<n�(������	8>��Y��P'�0Rl#s�%>��d �c�[E>t����>��2{d ��}�>���f�����E�x���G���ļ~��ތ1����i��brX�H
�M<���������2S�P�؃T���W����x'�����.-,}�7_f�-q��i3���En�F�fG��%M�
�]Y�[�|Z��D�E��`.���p��._R[�`#�9�撚�����	� �i:F���%�
̀
y������q!%��D�(W��wSp.-�`sS�e� ?�q+7��{Fd_.|t"���l��8�%�PIߧ�U���opH-��x����uh��j������Zr��25�Z	#Y
�����~o�'^��aT6��}S������X��/Ԉ�J�1�F׈&!�_�
3W�D�"��\#%�}Uέ,ɨE�Ow���{�h9�k������aS��t̨�jF��~��W#4\��g��J
5A���1?<
��g"�����k��!���c�,��P���u���,}�M6���ev㾵���+�#�3�����?_�ߏ22Q(@(���R̡ɏ>>��?/�'?V�zx'rSl*�u�4�V��޻rD��0
_[�@uw"��f�O�՟�z�	�g�V|*
x@�t�c����P�$���9�R�q�����~E���Y�	r���.z�h�����d��cd������<�7���1]��S ��,x熕���-Bx��+;�`��9q|�"���ة���D�y�dN�7�<Rop;~خ�r��,�+�!yU ����|�o7�k�Ǩ��[��C�ާ�J$�C����U�^�^���AW�'3g6�Ԗx["�=8Z{R�Q__숳6�Z�6Ӭ# �����<Ըמ�^�C+����b�k���ysc��Kݜ��p����>Ϙ-� LG���{���I3�4������C���+���#��,POek� l��a�d�a ������\kQ���vt�����VgSE�0�֌,5#�;�;�̗^B~i�o�oAe�e�����*�d�r��30/Nz�p6�v�L|P˺'u�G���GF0�����-Sm�	������
ޭu�R���6n֛�w�#i8c�:��dk��X-6wc<�{vEް�[#�9�~����?��W�:0�ٔɁݫ�](&Ar
y ���1����*_��H�5Dj�)��[����͖�ǩ�q��%�f,�R�,�C�	 ]��$�bX�h[�`&���&n�˨�'v�
A��B������b�[X������,���X�og<~;���A$�r/՟�R��� ��3��c���d��8󺛑L�� ���=�ӎ�w�����#�P­�RRڿ%(��ľ ����};��v3������S)SM���;(�@l�}�r�Q��T,	k�%y?-�#a#X	���F�
���� �߂�Kğ�ֆA����2��f�|��Ek`�
y�Fj�\�i�� ⦶v�/}� _�Ke�@�7�c�ވŐf�,g!堕"��m>����1����zR\m�]�r��Q�>�Xl���eK��e|�b��%�u0'C�WD�_�͖���� �J�;	{���7�h-v�d��O�"FD?�t* oVe���Gm�Iq�Rfz���A����ɂ��Q{jO8��r�F��G!��F�ְ���H�q+�pǪq��p��~!�';��#�T=t#�sr-����+���6����U"{J �a&�h\g�����|���/�_ēX
;��XfK�zϹe{i��mx�XCJ���k�(�-�m��LymWO�>	mǱGO���uDxS5��a������)�-�%Up��C�G�ì�c)�M���(�>k�D��H��l���]���\ҧ[:��*<���h���[4d��z{���V p�����	H���45�t펇>���M�C�S�Yq��0�l�"v�������L���6�NH��C���6i��A�J�A�����u4je�&��Dv� �,��J�+���P�c��Lǣ�
W�]����(�~�K��([T�Y_�����M�F�l�$4a���r���f�P�u�C���o���1u�YOg%>��$<_�q0y�:����}OB���S�A���c����E�s|4��ʽ7R呔����a D>��m���	���,9M����pl�ԇr�f���X�WD5b���}��n�6��8�M�J������S���hx�4��^�+�R=2��v}�j0<^����	�� �%���{oߑY+��kޒ���K[ޣΪ�4�H�4 .�t<��85�s�9}ǻ {�l7W��x�ϵ����~^��c�)�O���74�GLG�����]iJ�߇�yA���.6;+]>|o׿��p��� ����.�>��_��nȤ���]24��Lȉ���qٲ����������}��:����G��~ě�x>�w"X14�{fL�x�I]Oʞ��#D!Y7�\O;^���P�o����U�c)d\�G���7�w��L:�s��.w�{2(7�(�v�Ӑ�i,��sS���2)6~�rK�BOm �\R&%�� 9{��z�>l�M�XJ�� Ge<�{��g�0�O���M�#4��X[SQ�]q"��&�{ߧ`S��Q6}QC�)T��MP�;��*>�J����һ$ﱄM#�k��D,�_]��|,^��4I ��ą�)�`Ƅ�����0a5Lܫ<ʡ��+p�����<��j�b�:��\{�5���m&r��
\i���ra���r���Q�#�Kd#mg)��0[��ţZH�W��:k�p�����R�OT@E0����64��eZf�́?Pr�C��r����!�<���i���;j�U�G������a�}���1ݲ|$��3U�/$�"g���q �7�ӉA���T�Y�r'Y%Jm��w"�{_��#5�+K+��1?QQ���t�>߽Hla"�n	J����<�����K�7�H�XR �Ҝ�l)S䔠���Z�^���ʐ -�}��v�Tb6����4� *�t�|U�����إ���
��]����<O8>��p���T:Ll�{��`���)p�pO2T�LN�[L��y����Y~�8ޟR�k������2쾬<w2�������ڦ�KG��t�g%^^:���L����V�!q�|��U��/F�^R�5?q���I�ZݺA:�_ ��B���hn�B�J#��q���<�$�o��a�a�9;ݢ�N�6�jh�_p�[g1�vf,V��|��c��$�A��b�CK��N`
e��|���
�' ����|�qX�nF��
���K"�W�l��P7��T��vO����_��\��zS�Ġ�$�>3l�` �c3�Ka�?��6L��Eo ����;2��W&�YR^31l틓���0`MW���Y�de����s�r���ӆ�[�+dͧ�KY_�M?������y��m�@�t�y�*	�P�n㣀� )�G`�R������V� _�Q���n����U83D�����WY��M��t�Ŏ���/ƃ��1��4�nQt5W��(��f�>c{�������%g7�9�TԆI�8���7���c��\�k�{���p6���~,�V�eՙ�)lh/c����6?=0.��G�:8��x����G'�E� ������X��T�r5�|���i"B#.��F��P��OŨ���:{둯'�e���V�e:����\=�?M�(mQ#��� ���>��tY��d�MI��s����;�׺d���i�8�̻��zL��eۣo�d�jJ��s�Wo�e������YM��ƭl�EZ֚�Ω�����/:Є�J�g�����ǿ�66�7!�1��Ǹ�_�1����jټ�[��������;��t~L4�~��mrz��R&��y����%1��d�\h�9:�z�[aB3�x�Ǚh�����XFZ1��H����yX!"�����w�߱�L��NfXJ
藺�H"��xi�Po�y�R�I�Nٳ-������ /e�^^��$�t�5��_�&*5� b{��w_��#�9R��lJu�2����PJ��>x(�y��9�� �+��LeFC5jל�Qb�ǎ��G�3�~�!OFM3�͘�p��p�ȼףV�bB�2����PU5�O-�M@�Eױγ�'n����Qt���~S��R~7��c���	��\֫��>ϙb7�H"��Eȏ�'�((~\9}N# d_
�fj�0��q�H<Vb�wL�;��Y�������0�IbG�]J�WJ�4����Ŏ{��.�V��x����(�.@�lE4�h�Y�������B�	{�Ӊg�Wc�@����qP����s2��T@�2�$Y�%G��VW�T}$v��-c����I�ڙ�i@����sk�ą�c���g���c��á%<�b�y���K���+��_�rԼ\�ny�J���Ts��ni�
�:'h%)�~�5�w�u�\^H�#6�86��`78�)�4K6��u��&u�g�P}�~�w;�pڳe[lh�N,7�����L�Ő�i0(M�4i��U,Z���y�}V#kP�w8u�ϭ�(>b�� ��'�e�Dw��8���6�It�LKZ�(�n�}��@ ]|_��,�����az�#.3k���P|$ P�΃�r	b!`Q���H��!bg�3�Up�t79���:�2\�E��t���{�G�	�q��ڌTH�0�C�B��H�F}���ɠ�=�x�֞zt�ܤ�Q�p،W��,j�����/g���uڷ`.T���g�Y�"v,DJk����:=�$&��މ�p
�J6���{��>�r�v��R�z��t|��ö�h`��,L��r���-�vܸGó4��C	����uٞ��ED�_���qZv������v<�h��v��U�5Ξ��7ۇ>hȇ!�fa"�VB�`�9��"3ڢ0�`�2~S�B7	���F �A�|�o��S=�1�B��g_�A���	'F@���x�k�Ƒ
�A1\�{Io<�F}t8��F`��m��cФ�sqt�BA-��I�& ]�4��#����{^<�ˣzo!؋5��O+s�o����6��N�D�ޱ�>;C	�&iǅ�DR�npN3���B��k���-nҋQQQ����ĵ_eB/*���8���]��ԂD�Q�B���*kE����LԆi��	y���g�xs�T�Rr�)��F�*_Όi��h�MP˹n� x> �hn� �+����[��3hS61%g�(#u��vi���~�Q����G�r���P� �Uh�ɏ�)���+�tK�o�J`P��R߀U1[L�e�~��O�b�=��H�Җ����l���.d�z	#?@��y�c�AuJT�l�2��
W%��� �ѱ�����"t
�B ��,䁦�p8&�����%�=å>���)�����Bal���H���e��� �K]pQ�?2�k��ݭ�"��H�F��@���yn�m�>k��������N�l<�o��:�оAoFO�����Y���|b�e�����0މp��v�:�~�,����n5��|��b�!���7P�I���U��FſF2����w�:��
ڱw�A������}h�8]Y��?�}�d7����i�\UQh��2��yf�?1NQ:'����:�<�6bX�g���f��H��Y��vmhM���Zn��C=k�ճ��w�t�4��L���r��0N-~z�!��w�2�w�0`���l�k�\�h�<)��(��t*x��F�7�����L�R���@n�BLjs�zK��w�K�͎�
k���q�o�r�θ�A"蕿�Т��<�&~�ۓl�)%?��!n���o��"#5��:���\��vA�#�l`���/Q���L����� �U���w��UG��?�Z�[[�����澽��F�0�������Pp�pIC-�ෘt8�[kN���g|]CrC�qK�*rEO��)�������tD��L��0���#^���4]��pl����&W2�G�q�a�@8���.��A��SJ�	'S\����!�g�{Ɗ��kt_�u���i�{w�t�������e�2�\6a���e��1�z��A��XکKD��|�<x>c��6-U�>5�Z��,A�U$M\�-K�4z�T��jY`˶�t��6\���Cǈֲ��J!�`�v�7�<�������kP+��o{Y�O+�I/���y^�D� |�O�}��	���ĕICeI��>0�R���ԗ�ϩy�Um1�m:�
:�����������0��1a��������`)s�� ��ԃk;^�X�ߴ�֨�K���L�{�K��M��^���1��f���~��^�brZłH�ք�N��I#vi��.�e$qѾ3	� *kq?���� ��'Pf��<° �/P�N*�.���k��ME� �U�$@��O��5���7ʷy!{��2�V���.X\\�ϛ��7�m�t�
os?(z#�8ѮEN ���i�ۈ��i?_z��2���b�=���u�Yi �O�I���M��s,8�B��Z�Z�� #M�ڷ:�`m�z�X�	na#˿�
ư�¼1�nXJ�6�\���'��}�l-�EO7�DuM�q?oG6��I���l;7���� |v��$$M:��y��P �S�thAB�n$/K�ތ@������۞.�>0�����L+�|�S�yR���.w��\C�����k����t
��ڀ��8U�s|����l�E7��A#�߬����ΆdS���/E��}�����:��tuM ��ɡ���U�u5�U6i1����HC��`d4AA�V�A�n|�ʍ>	Av�/xL�e?*�8��4�'[�q$]FKlV��,��l�M����0�VzSO���ġ��
R����?汤u�JTvBp�X�ʋS�1�`�B}#�*��]ަp/ �qxY�>	�� ����.䄾���CD8�+!qɸ���\hK�4��-iiq�*q�*�wN�C�Ϩ�s����b��#w�z�Õ}��-�g�_0�g��/C�L	��1�tt��%����Od4��mi;���<v�4�/F��h�fjճ�+y��95���Y�|��ѵ�O��C*����bq"�31r�g,<6���8-$F{���)��l�1�H��jb�ց�� \�ՊeF�_�5����%.����;�' �Ͱ얬��l��f���+P�(kk�l #lf[�3��=�O�r���Qngs42XJ�c,��2�� 7er������_g��CN�s<��AT�������Yg�
����K���<�sSvh,���0!�	���#���Hw�L.i�*��g�^b�v�e
@햸��-�߽yvGv����� ���n���(�;@H�}Bݎa� �&	�ײ�=��RpwP���5�b���J/�e�J��Q�*t,k�E����u��ܱ�#�������o�p,3�C�1+���n���d]X�j���Z�|�Q�D-�a&��t���TE�NF��wҝ]��Z ������{"ýl�]+?L8 I��n+U�Vd�~���+����,<�����^i�;Zk:�y\<�'#���4Y,G�޸%Y��V?��VHt��j 1�X?��?��2�L�������2TT圤��m_�n!��ߜ�r�@������e�lܟ4� u�I��?O���y�V��U�2�*>9"`	�ZP#
��+zrw�Jt�/�3�K��l�R�C�c7�ps�9�[��Y$���J@�k0�gS_�P<��f������|�����iW�I��%�c4�vQ�u�vH�/H�K!=e4�`�?��(�Nos5ӈ�I���eh�����Sy�B�䪟T�u�!��^�g�7$�2�7I+��a�Z,B��s��(�m?b��o�zb�2��XNXvzV�b�?��[#4�̆�Ɔ�X��4��q��'Jf�.�c��׵Oz�<~X;��g�f9(A�/烁�u@�y�v-E�����P>^�ҙ���@Q�sg�)�}����J���	Dch���|񠮞��[?"�"Z���W�$e�W�Ng�$���h3{7���y���w��;\"��]8$KA���A����V%e#&�X�Q���
=at����'�5z���e�ĄX����ޥpj��P{��'@%N**�\��[p}
y�]����/�Bw�ඨ�[Z$�\�8� �]g�☵Z	���P�$�PI3��^�bL��N�D� ��z����m���yC�xn
2k��V>������cs�M;8|>)n�؂�0��y�.��/"��9=+�(���	�DB��H�C#�'�&_�IA��	��Z�O�5ڏ%���v>��9���9�*_��l�1��.�eM���w��v��;��*�,�$�����s	�?H����d��)��� �?D��e�
=����
ap�I�#SM������m�Xo8�"���<���]ʴ
j��9\~��`�sn���F�J��S����׫L|z�̠�e(k�����/!�� X���)���-猥Q�k�'Kc�i�Hv_Tz�W����?'���B�4;�V(gЁ�2w���}<^t1�$[v���  gV{&x	�a��6��88�Uk�_g����������%�f��U#��[�^�!AX���k��}��&�#L���O[��	�0=���z�1Wgr��=��)�;�O��FM���m�	ڣE�Y@ѿK��-f��K�m��j���&�_|e�)q6='�9|F�;
k����RoM�UX��.�D[?��4���bC��]��mųՔx�e���%��:�۷(�[9���������<��P���ֵ�_3��@ވU_��Vf�09D����&_�)|����٧S�Lh�I��xn�K���.����(�b"��M��2l��R���("���;����awL�߼�6p-X�ˮ&�=8� ��O��5�O�����z>!|�r��v^��s�7�-k#WS����]��Ʃ�I>�n�C Л�}���G�ߜD�V�I�5Ҽ���|NN��L.=P���̢z�$*z>(O] ,�loTӈ�A��tϚ�X����f�������Ɂj�b�5�?Yҋ�D^�:C�-'�	�XD/��M��������)@9�poʃ-ώ����yxwy�)U�&�[�ޕ>�d�ek��jeor��[�m^��pm��<~��D`�X�Ë�_G�Ǿ��5O��gh��c��1 �ϥ�&�Gu�=X�6^׻.�r��5t�~�e�x�E>� S���-�M��Yx=F�/�͖������Ҫ� ��s(�C����7�ܨ^^���V�`GI	��]&U{�D�-��o^�\}H���O �w� �A�J����K1��8�dQR4��J��N9(r��{�^-��EK[��"���y^kzJ����W�q��P�QHnֵ�K{�N��TTf��M���wkr
+�&0u+?ͱa[Yd�`S����1n�ѥ�-�}`i���y�N�3�X�݅s9>����j���RM;?�:��Ή�x�!5sQ�<OA�BGoDL������)���� �V����c��Q$W����@�>�[���۪}��T��>�E�����Y���%��tt�$�3x<��E�������@蘩�3�M_k�J�5��[h�~0!����������*�yG�S�=~D$_�������&wL;��w+;�-n�4�PԌ����]'��R�e�a|���[�:�{��t����� �+��UH(��O�X�̘��ꒆ���;)��o5�bwz�l�4���L�}b4]����A���3I�W{�I��ҥ[�J�&��x���H��e�I?X�]��G1�FHb��Z�: �J�0��m�i���R��a��3�Xo�fS]��$|8)�(0[}Oދ��`�T&�_Z� ���p2���6;l*��
��nf@䕦D+<C[�c���\�z�N5�֬��&L;�8�=�N���'0��c�P�����Wa��ʊ�d��|�B���gB)B0t���%R���g2N�X�!��6Jv�b�{�L�(�Hi��.m�W&�
�p�(&���ʤ�Q�S=�����:�b��Kc�ߓ�H��9B ����ъ�'����O��gps���<Wa�Q���IA��ϪG��ɨ�睲M�3����p1_���{������Nߘ���s�;�ea!)Ks��+d>zƜ��&�����WT�_揖�6v�q2o;�n������r-޻����S��jz��@ �w�J��7��vN��90��b q%d���ӄ:�a��v�?-f>,.����(�f���;�P�.ы��Ӭ���LKdE�������#'3g\P��y �	��*��cc�9#G(��X���%w�L��|,�b�F�3�����	_qm���Aw.�
h��Z�y-�e�M��;+}d��X���e%T������m�U�̺Ѻ?k
@���Z� �E����� ��NP>�[�i�0�o�;-�Q��l��rRT��?#����<D�@樓ґ���H{�Ҹ�}��Ӏ��N*�R�3<E��*�'�&a$��Ƀ�ʄ
�P7�����U4�Y������TT+��R�"���`�V�E���N�=_�wb	:��l�P��\�����?�7��j�� Զr��]w<��ߗX��f+i0���"!#��/�Vl-q��f��M����~I'�G�J��8���c�T��I"�w������^Oݚ�=O����>+
yJ'���`���}�'�4E�J���c+���TRLE��!?p�w��uw|�K� ����0'�Pn�=��y�3)�(���.��*�+��V䄔��t�����e��R}�gF���a��C�$��H�E�kW�M����b'}Bd4�8|*h�$M�'֬�wg�����y�O0��V���s�W@z<��TN]k���2�g���xpr���Q#]�E�q��q�<�~�������2&� xcS����M�'�i��Ѕ.�	D0�}/��۝o9 O�c���̰L[m�B�W�p� �RdQ�\0o��Qegw*�ʄ�2T+j\+����d=��c�urK_���C-;s7b�kjD�y�(_XI��f�@�[Ю	�r)�m{s��g�8��`[����C:���!`7v��:I�]��xKvGI��7�NOBq���@�`0c��Q���V&PͲj�3�x�1����+�zt�Q��KP�#ʒJ7��=\��D�#�6�!5b��`	�Ĉ����8P��^wuh3��7��b!fwU E��\��6tefl�{�N;iHc�i��excc$O@BC��"�Q�?��IE���F��_���F8R�{͒���bt2)��|�~鑺:��=��lcV���t�6�V�!)��� ��
�r�Լ���tؒ�15Y�?�|.���6���������	\Oaǅ͵;��^ar�x:xezR�QsC!�%���)���z��
/hޱ5���ƈFu�s��1�A��~uW<�i���{�9٥�x0+gAgb��~�R	�����9 ��3T���T���_����y2A!���I0[�n@�1�1��`zr��h����u�k�
x����#��«�Q�-�I��rYw���+�-�g�����]�:���E����3[8c]���a?p����]=�]�ZN:	�"��܄�)*���g�״d���h�o|tш���.���;����9�WP�,ɢ�@.��U�����Ά�ؖ.�/r��ϳ8��,V[�K�҉�Jƃ��1�m�d��)���!ɪ�\���ʌ&�^i{��WL${�>��X�{����z�r��	��AcA�<�:zY�/�Nh_-���y_m���rlj!��B��Z�s�5L�^�Ry�)lY[�;z�S���h|8����j]b��̖P+�yW�g�� >��Z�CE��7���]d�.o����gp����ի�V����@^�]���R�ދ��e��1:�����y$y���[���*�x/:i�y�1��,f']�ː[�9�X���\�{CE���.Ѳ+������W�b�n`�7G���7:P��ػ/F߷J��5G��!�h�/c��Tx.�-���&֜���������W%�j��������6�t�_L�����@�1�`�����׸�Q�C��$1����?��ڎ�:0BŘ��>�9Y�qT�0m���zR,���z �� m�H`�u����g�������I�L�gau99د+���;tst��� �!F���ko�ڍSVa�!���N�{GN�|Ҵtb%rn��7��U3B��
Zo'+&��Νb��rWr'�'�	b0�+go��4�kZ�G�)P�CY�O��8�*��  v7$����� Ʉ0A!�yJھ��.����?�-��b��Y3�K�:�����oDx�]`_�|a^�->�!�����yP�+x�qc�����uf��A���l���H����Μ�/0����$�J��%T�7&���N%$~=�qTl"�4�έ��/ե�$0����.*K��t�m���A^�ovPO�{[l&�y8骙�[����~!�N�=c�'���"��� d4�{���+ly��94B��FS"��3����)�~����C|,�#-�;xC�m�Y��	^?
\���:e�O���t<-����j!���\�����ֳ�g�ՠH�ZU�iIQ�r�F���0y�7/���8�@ǋ3���ܨ�ZG�u��$��+%N4@Ά$��_(��)�8��*Lo*��D�|��c`���=�Iޣr�ًXeY��Ba��~�H!f�'�.���.톉��>x�l"�����ڂa����U���ΥC�r���w�B����%y����a��c����t�$�'&����j�:�)�eygI�37K�axK�"�Ey�k�7k^>��eP�3-��h_:��gq#ܣ]R�Q�4#�1c�Q2a�!����tO8kw�'
>i�oa���	u�Y����ĕ���k"U�tie`�������;�5�u=���+_���$�C�O������@��/���Q�h�E�J�T�Áqa���s�q�SD��dE��;�^&6Ը�#���d�$���>"N�,�̋_N�6�#���`U�g���D�fr�~��J��>ߋb��SI��Dp�&M���`�W��yyxa����ƺ�T�kOA �xp��0�QI��E��u�Q��$)�A�N��Ä�^V�p�n,7>�l�VtY���iS~�:^d�I�Ů��S�q�|G�pb�3�j�w����U����fW�����x0k�T����޾�s�~����G�Y��?<~vM����^�������r�:��"�?�]=���	,�� U#�Z�9����~���u�S�q]��7�wh��`1V������`�4T��d�G�� �.|#Kp�}��vp�����z��w��4m�/�H1f��@,Y��?���F��Y�xGJ2X2�T� �����P�1�����a��C�B$�7�H���z�}Tm�� �U�k���
d
��ֲ�,�c�?|�v�u
����-eX�M���h2������͑�~�E:�4���Y������#s��߮]�������iskV�d<���,zR�5��c2������lƭ���ɻN��:�o ��8�_�o�N�֦	�˫��b���d����zX�c��� 
s�����$�}ﱎ� ���.�6e^��������0;)
 h�Rg��i�k� 2c)��������n&��v�J�+�u�qL�~����e��"6��yH�M;��(t�ղQ�1�SZzO�u��=ʕ+��W��G��%$U��$eh����$o�4.�<B UqHa'v��33_}S`�XFDR̉Տ�]�0<ə"��ҋ�Pc�z��u"�0�\'��JS!>�̞s9� ���S�7LÛ��G��W��i�����oi�U&��_���O�9u2���u�-h'�.��"G�.������0l���7nV�}��;D��v�0) AY�Z��0a�s��э�A���w����Wa��#!aO`ed��-����`z\8���J���y�o�7���!�)���;wvB��禈jW��Vڀ�<|aNB#�u*
�
��8���{e�H����b�[��ଣIS[X <!'�ګ���-=lU��vO������EW�.F!^�O�|�(析?Ii��܅ZGQǕ�dkR�K�0�R�1��$���6�g���z+Jkl�k��oLYo����8�C��l��?ꍩ$VBT�+����z�a4��=�f���˴2jH�O�Jv�س)�ܬ�D��=�g\� 8���S�n1�?"��B�x�
�-�8:#F�/F�
L@MK��~3��nGO1eQ44C��㾕�k~P�PRG!��41�_���<�[��Cz�ۥ$q�u\N<���ɦ����@^�mſ��z�XDz�囎'��t�h��n|ݠp!������ݘ@5V��R�	ͱ������@LQζ���%��i�ۓ�4F>w\*���'N�|�4Vr����MZW>u'�9��Yl�4��m�U8wA�뮼�	�銁��?�� ��Ne���yL�Ta1 �����3Y�5σ��qvd\�������L����15��t��Gm�*��H(0�${���/��P�+ A���ʚ"܂�+�6D/2�T��S���p0���i˰�t&a�t�8�h�����W�C�R7h*e��f<���=������@0����Y�r�`�8Uw�&e�QH�����I�q�4��F�%`N�7c#|�����_%�O�;��Y��e)VpJE=Ф�|�E���D��R�����60��p��S���3e�;-��}L�ϾG��F� lg#�? �r9��e&�b�[��@5A���O���}� �ꐴ���0%���ʭc$�_�0���(���F&����ܱ��q| ��ȥ�D�� �C��7�:���V��O{��� �>u�(HE�m�J�d�`���rRpf���-0+���"�R�i ���^����:u�6F���5�G�	it��tq��;t��T��xvB�������I��R�zF(����
�n��W��)�̞���Є^���m�e����Nx���`7̰-��f� �V~ԡ�xi���@)5U��[-����9Q�yM|���=R�JH ��V�����'�uv$l5���Tϻ�Rj�U�Q#��/%�*B[�i���5�6�|$0��n�e)����Κ�`��|
�OY���t�zj�!�����<jvB:1)Q��h�V�6��Is>�y�$c� ױ3:���*�7f��S f�y�6@�A�6zS�N��U�DOU���v�5�f�^�`w�T\�}^��������_��w�>���S��ݿW`�s�L�x�L2�mY�?��P�8��||�%v�GZ��g۩���G�����W=g�L#= �(��HZ����R�6U��W�`TB���*k�	�ck1�8u}q��ݔ�<5��I�9 OfY-^B#ghl.�3vgsO��%��JV�6yQ|��%o��Ò��:c����S��+�£Y����Ja�}:vª�J�������͙%��������w�]:�<13 ���Ec���p�^��� =@.�2Bx�E�f뿉i_7�"�]�,����V�����,R�)@�H����)�%�0�O�Y莀�Q��[����[�	q�J�)_Vby���x��-�4t�>��H摜�~c�ׯ��t!L�������v`j�a<14&�sݙUF#�%���ژ�05S�<�L����Mo�;��ߔ�X�~���C�:�VO�u��AA,^(9�>�r͗:�v�v�հ�%}im]Z_��D�nY����ѓ}���	�n��8,�Sq�1��b�0����Q�7d���8�)n�piE�[8Y��>�KjgDc*ǯZc�ϟ��4�_�aϔ,h�U�i�̯��?�c� Q�e��v*R�g.�=��zh�ug�N���
�*[E�.���������ug	� X�M�J[�J�fQIb:��س�$Wq?ul�wՀ�i�-Cݸn��bde��4�
$�����.���H,�����.��E3��t�M�e�ca�p�=��d��P��h
�;-�U�q�a����XT^�!F���&B����tE~Nz)������2;=�D�m�xHn0�����6Z�M��Ӈ՘~0|�q�$�Ii��j9JA
����jD���ն5?t��ţ�?�!�^cˍ�^�ԇ����J'�G�K��
��ݮQ-}x���K��I^e<��u�"�W7�@#���/���|S^�*���q�>$�g��@�~�i�<�R��������yZў�q*&�!�������f�d���H<L|	�k�X��h����(��b���t�u���Y@W:�0>�"�gD���,�
��H�ru����8�"���-<��x��-�����ci���Xk�Mś��Jh���;J���3�ȟ����M�BB�V�a����Lb���d��^�;B�������
���g�k#�|Z2d֊�8&����B�-�0�$�6�].��x#:)MA�~zॶG|�<���w��_�̆��G���ײ/�y�iTT^�׷~	�i�S��x�Q&���h�[R����	���G��(��[9P�:]��lnʏITydy^.��$�V�,��6,�����8,MZ0o��h��m�(�u��A��M�Ձ�i�@��Gw�U!e>.~��C�ߌ��d�Lgd�+��¶�>=�ͣY���h��/gH�����h7F�����Q� } �.7Uh��qp^:��5R0����L��+�A!8�u|k�S��t�
[��~*0�W��>���zܰv֦�D PM>Trɿ2��d!�l�w��4t�O[�Q+�����y��J|;/��[_�����2��D�}�Ǌ��1OZ�ҟ��HH�rI�m"�X:Qo�~�YV�h%܆��(��ل^Y�p���R�c��JAg�W[X2�ߝ�]�B�{�L�����Z?3J'�(C���KEk6d���
Ow���#<]k�G�4g�}ױ�|1ĕP�qu+��ՉZ�h�6F7L��h��'���x��{�ҵ��
P�YXa�]�J�y��{\��K��f�]�$���(�4�n��vڲg�Z )|4L�]��@1��_,�*z�J�JT�-�g�+b2g�i�)��+�,q;7�>�$���ep�'�(PE%�.ˌ���e��1A1ƨԗ;�"���8�� �e�~�@�B/x[�ϵן���O��[-�#Y��UH���/W�<@L���2�Vu�O0�!h!g�xQ�qƅ2P!�t��,�8N�S|��u�v�':�G�ȎY=�o�쑛�CrN��U����:�.�|Qއ�z�E�B��F3�;�lU%�Ȓ顖Z�0"}���
2��Я8󘼲�l�ɋ����qA��k�[��Ը�h4eX>6�K%7Ďw��맗5��F���%�u`�â�lP��9l��}Ţ�qi?�7G����u��F�bO�۲HTϤL�������a����LS*]�<t3�ܨVwzCP��2ޞ5��i8&����Jo�����S��q��Oi�q��!��Pn�D�X���ϩь^<a�2�}�w�i���/r��\�J�n,�My���ي���� X�Ux0�k�g'Hv�3r6���afq�e���T��*���v0 �� 1I�W)�w�)�P�k�Ѹ0/���D7!4C���3��B˻��<Rt)9CԲ�L�h��;vW ��%�X�V� %#Ц�q�Xy�nf �}&�q����8�	�d���C����2�+w�5/���{dh�Ɵm��膡�s��Q��ջ�u����r5	<Gӑ���R���-h�*�D�)6ӂ��Z+f�i�*�.�R��y�i������oG���9�<�@�*�����}�~���g֮���� �?��Vv���h�u�R�e
f��ǲ<�Ӥ��iH�:��J�Wy���
�
�m0�I�����=��9�І���>��w��zkY��WCxB�2�&�?��{�/��	�j��}�`m^��8��vWL����k�]��G�&O#�/���������>'�v�c� eOܧ&d�T��+��y0�x1���x.�d������;]���~f�^dgImWÙ��~�s�y�G#�.�{�f�+�P�UX��~��0v0����n��'(l,�2&��U%�����5"�����몉��3l���XWB �o��P>S�W���qy<O�ք��f��k.�󶗚��*�p������a��v�<�u�����it�M�������74  l�J�Ѻ=m��p|�n)R����E �a�s��D��wA�G�3%N�M�_��>���*���j�fy�7:���Ў�P]�����V3�et�/��'M1ф�Y5��n+����D�Ed�?�w5a�`~%ay��l.ɽC�2����F�gIrKF�C+x�\�-�=�o�E��~�1J+u>΅5�t?��^����7|�Y=Tl*��O7?����-����݋ WZ��7��|�����T�Kc�T�T���z�VPbN����I�e�v�o��(�f!hZ��z�����zpr�_ɤI2������H������i�+�W�v}���{˽�rw���	��kM�X::H4Mqu�X�d��g&D��qd�=�d�B�z�@čv��D�2K��#s�i��╮:�4В���Љ���}����y���`T>�I��Cv���!��|�Z����>)2�̗MDaW��X6�4��O��[:�-����7��L�	Ho.w��(�!b�h�����V�P`��&�1���9�7�Wo1�m@�o��/����M�M�x`p]�n��	nY%�> ����>c�+���8�+��v�=�}�x�;�*?����N�荭h���^���j��lhag��2$ߕ��D��|��h���S9f��j�0Y=N�#o:�M�t�&�����p��_:�e�]��|��>5���VXW]�J�I�U�G�G��6����(L�w���)�Q�;���e��L�r��ޒ�_f��+���1���Gsݐ͞F2� q����O ?��*T��_YM�Jo?��L�ݣ	6`��<0��S�%4�{�I����qag���s���/����p�j�ڴo�/2n5u*E=b=.of	� �8]�:x.3��� ��ٗ
��F��ۂ���)�Ġ�&��-��T�6E�Ԍ�!�̄X]��`� ���q�b�,
fͤI��E�����u�fC���0�R0�TiOK[�������3��B�҈%�/&��f[��VW~D�)IY�y�:B0;�Kn�x�B�BR:�F:��p���>��]�[~�I���s��g�]Y�bJ��Pkz���ⶈ4H��P�5��	8��ń�Pg\X��	
�����W��!������Ӛ_u�n�����!Pd���#-��2��c�����@�S��@�Q��ߒ��ʻ�`��L��(�����~�z/��mb��.S)��藯40ۉ�A��g31-�%l��~�L�f��+����g�ou�q���?�tp�UB�X�BZ\�Ju�f���B)~
�KT]	�NYs��W8EqiQ=��*�)�'o?ë*@����KQɐl���P�6p��`��u�i�|��<I%�d�̻�z�����C�w�4n2ZjMIVw-�B�PKlNs��eg��.6���sF�0l�A�v����xT��5${\�B��Yt�4'~[�u�Y%w�4ń
Y_+Qu�-�'_v�������� �ndwӔP��,�S���t����!���3d���[�m�|�~A�!�@�e0Z��,�b�s[D_����������'��G\A���	G:�ö��d�Q�h `¼ɟ	�D��ur�ao��#䞿�?�X�w�235D6&�#��)KX
�G'����?N�M�BOI.�uy���&���J���+��-�Ơ�P��b�&/��Nv�7?-;)�<B\�p�Zv�nT�Π�Gݧ�ړ��J{+i�]	�[�S|���a�7�PN��7��	�8U�{��
K�.07'nq��?6h,R���"**��7;K�zd������{0 T�Q�EMD���:�H�Z�#��N�mc�����^CH�ߞ%�r��"�_f mt}�]�5e��>��l�םQ/3���Ɣ�wc��럓#!�a�����kE��G��@�1:H:��e᳢�%*K���wCQ,@��KA��<Z@��,�_d8;���o<�%3q��[��6�A{H��^�4�y���i���fw���/3^���k�W��J ��Z�c�8�RPA�P�4���T����~��	g��p�s#�b�'�����;�`�V���*�nD�zEu��}��P���
�;ߐ�0��3�R�>�g灌tG�ǣ޸Z]m�b��((���썘��M��&,d�=�Qg*-�*�7��'ZK��B7���k�"�֨�a�W7ep�΅�'��Y+��wq����wM�XZۻ�"q`� ��˟M0a`!�����n�/e��9�� *v�2)���yJ��/CC��}�Ϋv���#�\$�TK��#y͟�FC����\�y3�ʒZpYǜ��	z'�'�G�8@.lH��C;�ݘ��r��"��P�XG~��j'�T��Ց^,W���7O��}sщx��b%ȕ�/�=���W��
ؔ^��"�xhj8=�n٠��G5���v��&ѵ/�}�n����q��s#��(�'�P=�/���D��m�`AFs�7���q�j�&��G�9���
��n;e�(+
���n��B1�G�e�(Y�V���xo�B��K1�MQ�z���d��f{$s܁7�MAdwV�j�,��l����Ph)��9h���|����d�#x���Ok��IO 4���v��~^{/����%h���!�М�;�E���Jc%׫��G�b��Ƹ�����Rp�Б�.b��+�vz�H�z�D�ُ�ݵZ��J��ʣr��{�
��0�q��^�|iB$�� ۜ��Ш��KJ
�;������'UFm��ھ�?�HȈ�U����X�|������z�U�p��`�M���;L�m��D��!_5�.:-���;Iyf��K�SHg���zK��츾
ݒ4��`OX���\���#=r�K�;^��k���=TZU�	���@�SkG��1P�ʦ�n#���5�b�fm��gOe�}]sRfg�s�fE7���qj\��1��}(h��f:�b[�6q;t)�Ɖ6LY��U#���K⡡-�}�;�F��aH�Ø��Ґ�#��WS�J��~_qx��ۛ%2:m]hg-�N3fV��HD�,���,���#^���ޫ+�ù�A��g�ڄ�b̝����@�B�@K[Z��9�#T��LL�4����:�]��d�v=�H��Z�9K�l�okl�r�8LR	f��ٽ�V��-@y�3��"����!:�E�A�
��;*������ ~�'6O�ϑ|�'aH!����#��5�&��W�S˾�5d^%Ϥ�y��'g�����o0�a�j3HSY�`r�8�����O��;�[1
Tu�m��y���+@�'��a��O��T嵮&��RU��zS0!`��p�RQǻ��R��KM��C&�LU�t���K�/5�F�BEn����7���� ����g��ӆeS��'���LTؕY��vC�k�Ls�v}jg�e��h�_b(��=q)�@��Sކ*uZ���_��+/=��]�"�}��Qi೺'�������$�X�ݲ�f�lh�;������+�C��k_">0�R[���l�tf=}�,��Vy㽏X��A�u$�����W0�"��~j�y�ϥ޻�H���̈�K�{#WB��\�	���;�GSݡb�F�q�լK��S\�l�z�L#�#B���f�08,�vii�� QB>��Ȅ�zn�/'
�5��}�0��Lki�6gDP�{[��W�"��)�z �[�\��k�cw�(l� ��{�}+!���,�A@
-p�8:ٰ\nPZ� �$�)!�4|��QqK�٪4
�� �����S�'����|�9���\�n
�	��Q�O9�@��;ߨ=�Vb7�Dw^#A�AH�6';�>t:v�!𼡔��氒�]� a�ش������;�N1��z�4�%�6�a�hے&[�:~<�XqB5b���E���C�H�VzT}�!�aځ.��֍q?�/��S�S2z5(B��:+��=~�g��m P��0�wԫ���@�fL
��{�]��	~�>��>�K3z��^�m;��R��	�K����O#=�}�G3�1fX@�5�NY�=NA0l���4t5�P�o�Z8At��U�)#�w���@�ۤ8�4�|��w)��Kfݙ�4A�˚yw�b�#��؃������c!��`[ ;�/#C̎�I]���ى�����������S�yK�l�E�� �;%`l��l�qT�W#�we"�\��7�֫���: ���(R��)50\7nn�!
"���p�
�T��f�9}×։���-ނ�W:�ۘ�8��VL]eh��t�^ ���*�5��ې�7�K�IÃ����������v(�N����n�ɇ��W{�D����A�E�Nk�@�G^���\�"ҡW����s_ Eu�W/ż��Kߋ��/c�m����y�Q�)�wl�q���܊�OÊ~8w�/���L�E+E׹����_R��K�>���vOL��0��J-5����ks�L������COr�T#�K�	�>s]���|ǁH��$$�^�/���f�:��2����/]������E.6���C��Z]�ݥ�^�Aj��a'���/n�(����◡聾rK���uOd��i)�@���V�Ό4���urD"E4��L��ŋ�����ݞ��:#e�1��=���|�����~���]��:yW�����ң{W�P��<�#Oq�v�~å�^/���;Q��V��@�~�h�A������i%s�F�a� +�о4��lF'b���m[�^B�ϸ���(�B��7V���B�uI�8[�.v8���� R��ba�͌g蹈�e�F�?��Q�,�6�� � �~����%F;�L\5�X���Jt�'�2��[t�TQ��z8�Н��:���Ua噁��^J��'4�JG޿'T�G�a0��l���^��=��v_z�Pv�c+*�%� 2�)�`�!�*}�l����&��M�< Z�;/m9ư����m^5�rM�p�Z��C����ػ��l7N������o��BK����)cJ�F�T��*��b�:qr�xu�-�wsĉZ��;1��*v��NUnP���G�}�E�d��N�a���c��vdu����д�q���=�� w������jo�O�1{� bwr�=��"�PABa�4B���_Q��?�(��:��d]�����x�b�yn2��a���ى��r`�v��Hk�y)��t�:;���]���t\%IC�K-�����u�MdY��� ���
2�2��Rf�I���]X�����F�n��d���MrA�Ça����h��\����6e�];��LE��Y|)�W*X�A"�MX:�C\���OZRj��V|�u�Y�1��~�mZlP�3�v��1�X�~`x�R`�]�~6f/��&z��o��x-�)4�P�!Y����<ޛ�� �[ou�YW��9���!�,�z�C��Qw���%(�fI�L��YS=�Q�%�E%��r��d�VO�0jN��O����r-٠e7�ؐ��"��6�4:�_�QŇ}��$p��40����݂z��r��n�2�ԯ��`b�C�&v@puE9�I��_dŮ��'U\����y-���=B�(��d�zԿ�>{���N^���\d(��sC����!)$d!�`����:��e_V�5�xE��B��b��$�Ӷ��^�/����V�܏!�f��î��K���Z	�e08���VM�[z��Ha��o��c6�f��gǊ����l�7�<�4��5�����r9
����k�	���*I�/OQ������1��lX��(�^{��>��YDx'���6/�#�2�>
?�3����2렛=�����4�_��o�X�hŏ���Uw�P=�Hw���v� Tz'�m����1I,<�N�H��������<�	Ą\.7'
�������=	����l7�6):�d��1��b��ş�Y��n�H�%��zs�A�zY|��n��O�	t��Sõ�z����h�}�r�ؑ$��fһ��I�C������*!n,��Uo�+�~�	��(#��ū�W]�(,��_�����渢��ez��.ŸI��H�-Fr��m�]���K����ۮF����!�����Pv�̈�F<��f��-�Z3�<�d<G%Q���	��eE}�)^�Dlu�mģe3:�@0;{y����o3L�
i�o�4\e|��ߠ�F�?�#d���Pf�J���9�k��/e
��@��c�#��HK�CH[.�����]��3�֞�=~�f�$�T�iƻ���D���B՛��5�n�hpU=g,����嵓{���&̠1����YL���f\%��٪�&@�XO[jO;����M�����Z|�=q����BVདI��ϗ��3�7Pb��s�#�
�����w�Q���0���NQl����ķ[�1&��9�8�������oI�W��r�E�82�{2�z{am��|���\�_/�'�n�L5b��Y���} N�Ov�R���y<>$����o�u�['���:��S$7IPP�������P�o�㻪�jF!d\�V��\10xD��>L�p�'�$$�e�2�9=�h#R����X�Y:���<����g���1ȷw��Α�J��P���%y��������?�����#����3��3v����?>�k�+�����?�"�A�x#�"�����S?�c_��n�s`6����V)$m�ݝU�5�eYo3{���?�e>�0C���(��_��JLuD��˰�H2;aE�\�Ql�����z��(`<~ة<��L�Y S�������u�ۑ�XL��cMS�]3k`���x�<h�����:�4�u#�ֳ}���C��s�)@�}�S/� ��0���XIZ��4YMd���%E�o/,��#"�
�/"�K���t�*f�=����`�!�����%(��/X�w���)����֧O}?�PX�w "$`�� h*|_�5���B�a�Jo�
?&v���5I�&A�a5u��X�=���q�Q�Aa�җ����q������k)R�X5i���/���V-g�l����	�rR�E����l�:����!o@ ����]�X�+���䩭"�c����w^��T�����|�uw��)�������!�t:�Ո�BZ�~����n�@+տ���n��˵��.�Ӭ�4dU�h�>�"A*����r����M��Gc�+-ƙ�gRN�3�l�~�D�5gUaK�+���%�uWs�۽8��I�^=W�����9�5D�e��F/���Wm��繏��!!�ʲ�����7�F�Z	��k�'����0^�g�xC�y.�F�����t�g�&�f��,�#jڮ@^6��\��]��t�v6��?�[/�b������0�?�m�mݽ���r�"�#���W����1���W��ղ��b���B�Ton�'�P��g�Y��p.�B�����fԇ��$XEA�+��"6Ҕ;;�&�oaI��N�T�ڈ��$V�d�{�.Q/���Ф��#�&�����{�x,���ͨ��Q����U
qe��{�|�9qt�UՉO^���(�*f��Y�z��x�s�_)�a�#֞>�oڜ���I��㉂1��LM����w�x��xT�iM�M�����՞};Ў\=�]���^Z��@1Zp3�R� ��.�O���wn�2F�Isd�#�OcʹQ�k���I�/'�/�;ׁ�N��h(�%C�!�����Q���"�#����"�NӗnJс�L�ȯ���f��,�����|0��n�y)�ig�����:��ݹ�i�5�ä���NJ�u��T<@������3�Uц-k�����]k�Fg�_���?ȼ�[�@I
�(o4�.��}��a/X>�kx��Xu�h���9�vׄ��%.����no�ڇ�\��?�؏�o��y���I�����m�ҩ��Ɨe5+��d�;$&8]m��p�iE&a�&��4|�G����z�/yZq�:�^B^Z���,;�f����,l_L�3 p Æ�RqQ�tgչʔ
w�@�)J����~��L'?� �ˍ��2�xY���>���=���иV#��c�1�Ӳi���}ݲ&<I������vZn4�p��]wPU�r#�Ub?(:�lA�a6I<S���i��}_��G��r�u)�І"�C�����9�]��P瓊�.��j��7��bN2�d�YR ��!jZ�N�V�pȆ,_y�M.S�0�"HzG�*�,N���R��d3���9���q%��'C���<�%s8������Ѳz���?�2FI��Cp?X
*�	h;d��8B��F�ն@;,��Ϭ2�0B�&�@�/t����<uu�O� Br�k��$/��X�!R�q5�3S��[k�s��8W���Tx3}��C��9$��O�C���z)n(L밆)�tЂVi(PU
w��vF!��Z��f�j� ������I$fr�V+Pb��-���ဝԗ���F�6�����������]�yiӻ:�f:q��ssZ�.���F�c؊�D���U*(�nR���+�"���Ώ�*������՘���9�R"�t�Ή�Ϋ��{�6S1� r�:]�H�����ku��-[ӹ�G�i�q������>#:`�)�}�L��#S��O��zWY�-u�eH]'o�	����kX/]�ʫ��Y�����E�(��	�V�B�eC�$Ad}��K
0��3  ާ�!��^��ދ�@�t��Z�Bc�8����ZsL�n#���Y }LUu����aK\!ٝ�OX�&��p��y���=b��.}u=�FH��1'�yqe�R ��wU_�\�>/K��N�5@�#-�d3Վ�L�4��م׼�yXX@݂���h���/w.�]7�w �⫲�>y��J<z�F��ȱb#)N����>HV��myf� ���{˴N�!��
�7���;B��]��
����բ5̦�&��NИz߀[�>n�=��a�U!iR����G��9��VF/�bE��(x����2O|�]�'��7�%K:uh���e�yl�'�
��?�6$*Ȥ��\��U�J�����C���-vֳp�~pY���hҎ������d	�G�_1w�~�ɚ�9ƈq��cO,I����/K�_�@g�f�%���ZK�2�'W��@�d$V PGmƱ��1��ȗ���F�}Tߖ�F�٬B����w`*P}��d�]h!"ۖ�!������4E���N�p�����4�ᛦ
���7n�R��	��C(�Ɵ�>�aS͚�d&bPT�ln�m���C�^3	(-+^��3���t�c�+Zj��	[_IS{�`�:( Ɩ׽i��|�W^}�	��FE}r�e���C8��[�i[g7 _�xѧ��8w�;w�Y����6��I��iYЛ>���L����G�{_�œ-?�.��K���F���z$��j-*���BY^��Pr\��M��*�J>TA�J�掠#��&!�H�G(��*�� y=�:J�	?��k�3@.�%^�k+�����q�<�k�d�q��qn�ַ�����!l�ϱ~�AYe��"j����T���T	}��et�bU�sۨ�y �0S;ne�"�v]7�R�͝T�V�#�ӵ� 4�6 ��\�!����#Cj�߱�+����o��� ��:�ճ�]<Nc��/��L^�h�	�c��n��n�c�Q���Ealr���������,�I��r�Q[��[aM�/�"6���O���2@%�8��~��0�JMOT���?��u�,����^	�	=����a��pN�ޣ���k����PZߋ���%���۬���G�z;��R�b�T���v�/T���`�n��ͮ����ty�`L�D�2N�"!=S55���K�;��'y���R�0QU1Yw�7 ��_�!��K*�����ԭ�,�z�A�L�ꀍ��d�*f�\�:��W�y�(��m�����IM�㣖�,-,���h�4� �O1h.�BQ�;(qpЅ�TpT�Aeuf6�eKm���v�A��9�ZIA�K	yPo�^�ߧX��k����Ƞ^��A}V��S��8�͜����ȃ�q��.�P�0Qg5�Z�J����Ơ�_Zi+�D?f�,_���|�A�;J��X=�W�S�;�'zeJ3�Kb�����O^b�U�&� 5o'����6N���\��,���&^g�K%�8wS~�]������%�c]� n�օ�8x������?�o
�򠆨�J037噻�k�	�3Jւ;Ԅ5NwG+�������L9򎋄vϚַ���6-Y��R7N�y�g���/<��'\�Z��/i�@�x��~��	=���4d�=`���R��O'L���}U"�Sqʳ�Id�~ A$���A�qK��Eٺ�>rC
�X(��nԄ���աa�����U����.e%�Xj��J��V��fZ� *��K2ޜajC�H@z��4O�Q�ύY�����j
k���~���KV�&���WL�1qo�@DJ���Mn�1��]�P.cLFF����}R��}��h裗a��c��e�d�9pN�_�����v���F���x��0'՜歗]�TI�h~�����faB�=��<h~�x薞	_נ��N��J ��.n�L�{!p�+[Ҫ��D�[�^�6�4Ȫ�c)��
AJɿ���a�D	W����_[~EH���G���.�D��!�����k���F�`a�1.+����ǉ4ƓߗG��Ds�6	���.���WY
��Q�Adp��,���+ ��.L{���.���`b���Nňtȣ(�Q��/Z�T7:�ya�u��~ ႟1~�V�iCEU��1�@@��)���Mx���,�����\:��I������<w�.���+!$�W[?#���ڔ|(�����Z� Wك�Cڱ��;D�O9��;�a��ߊ�@H�����	'�Z�id?�⵮V&v�5C�4���$E��}�-�����1+%�}{2=�"3���t���{�o����"�S�5D�P:5:���'�zbUhtN��;:��>�B����p
VM�j'��O`UR�Gзk������Z�?eR����`�fq�����}fht<
��w�%+o�Du�UȈLVԞX"t����:#�k��oh����Y�1�ÉX4�L�����̞Y���@���Y�����S}���+��v��(�o��7u�bV/����xm��-p�^h�8��� ��$�M�
nK��g��>�&~�x6>D�/<~��-�����b�$4��N/@�v�Lܩ�e��B�,mZ�^�&V}Ժ�ˍ���S����m���ծ�ކ�/!�D������=T����D�e��JPWkT�{�ko/<��>�t��2�"��E����ϛ�"t��x@���CMx�|_?��'@\�����T�{+�~� X-g�#I��J~0��	x��VHgn���B�?-�*��sl~� ���jȠ���I�܈Cl�ȴ��"�1\+C�l���Z|���<3��7�酴���F�u7��i6�>  �7�e����g��! Y|fJr��
�j"j�J����Qӥ��7����#�q�0��@�r���H�4�E�6�D�h|�D"Km��a���n$B6�M�!}���y�C=����β�]Ӎe��4 R�]ɩI[
�!�103�#�!:��#�V�+d�M����z�aā͠�lc��Z�g�~@@�Gz�'�sX���G�H!.bJs$8����g��������p�Y�Q��ȟ��
1:OI$:�Fˑ <�B�r,���?���B�P�L9v���0,�l��٘�V n�� �Tp{h���nbr��u� �^s�I�AKؾ�ܲjB�9�?i�` R1�'���Ec3#�d��np� Wj[��O=ݛ+��Y�1�g,�Oϵ��ִ�a�9�R^��,ʶ�#K�[�g¶�8a��C&N]O#��dg7_��
!D�ӷt���ܡ�OO Ⱦ���ˍ''+�:y�/��Z�'��`dws���w)l�s8t�%?�}�q���-Olr3S��v>�-x|�$_��e��R��1�X��~�xdj���
�����/�͎}%�ݵabK���\6��`۞�|��m��}�J����'�a-�M���R��;��+ּ� d�Pe�	={��X_������؀��%�P����v2}����0���^/���zB,�.���6;B�F�����ӜY-/^ͼ��Of/'H #s�{x��iܿ�<ڙ��_؝�����c%�#������/^޷��TZ��pd�Y�2g�>�(>>����&����H%�a�����قl-@S�����?'0xF_�򲕴(��f?e\(8���K�j�ėk�rk]��{ղ~NW���W{�*&��@��`�A���2�����J�rj�h�6@5I� ��L3B�.���sz�(��Խ�8;�Np�3{�|�0ՒԞd4�<����f�]�2�W6���_�'���eS~�Q�Q]�{��>�U�_�JZlN�o��mT{�o�i**����S��th�=���=��9^^�p֫��B�
,��jTI��u6��`˶��.��WJ��\ D���~��őU�j0�~�T� ��D�`�,H�t�|M�;_0������]����m�3ϖE��>f���H����P������j�)Q���:m8��'�W	U�+kR�V6t���z�W���_�x)�����]W�;�ڗ��I�FZ�)�^�&��|�����ߐ 0	��s�n�գ�6?k�M4iدQ�aT��#�Ps�����떕�K���Ë\^e�ǿ��<y$���=���l0d~�*�}vW����:^��?��!�k(��C�Ҭet��09�pwI#hAk,v��?�-�.�Q/���/y���
i�29����1�N��*QUc���#���f�!���(֟m�B��؇����
�xU>8�D�O��||��AZ���Z1�9����C5�x
�g����o�2Jd�JN�� ���H��v�HO�����@�����K;��pt�� 'j�4J/C��}����Ƹ3n���5N��^&5N��kz���NK�T8��� +��Q�iA��P�i�W�Z+ү&; ��-��7 W΀��Ҫ��!{ӄ���n;����mt/v6z�Wخu�䀶��V�2r��U�r��%���<$�a���`�>�(J��bp!JӓzqS"��o� {��z�3�c��0~yzn�Q �Q�଼���n�~Uf��M�^��GP�H<�O�S�����сSW�6\5!�ft3�9��Ș�K rb�̉}b󾒰fsH%��%,��=����r��!W$��&|�A���*�]e����Պ���a �\ c�th=p�[�!N�'/7w����_� �A�ֽ�T}����f'(����^S(Y(�, 9P�j%����H,��w�k���Y�x�� ���T����t�_Nr{7��z���.���WƄa������s 4�L�@���aP����9�,#+a�-� |c��N��)����������F���b���v�$t�P�Rn��]�UN������n�q����:��D/�}���ʸB �3�⒲͇'-;u�G�٠� �iX=�m��T=sRN�a�2�__��RY�M�0�����6y�g�/�Ӂ��I:���DU���/�e7C��U4���x4��"��ud ��J��c�&A�7g-7�z<���?�G ����3���^[�M�DeNK�%�ƶ�2�M;����5LӼvbʃ>D'��nK" d�]Ih���y�#����CY���*r*�.�3p�!a��bB��J/#L��k�w<���\�b����&,�iL�<��z��?�PUצ�U�a��e�*T?\�@�=�Nɺ~<��I�j�U��0�z�v��WE�-o��(��c��D/@��J�f(������a�A���V����r.G�0`-��݃s=H=~��T���	�y�J�/wI �*zI��yP1�݊5#�b(���R}�53ڱ}�b��@ҡx������V��H��	"�������>��m��2\H/V��AVCm��4Z�3뮯K ��,c��1�,7k�J�SGUP�t<��F-?���V���W4$^��B�bMPn��(p���=Й�fMֽ��O*y�%�D��C9�F�ٯ��:0<S?�9a$߀�>���A�`Mz�FǱb��v�EF� ݯ1��0������KC{D#*c�xu����ы�b�Ӛδ��`sLF|��$�&š;C]��D�������{:T]�3'Ɏ�HC����."��e����-gg�VO�K�����(�-��OA�Ɠ�UN{�u�hF�n�ƀ~��_�pJ��sУ���Uƒ�h���*:vbJ��V�_��;��>��(5+$Tl���|�y�n�7�+�N�cwd������ݜVr��;ty]��o��2���ܿ����c:3�:p�d��In;Β㈱�H�������|>CU��H�!��s'�x�ݐet���_���E�Z�����V�<�ge����6\!����u�4`����~�ܖ޿�A��)S)�����y);8+%��}�4��g3���G89/x�
�(̛:��<:�mt�
�)���/BZ��B:ʥ�'��oȆ>#Y��"��x:ϗ��fvj8=D�7L;�F�c"#t<ϦpaL� �&!����Ά�2)���� �:��i�k��X�Och��q~����ъ��?��I8��@_�OgA]�	�8�!qdƫ��k�������_H�Uh��6�'�r��#�ݮ�́����O����cgk`b���i3������>A!��ᴝ�(�.����S�^��5x�8�G:�XF�xc7�y���+�pP��t�x0#��M���h��ɡk�v�u`d�m�qW������'�#̍��^�|VF���=���l��x`f��_����8�Q�WT�9�+�#ϡO���!e�(�[���r��p۝݂ �y(��R֒j���;-���(o9��y&8�A������O�Є�X��S�-�5���f���/�	[���j1
�3���'��5��Y�?/o��ͫj0�YG��gq�\+��L��Y�"�0�0��d�F� �& �f�`d�WM^D^vU#g��K��Ț�����P����^qÚ��Z�2��0�j�6x�"��q./� F���Go�F�	ƣ�D�bv�ϟF��Ԁ�Ym��5��� j�T��fw��&S&���˻H�#0��Re�e^l�Olm� ���:������ ء9H�eA��c��?���+����eBE��ծX�n�b��9i��:��{Ɇ�g�Sa��-���%Ӽ���[�(~�SmCӲ��a��u�*����-ܢ6%n��'J����678zZ[jQ��`�~Q׺F�K�[�o����Xj���ɧ��Cwc���L&�D��m�U���`׻3
[+��
7�%m�)���0�H���Oz1���K�X��
���zW5A����K� "�^�����x�op�$#�D_�G`��)6��/��G
���]
��W��Z\l<�Du��a"r����S�f�P���ځzO�#�)��*�PC�hre~���!�}t��&z�z�{�r�5����] ����C���flaNJ��e�K�m�P�B�E�4Mw<��S���_���!3�OV��Ĵ��\[��I��E\�rH�
(5_�s����Y����~XHY�:��K�쀋q��굱O��*#�x��2?Y�神�1�c*��ι.����P/�pdC��S�Ȗ(�08��b�R�.'@_h����c`!�[��6o{��8�q	�%���y� d)�O�)�F���+$2�p�ݑ�}<Ӌ&W�\F.��%�λ
� ����e��>	y �s0����|U��^��\^~��sE��[ܼ����d`��Z�,/l_�����'Ѓg�����i�#�5Y����R��%�d Pr���@8��r
3Ԗ����סj�+�wO�a��'��t?<�yr�Ҩ�~�sukQ�	�`�ˈ�H�}���+^O����'��"�uB_Q��ʸI[ d�<#|�e8x�^B5���c,<����*�sxWJ�=3��8����!,ʟX��i?lsg^I� �c���e��l�RR�9 �W���M ��R�tQSp�+��њl��EI-kxq�DvK�3�1���?��l"I�y]A�&nL!�����>7@�7�w.����І�^���123�ϙ�T
z���$$�/QH#h56p��Z�s�׀��Z��e������y\A��V[��b@�$�����故�	N�Zݬe�!,Ggc<�>�=ޙY�w� ���h�CT:������0���o�W��;�<<��� S�3���_�F��Ꮈ{WCGA��7�ƚ���YN���'X�Ņ�w�VH�o���hi3�0��|���b�}�5j&@oX ]x��������Mp���n�d�����dk@�M���]w���WM 'YL&ty�F�]X+���c�q���3|(���3�|���UE{q-���뱉ᗐ��+�aX ��O��I�0 �����.�����'�W��1ɏv��	l.Ѳ��Lw$K�A��uM�ˑ������,��x��ndRw5���a���pA����5u����A`9��&���Ω���AF�����!$u�9/�Մ���"A��a��Z��z;�F�X7�!jvf
aMXNvfL_ W���R�������S!Q�F�;��S�Ds��G.=�ZJEu��*;�/��<^����A�� �2N ,&ɼ�QzY�*pq)�����Q�r)�������ƴL�F�R4��pJ��0����0!�_*���_m��=1m��8Q��"��t9�h���ҠΒ���3���]�������[�D3�c(Ee�Ҝ¼��ؐ�rE�4EaJ�:1&!���7�(S��E��@��Z^��F��N�Y;�8A�<�=_ߴ��D'�*u����P�q0
�A+cV.�����2%olNb���T�1�8�EL�445�K��t/ۥF�t������J�%����EI3�y�J�h������㈽�I�i�z���w.T�	#��=&�����%�+�d��/2e.�����<2Y猖 UO�z���#��љ|$��.��Z�rSkFg��+�������HN�l'�2tBCBW���4�b��� =�X4��qυ���7u�8�[
�%O��o)? 	=1O����m�P���R�(H⿤�I����m5���4�a��O�b�9P8�-�g�&�}��`F��tZk�4���|�hBX��s9�71����X�У�^���`��Y?t�@����y:�XĂk��v��%֛��xeD�+X�]F�������þ�#!���;�w8�^����3�"މabP�4��"q�V�S�ж��w瞚1��AuL+����(:`hkj#�o�P��Q]�F ����D���$�G��u�<�GX������S|�˞~�]���$��u���D�:�!��]ޟt��W�B�ZB2V��<G�ě���mɛ@��tJw�b[�����a "׳��!R2�EЛ�Ϲiu[Ţii�VU�c��qq4,��_r2װ4��0�&V�{˨p����
��Lq���^r
b�
���HL{A�{mdy:�|@Lӗh��8�Ӕ˴t]��2PD�x�OL�3t�A�U���MOy~��B%���O3*T�h��Ƙ���O�.�rb�ez��^�~�r��C	��gFW�;��-=>�i*D������R]0�gv�N؆�[*��OzS�E�����"b�t���g{޿��x�1��\��%#B(��f�y~}Mw��i�7�i�[�+�Uk����T=h���)��ьw����������E��Dv7(4/]w)re˰4x��f�i���M���X��6��g�`�h�Hޅ�8hd�W�ᨕ��=z����H���L��{|Ћ11Hԉ�=	�x �)gn��i�t(�\
��\9�T^�c+y(U�o�/��֛E7_g�[�SWS�a��@(;2C�J�S�tQ笨�[���vx����'N* {Q��eu���gB�tق"x�]����ҳ߆vӹ���ΦV�<�⍇7��˰
�O\N�}����&�*8��tq�sb����VU}w��F�J��ع��(�L$����U�����䢺�0 �ê�4�"G��ӥq��hV�\���?������0u~!Sn��]�ѥ����_��␳����Rq2��/lX��\?�tu�}�0?��7a�]��zhO��鈓O��;���IPx�'L�'$�X���$�a>�����T&��@��R�ܢY���j�B��������.
�V�Ϧ�ё��;e��ҷ�l�'w���0�q(�߯�6�0�Þ���U���_����KǕ�zAMa�4f�B��_~��H�>�r2���T�)�z����J}�Z54tP�w�2ŴZ,��X˪w:bm
�X�K��t���������J��m��F��t�w�4m�KsD����L�îЏ�b{�ҒOr��vG�K��-P89�ħV>��m�N`�����B�-[:!����ҿ�m[�Iv�KbD�S���#�2^�_NYf��{S]�\3�c�?�w��[��.�I�w��ix�@S��A��i��=�74��?�EKv���R�`:��i�"=����;��9���0�Q�T}k��Α����"�
L4�ХL{�����L��������bET{~�	u]&��{�X���y��C�H(�IO�).�8������z/�v��$�.-��^j[l�CRa�#�햅)yO�N��,��e��m��فyO"�`�MZ�^@���`���֋f�-K�4^��{��С0�8
������|d�ݞ��1�Ĩ.ԇ�����K�_Ϧ��V9��2u+}����{�d�R|��Zۧ31��l{�%cĄu=�|�p�4�';�(zrӿ?Q�0�W+pÔ�[�Nq�a�v��dRBg�����9�z@@�>	�OPmb�6?��/M�k��H<�З6��θˡ��0JJe������ޖCLr5Hu鑾�4����CF��f�
�VE�&�h5�Ti�E::޿�����	���G�M��ƴ9M]]�B��N�������#���X��JWR�7U���0܎�/`��T��,X���έ�_���z���^�ɃE_GӀ4�E� ^D%�����s|�\9~�Q'�F������R�0�#Td��Zڐ���)r��y8��E1�YE!"�~�����V@�ey7��rIGy�[���!S�5&�j
���*U>@i�/�
�G4-��g���8�Y ���:-��rN2E�� �{�X=�\Z��M���"X_F�a��.ް0���y�Z�R�B
"���k�2잺�iMkt�:��.cw�[,����
*��������Iv�7k���	9?~N�e��s;�zS"d����DTSC4����C*5q^�`�q�$4�n�0y*�`��S�1��������	W$�A9���\���S���a����Rz�Av�bi&��R�܍7ػ�!&����Z�k=]�.k�..����-r������K�D̞��7�F?�ԉBe�y���w�O�^���}�v3[�V�h]��T�ҩ�����.�,�r�)�Q���/��x
d�p���Ŝ�)$5>ERa�L�AW���QA���՜�1�H�a�ed���z�w��io$�`*�.�-_끩���!�icT�	� ~��a�Ght�*��*����Z4�O�3J:EӰЯ�{�*�ؽy���g#���#��~�j�{���Ҥ�Y{4�ޮJ�_<���ż�!�$�G���B	������TbX������G?��O۬1�S"���;ƾ4IN'S����|����BM=bD��K �0��U��V?E?�ف��O��H �>'&�+3|_U��5��hz�^�]�yB�l��#da�����f��4$�� �!Ѵa"����g�ȭ��W�߈�nh֐��U'l�|x��\����H�1��c���Z :�+�V�=/>e�c ��Q�]�]�y�*Sk���{ �/Ad{'���>6�67(�5�K�O�	_9)��!�7p/����;b���,Q}�'-���c�b^�]�@���/��뢳�𛰻n4_��~(s���d��s]�2���t;�:]�i��L����D�`����j0�$ ��_X�`T�*�2F��[�B14��aZ��Vix�]3m�bt���"�jO8(�^�f��0�w9�xLW��obu�F��)�/M����RH���u�� �V)ϠJ�N�`o�Ѕ��Ș��Rl�@����,NZ�W|��ϊ��V�Y]i�ϼ�c '���O���"�f�����:v�p"��|�$��7�*��;�pW5^�U����<�#��q�ebx�DJ?r:�3�=���V�r�O��&���VՊ�}]W\�Z�}Ƥ
DF��|�g��|#�٩���F'��=>�w'F�7�i��粆#���8Yۭ��g>��^����`������E ���alq(���\��N#јt�unL�����T��1u�8{��m���n�t:����c���RvP���L�G��]$XꙸI����R��?ԥ����c��t~(�s$�C���=���B`&���Z[�H&Y~L�JF�	-�OD�Ԣ�A�݈B"$1��D�,K����WR?�-���_��C2�F�4��F"�<���̥<	�q���ɦ��]9�:ߥ}~|۞��)B;����(5 *}�*�JA%[����є���'��*�4�*owE?ﾛb9��ً����AiC������*��6Yf�.��@[����#�Ӛ��l��� O�+e]���|a|���"\��e�Y���1��5y�a�1����ɽ����0�nw�:�/�UfR�פoMG���{z����xz�a���n��6��x)-��R��eM�x�[W�<.��yF����7h���* 4��ET(x�/�.��xƔ�5Js��;_:�Ciߛs�"�0�0j0�\�	m��]����f�`��/ߑ{U֮J�����o���C����O�
��I���?�+��Dظxa��9����u4����G�~��%$��-aaz�7<�>%-^@̛�uL��<F ���Q����_73�ޜ�x�č$�σ'Ԭ߬} ��y͏�W��i��0Q�@R��3�=���|5�n㖫`��2.�'Ķ�΋ɥN�S	�s��bQ�%���J5X0���O��Q�CP�������	�Y6k&X�)CY0=�x����n���sHc��W8�z5�p�Yj�)����be|���hȍL��Ps ��U���&4��[)�!�f"�]ʶ��v���y������	�ݿ#/���C�w�������ds��c�] ���;�6��:���?}2�C"�-��n^H�(M<��J26av��j��}m�B��w!���c1�s�����0�k܏۟j��]n���o� l���+�
"BM{5@׀����
�r�uO ��"ҥj���ڢ~��2��r�	�2T @gm	�#RA�X��r�����#x ʫ�0� /j`���C��7��N��n}B�%Φ�Hh')����4�3���n��5SHf�W튽��/�b��Uf���p���y�9��������X���q��2�ֹ��~������A���5�C�
���2���B���L��IΕ�FވP��rt�ۆ��z«�{Kq=�#�������EX�%�2�X��M6��k�c]5V}u��:��h1�/�p�K5��@ m_Q@�y���NC	i�m���G>��ͷw��(��Q����l�dYʦK�fu������������(�4�������V�GpM�J�WW_�]�3��59ɠj�~�oE� Tܜbd��G�#	������6ť4�����-/Y/ڦ���������T��I�����~�Wܗ>S�s�/(/9;��io��٥�q���F���!6U.�?�����J���j�Q�q�0���2�n��;�f�/��Cwu�k����׭���;���֨O9�d�wB�V���M/vݶ��A�yz����ݚ�=հ��W�Q㰿A6\���3O��J梵����R��lRk���P���PUvF�d��3�k#�MU^�Q��YCܔ��p�ӄ���S�7���E���B靦���/������ʫXNu�LT%�	2��Pw���U�V�]ϐ�?�ڲ� 	l]��q�*��B�a�.��FlA�f(@��i Q RICO�w\��s�<���U�t���7w=Ҁ��k��k�M�1ʮ�ձ��[F2���Z�u�E�+>
���d����>���Z����LJ�^Sb�%�Ɂ{v�"P'V"����[^`��-5��XR=���Luz�Z ��3IC����2T����qq8)1/�X��L�9����`���k�?&���oe��_�|�b��4��(E�����B��2��g$�6�sz��FG/s�ő����O��O�LoSa��ey�͚⪰���|�@̷؆V-��x&�U���9�S�xf6�	���/�wNjhj#d�������D;�ݵ����Z�`�j�$x� �݃ۑ���)1P���mˍCIY��6��N!œ��ϛ�߯�(�
��i,�5 e�V��*����M��;^E�B��/�{�����9�� w��>��n����V���}Kj���APlZ��ަ�u,��95����g��?�h�&���Z�ګyH a�u�1ח)�su��\u��?�Ƚ�B�z��ӆ�^��2�X$�k@腘��.i!C�o�t���4���Y7��D��lgW&D�|�,�1W��}�
p^fF�5l�t^�=���EUt��#��@�Lzܻ���ܺ"�l�ƍb�gt��+�y�݂�QMŽ��J�K6e~��oܪg�^0B2!�Ɏ���޿�1��z��Hc�\�n^��a�T���.�ЛȚ*���C�F�7!�0�P�DT�,�w�ѳ�e|.1��&K�H6T�B5i\�i��^
�E>�cּ�]	3��m%��������Zl,��;E��ޅ���ʋ�[ǚ�$�~h�Y`�[�+�Ir�-J�f�?�I�~��@����x��	CPROܳ�ǌ%,��s�(�_x#������[���{��<��S�;�%�jwP�y\�ԚC|ǎ��bLf�x݌�:H���Vz=:;X�,wOOZ��ĝhRsW�q�9�%���`s�l_��@��=�$J��V{/�k�Y��{A�U�@2����4{� '��E
�}�����	p9ð�6?���=6U$rj���CJ��0�|�=���.̨r���7�LL��"[>��6"9����zŝ%o�8E��龁�� UJ��w���iE��V�<q_�Y�9|Emnc�z�e���au��m�[�ɩ���|7���h+W�g���9���"��oLx*	�R�JqB��Q�
��Vf�Nǀ?w��R\A�y� �>3���/-f�t>1���$�rm^4�*������%��v��t��p&�3�;l���]���9���5_R�0��Vh��i��!|���.�N��,�P��T/7^�I�N��@�2�MHWZ���*�@�����%����8w�^S�ދ�� Vh�A�b��O�K�j��-P\�l�5��[�F_1�>�'����/�DVe�SA���|
7�f:�����/��5@�r5�lx*�S��v���%Y�GV�i�<�p�h~K�a�,aM�%[sf��������0��O(Mae�bÈq))ȣ�D���D��'av40�`K��}��w��1��_C��+P�J�iC��b���E^����u�B<�x�$��&��*I�%��K
��f�u�����|��dM�.�Qr�����f��w�J�x,��4�ysZ�YuT�U�(}�3�&̨�((�%<Uxf\EA�5]��0AXM5��HI�up���%�ڨ[���,n�������.?X���}ʹQ�$�I�:S�Q+�up� ��#��m� �^�����ղ.�[��AN\@FQ���^��/jL��< {�h&o��d�LF���c�v�c�ˈ��"ZL�T9_rD�]rF@�*���P�]��꺏�n�93Q����6a�T����7�����ǩ��:�wԫ��>k|���7.� �v�P�������i�J��2���eCI �ٻ�jk@#(jn��v� E��1vp)���s	�����t��-�)>��$ن,B���5l�(kEro���*�Y�� ��tlT<0�FN(�	��Z���oO45��,Q��KK���9��+8&��p�.t�IVBQȃc���#f�&�M�9:�=�?g[v�X��\Z{)�$��#Q������z���L��-���8�/o*��޼%����5�O�o�Id��Y���1m'-���ê ��v��p��U�W�o�5�K2���.�5o&�6Dt��n�N�d��C���`$�?B_OR�u~����1�����$Ըvu�I-�7��_x��\�����]ޥ�ù]������5�P1\��!��m<|�;m����VҲ��a�,/�@�RagP,o�+�����.�����>��36��|�t����r�aN��`��Ͼb*?�^=[`�%$��R�i�&Z����h��(w��-}������%��W�l>X8;{��l��"Q�/�B�]��\��i���U�Z���7��P ��M��mO�#m	��lU�?D!��ZN�n���x �"��t-�u%�=��4��9��R?c���$v8��:\��>&���{Mrd��0ʯ�!;�	�j�W9���wѦ\���^��e�\��QvL�ˏ�C\}�ulI���#t�ݍ@�m�8��ɲ����W� ���w������(�  �Q�R�(T"� ;�4t��on��鿐��^�	����35�ұ BE=	{K*��uI�~�Q��f����U�)���(�6Uѿ�t��R�tЏ�[c	��`Z& �_��,�`	�B ff[u�Ù��K��ſ0���C�ɮ��7Ŗp7�``.`P
��
~>���@�Fs|�}�W?���� a��9Z�V����<y�aȈ+Hf`�����P�E�-��[@BP���qf%�ƈ��/��/F?Ԙ����.��v)1�)kM���Ы-y8�6��l���[���7eo��vju�o�@�.�j����T�L9��A�8`z�o��|ܬ*�Z �[��Hy����x"�:3� {W��P��?����ɬ��I(�R����3H:s{��-_J��d�?@V��þ[�i��#�t*�a�����z�y2	�ȑ$UIP�7�ϝ�8��XLӶ.ap�P�b<�D�Ѹ�	tR���h�{�H�d���$�v�*(��т�D����h9eMД����5������6�Dˢ	���)���l5M;���p�ড3��e�j���"��yK�S�E+\�QW�9�U��X����S}~E���Yi�Ʀ(gڊ���w�0���KI�
?���}C�;��LP]�9#��3TycH����@�QV4��q�<C����s=_�]h��b�R��Р�C���������������gXq����ͥ��	�
	��(�R�^#*hyR�\l����,X�~ꕒ3���S��t[ԫ��E;'�g�*li_T�
�UF�W}vii��l
J���@^ۍ֐�tO&n{i\ �V�{�?ڃ`b��JX3�?Т���b�־��;�氫�a�;�Y�j���<�M��xy�}�mƀ|�O�������/�N����L�g�p�"��x�\�Z�Q�B�HZ��2�A��9unKmu��t�J�Т�c����[��n�YM����������Z�P��N��r�	�,�(Bv�)T��J��[ _~��el�̧3F�"A*H���"�Ŵ�ju�*� ��H��?rYi����J�L4"�`F�u&�KآU�&',u����,C���}����N���]h����%$�@�825�>M�9C�<<p�����W-���t�Q'�{ǎ(_��a�m��づM��S[y3c�ZUn��B$�	�"��}H��# G|UI�Ǿ�J>	�見�@e�U�����fN]�q"+j�m;���O/1L���\Ö��k3@�%�*���/�ϋ��B�!Õ#�b�.��a���N���h��\aQz&���a|���|M�qa�#QhAٮ70�E���)�����!~�� :���z6�h��⽆bV�(P��
�7�Fv��s��,��i���>�d���	O�/�F&�7 ?2��}�����xA�Q|ƪ/1"��mS�j�[�T7�P�y I�F��6�I\�lɟ�~�����6فALӬ�`o�ۄ��&
��2�[sL���s��.|��(te��v�^�������<.��@`�4���w晊Cc�T�~�^Z�Mk�_,�)��ei��/p�r��J	��Fr�p���)�?S�a�:��DM��{]��(%!����Z$|���M�-1��� I<��yO�V�����
�
Q���"�"kbu=XwY2��Z���8�u�)mT�9�IڭA�2��,��&��ʪH�2>6��C�������٥^��lͲ3�k��8�2�� ]���	·ݯ�â I+�>g���p����w��W���
�5�34�?�C�Cnc)�깶�:�����S���M_l�%]���|���������"�n�5	��O�vͣ 禓�tBJͶ��)�ۇ�:�8x7�%t*>#���:*��+� �;�Z�O{�&������iy�?���W�b�)���H��y�G~�o*�K���!�tE��|�@&�|f���Y��<�+Y�)���ӝ�1�:� ̉b��=��A.�r��B�џtB(���#�*���7�#�KG}�'�t�o�����l����6/�V�V�J3#��"N��2��A����=
M�f.����L���K;�oT��xy�EK�a��*��j�YUjpY� �D�Z[n�S	�5�D�(˾K@�]�Iyz� 51�j���7n��G�w'	Õ����zb���x�%t\�y�Rv�2��Y�?�`�+����55��4%�p;Qn���ٶ��'�����_���B��h�0�ÔEY���:9q�[؈��p�2>?OHOl������v_�_�X�"����l:Zo�I�w�_�ҍz���5˥�F���th
�q��f۪�[dM6�נⶸ�@�"R%x�n�Wr�h~�k?z�j���j�=�o�=�q���}���sU��/g�h�E�!�cQJ��ktDl4�@�|�b����5s�r����AIp��:O��h�?�s����*z_��-�u��k09��(��T���)�a�n ��z���l�]"�wT���Qƣ� ,b����t��'A��e���fҥ:�Ҋ��e/�̄��J3�ElΆ̬�G�%Y%�k>b'�,���c�y��e|31P�
�ef9��-�.ϧ���jǳ���9�=���Y� n�W�$!��Ɍ�5E�D*������fZ`3�A�S��
��HK��� Gչ���o�P6�U#�U�=a'�B��:��1S*3��	�JeJ�q_��)��R���h��p��$��~Fh�b;���|j��=����
Χ]��N��O������y�Cl�b��[5
��Ǫ-��k��)g��W��"p圎���#vy��=�ɂ�.u��\�������+�ݟE�ʔ��xS�����j�N9�M��*�ޤi�u��Yq�ю��Z���b�÷�F�ˬ�éT�H�&�A���"@j%o-���{G5+v��X��x#�\8-��v{J��L����
4��N�`�:�Cɤ�ɍ��"	�몝��:�?��U��
SxmQc�3�?Ξ>[��tF�ˠ�G<�?A�H*��U����*Iʥ�����pw�P��������*R[ '?�+g��ǣ� B(�
{J=a�&�A[k�K�d��Ń� 7<�pόEmn�Hf�Vty_Z��.o
��Ȑ����&�H_��E���q�AlR,�Ye�7T��.O,1
�T�d$�Ž�|"��P
�b�t�TN�Q~a<��f����}��JF�/��́�k�(�K4[���S��d�H�uL}�,��d���uɀi�ÏŀO��wW�f�c{q	�퓡@(��1�v;�֍5�����^F[������5z�C�w�n�T"�ђ�Y;O�w����H�x�V�P(P�߽]�%:��\�����*��Q�p��p6�\��;p�iX�7ԱtC�7cc��ǳu��{�Z�$R;�tѕ��/I�-@nԳ�\�]T��[�� ��fK���$��z���Q���z�#�����Oq�� �)��LM�2��W��2�C8O;ĥD�^U)"8��ٵ�N܅{D\QC�v4�	�i�,�{����3L,�J�`Z���;X�oD��{���2�m�����ve��*.P4��en��=��iݣq�Q�����&���� ���ȿ`�<�J}�ͣo$�1ѭt�;�-/k}�ŊP��B�k$�5꾛Q$���f����` #d���LOX�x�F����ed��M��� X���9 $�����VI�^���X/�[c}��lE����B�L���O�hn$Nu��k�����D���J�C�ق=-*s�ce��$�;���ڧ���(zݶ ˉ�e��K��G��#���'BY����Ie�_�F��)'Y}{�$XU�W����-S_ra�V�[�'��ϕ�L} �!Մ�N���6B�Ah��m~Ȼ��'t'v�[�vo�a��6��ϱR�I��m��N�na�����0CX���<�!oa�A�u2�@���1�����[�A�MV���� �		e�e+aMh	x�.�ax���48��E&�7E��qGG�� 6�ӆ�O��̀�y�Y�NQ�`����`��vSP��q$Ŏ�g���0r�1g�5��<�YN���Uϫ��L��{��,#6^��E*��C�Q��?K�	� R; �<��w����=��a9DV�'Gp������,"dP�z�Z%�P�0WգC�]m�=�����8\�����r��D���A�ώH��"��S��|%�c
ӗo��;�4��ARhBFd5�8��(�����1�m�g]-��Kv��p���G��3�`����X<��^~�n���WUV�'�lzb����>�WO��qk�f��JBM��m���0]��/rᚿ�Gv@n�8̷b��?�����u���7(
 Տ g1)F,`fNU	�:�8��i"�E�8&t]��
6[�U��S�-`�ɒ��Ђ����P��p��7���R/:�� Ə�}��%�Q��e�IeD��dY	��(��[�`U�s����*G?$X��g���Iܕpi;�x���$��b�7%�pX7���)z|�
�*�y�@�*�'�o��A�1�>�Q�@=S�96�g�@�J������e&E��?�ܟIa�(zW��wCo����8���#Q��F�Z�����{�W@4k5KW5>����~��w�Xy��!%�ɱ_I�a+ڻx,�[j�IK�}T��t���+�0���O��'ˋ>��쬺p�-DY�wa&�A�W�,��eY���P���fd��{��F���i~&���� gȡ�_�HU�&��>�PlRk����f[�T�X���%�t� ��_s<mƬ��Ӈ̌n*�@�'j�S�{�A'���C�7G�����O�a_��dUs��_LZ:`���p�]� ��/IZ�\����R��r���R(0�u(�"��ZH�e,q���n!^Я���a攀�I Q����U^�xy����;3�{����/e�!�]4P�i�o�$"毧��{Y�*$Q�����գ��J7�g\U �ܷ�A���jn3���5�������ұ4�1T��+�-KZ��,H����Ph�.����t(����M���<7\\���r?�}�v)4���A �����
�[����~���������^=�H?���w�����Y8T���T���Y��� �����8(yAű�?�v� �3pv�9�ڴ���D���D�!ɱ��'��-vQ����AQ��u����_������J�)'����<FZ9?$,��E�׺�oH������a*��1��^�d�Q1�Kk�-���p��+�&X�=���MY��K��ZfI[h�d���`�l,�]�1���R[�s��]�PL�]�q^>��;4Y%4�XA�n��?D�l��P�jO�s�C�R��v�G�z��-YÛ��L{����=�S��<�"5 ��!p����w���>B������R��v���&�؍�^�Y=���9�d���͎�%�� ��eD	m�>H�ܴ@�bx�X���al����"�i ��8ƜSY�l�1=BZpԙ���y���;Z9X�w�IKs��{@�A��}=_���⥌�%Z�#�X�J.K����N�z�g��i��\������EV9�>Ď���v���m�����4R��(W���ܗݻ����9���-���V�I ��`ܣ�>@�+@��\a�js���V1l���9�n�&��Y�,oV��'Frh��pS�ך^ܹ7�U4��4\��>���R�m.Mq`L�l�>��m����l��=��MMS&�:����|3.j�F�߀��n�_�KG�};��;��%�툼A�Ϻ�C:Ex=����?mm�R����@۶l�w�#PՆo]�lr�ގ���b9ٹh�^f�=u�n�G��H��5�����g3E��n&���0ck_��6#bZ{o�O�i��M�����m`��96.h��M��hQ'��g;�C9A��X���v썅��G��Ϯ0uc@q�I�LM�xno���<i�'�[���\'��Ex�b�N%i��Z��1�K�(�0𐜬U����0�By�U44.,��\'�D���꽛�\��E�����-wo�IBU93���R��W�Yqm�qUK��9G�>?O��X`���[&�F%%�"R�M.(�L-p�߄T:ʟٍ�U=��NhM�rx[�\P��ؽÖ����_\��1nh������ӹ�q�����	�S��-�ՙ�h8\\��6C��� L�)��++���7⤛��q���$	��'n4Ԗ΀��q���b�	���.]�v����pҵ���E�}��Հ�j�j��Ke����S� (���0@/� ��������^�r�FTζ�I�'�F"�n%���y�@:�z�-g(����\R��H͕�C��ѥ��n�E�����!�Re��4��&2�4yR�FJ��Cֹ�J��QO&��)cv@�Y���q�C^�\�/H��WR���Ž^��N�-�N�W��� ����셒�(\�x�z����	̹06�qI�<*̶Z�E'��,*H��n�y.��(�=�!���I)�,�XY�c��9�q"�ҽ66]VЏ�ܛ_^
��zB�.t�A��C�����hm�E4rM�7�l��c	�v����Lo�*_���Q��Q�`�?�U�B��&K�X'l�hZ�e}��`*De�0��=��LS�'���?�}�9�M�I�&v0�5.��	~d�uh%�복����� r����`!Ex�0�I�JQҟ.j��R���DH�>��j �@�v�#�&�f��(�H�K�8�a}��N׆QSM��C��p��	Qt����E�kCH��3V�ȅ��+]�E��� �!��X��j�?��ke�3q�a���po�R@��
Q�f�Fx!�:����k3`^4s�2�B��>��	�e�q�8D��P�k��Y�߲�����tխ����A�%Y�:$���}��֫�����?��'�e�ƾ;�)�q-h%UT�8<n%��z�1,pB
���uVi�A
��V�п'�"��IV����1��W���ԏu�	H�x�����գ�ȭM{�%�KLF���X}֬̒�,��ē��.��2��������Jva�ӈ!���:���lͳ){5$+
��s���}m���zoK��x��l���Y����Q����wA����m㽎� :8>y"Qk�q�l�J-jR����I���	n���c�x��Gz*��`��.���!�ѓ�b�4u�)Y�]��l�Ķ����G&��g$�U�	m$v�A�5��"�B͊)�x�a�K��\���&��h�����X���Һ��*3�D~~�S����'qb��E˜���x�$��@��"1g��U�>���@���_�5O=o�i>��� �OE2��)�LvC��f��I#"��\�l1�t�y�Z$do9o�.�⨊������R�
SL����5����bi�S!�y�cVH&��~�
!�g��
��Ӱ���v�a+���v�����>�����ɛXV\]Q��F���c��v�n�Yx�99�*q+��T{1��ʿ��+��@���xX5����{M)X+f8���O�2ZS�:/AO��M�O �o����Z�yOsd��	��j03�T��V�Ȥ-h��+b�B���C0�K��J��3T ��q��0��
���W�e&	��1�	��XT�!bH��.���tW�G�޷�G~�#�"H>m��C�;�7�f�I45���+���E>��oA|��wH�'����5V�λ ��7
X�O
:�M��ݪҪði'���
�O���ʳ�OL�����(�ER�>�c��Y�qʿ��"��(���f��)j;���[K.'�zy�ỰB�T���i��׼/��?��jY�@d��Hi�1?��c~��`R����7�o!�QA�l0��ׄCV�=�
�J�E�����e�ݯimF`zE��E8��O�>���L*�|mP��O�	����>��g�C�,:X�՘�U ��
(B������dX(K��B���w?��s��BP�X�p���~=��Ҝ�sv�0#�c��OZC����1���;}�.sp_��D>���Y����߇�
�ܛ͏qdrU�ʑ�n�%��a�[������{��$�
e�X(�Hf�-����A@4��#9�؎>t������ΕD���t��cƃ��iH%A%(���o�6����g�+�~>�5F�gEr�ӟ�f���me�6^�n��UX�����ܱ�@'a�2�g��I6ģ$�w4ņ�����s��D���w4�c�JT����פ�x�aK���J
�$AZ�1k�|���� �W�c�L7����t�@5�o��.�.��Ը����W���p��r5�'>6���TK�Aq�|At��2��@�)�b���!�9��_/��ê�X�QY3ge�އ�h��z���䞦�up�-�0��Ջ�P��(�� �?�/�;[��#��1�D#��9�Ӫ�r�-��_ײ�C�����Cו���1�����My(�f�P	���X�2+ڙf�Zo�Dd���}cc������_��
ŏ	g[$SP����,���\P��w�w	�/p��]�!��j�w��Cn�%�t�`��A���b.�Z����Ǝ>�b��Y\��
K��t&���W /�?l��Jw������a����D�_X!�Vw�,:������ �?OI�J��p&ÙA��9*B���C�-���a�v~"�������0��Wn�g�{u�*�ٻ'PO!T�a��e*SI<5�wᛞ1�d���# 3�:c7>��s�G�]�A�]��*�J�C��ky� R̛��;��)ĳ�͎��>��>�D=���Ʋ���N���Nb�*oYhװ��{���p���P�r���.��
�8�ҹ����Ph���)�!���܍ei�O';�R�F}�^ Z�h�ӌQ'�C���.+3�T6����ƞNv �S2�RQ��k<��o_"a���������|��]4�m����6عV��8�EH7m��o#���e�x���;��M̀82m�ݳ�N�{�h�<AC��rw�y,��Z#�f���%�(�a叞���bA���,p��C8y��cOzAH�Wz��<�z9	��R%b�6��o��Fպ9ͅ�z�1��]�M�N�Hܿ�獡-g���%rӎLgh���k��h���rP��0�&2��;Ó;HT7���G�|�M�bH���2�X1��-�[�2��C������ـf� /���5L�v�PM#>u�^(D/���ex[cy�Dia|�l�k(r� �Ĺ�B!�;�[�5�����~�l`����%L�e�ͪsCz=���L{56�+��h{>P��1��o����j6����s��%�����D�\f�.yԋ*�[G���+��H��^�}�=X�\� T��ʡ�]s$�* �0z�g�|��ܯV�]��{��t�:�V���`|--b�t����>eTA� ��E����H�I� du7S< Cwe;�O��d�0cǥ�/"����
6pg=�^��|r���T0f p���Q��x��=��$tL@�'�0d�H�������:��x(l��FLŒ��?��68���8BO=mꁋ�#�w)��G�1��G�^��Cy���I0���[��UV-:�偹6F����-���2����̃TW�=w�k�儿�˽a��J/ε���֡��[U0}7sLO�bZȗ���G[��f���Ǌ�\��r�����X�tCF��ύd��9:��yE�qr��|��R$�ߢ��j'-m:hU�Z��} o(U]�ؑ|B�\ƀ�s>��)TiP��-�k8^C�NIQ��v�	�-��
���ɱ��5<4�����:"��a���ݾZ&�\�j� �W4kU�	�k#�E�!��-.�:@�ƫ��u$ʡ)<}��k����#`�vC��*k�VYÂ�g���+ʠ�K���A��]G���ᑫS��7���NM�.<ix�KLZ�����V�����"@�%)��i����#hj�i2��b
jC�ղ���{ɫ(
zs<L���#L�n���^a^j�r��	�V�/�4�̟��F����K@he��c.���%�e7�S�(��ւS�6�,}�t�����:IlXOJ�x�iQ:?����?�ѥ�������l1�.���\g+UC�d�@ݵ�ۺP�2^o&�ʼ�T�Rx��Z
�a^��E\c�T��<"ce�El��̴F6(�d$o/M����Gݼ��^�a'5��kpY�ts�G��3�|������O!P��E�Q&U��M6��]��/"ǲ��qLkG��n�+ۭ$ܙ���
���s��RC�����nM��ef�}�r����;1�۽r�Vu:�ҿ���и��~�S�LE?�^zI�p6&�4���LS@�̝1�h�AqE3�Xt�Hҍ�[vA�#kX���j6Ф��:��d�ڌY�c2a���s��e3h]7�v��@X�m�`�ix�������V"p�;����臯�w��^�-�{Fs��P0���	���%��ivp�v��������k�:~�;��\��/���ah��7�T0���5�$u"֊�G�rE�NJ��	�QZ���/���������M��t��C��K��tI`d&E�.rl�P��q�ML�6�Dv�����!�� &P��3�H��8 !<�Qy�4��獉,��'5�|;��b$k��<ci���5Ʒ�s��3}��ҏ� /�k�d+�)���u6�v�k�Z6���Z��m�B$.U=�M$|��>M� h��x�Nb���n�(͗���z~w��<�f�p�{�G�Q��%��i���a�Q���d��p$ �;���G�4���wҴ�~��}�eE���E"��w'Wtyq�+��w��#&"DR����>���A����̯���TJ���խW?�n����&�M+._��9��I^O%�! �b��
L�~�ʿu>/�R�)x���cj�Ҋ�<���������=� _9�[j�*�0�{'�f���r���M����`���c�y�-4�*a<��9����h�$x�=	9��t�1S =V��T�'�z����Tޜ�ǘ�
`ڵzј�ń�	&Y����NI�9�v����z����[���W�sh���L�� ������ۿ��R�������)X����Y��-#yT�:��v|	3�Z���N��#5Ol<���O�iY��㵤�I-��@Ԑ<sP�GG;{)�1G���|nf��d��/z���&j�^N��;�9�&�S4B�.���w�ٛ�H؞F��s<=[Q�D�+!X+����B����,]
㶡� �E��òĲ����7��jO?��BH��&f�
.�0�\���T�7Y����,����w)rn#���]�E �d�6P��w
Lc�A���!x��#���>��(~_��ވ�����=hVDeȎ��XM�O>q����F�F�t1�y|l���|~Y�3k��1A�C��mS-@��d����t/ʽ���y��lp�	+I���u�R}��o)����W蕢�Z\�|o�z`��(
�j�E4O�a]���ʆ��2�c���F}߯�-G��� u9f����@�B<,�EԎ�
\����o��؈��I7c@�IIl�<�����I�b:�����]�d�%��RN�%^Z]�O�{F`-�C���r�NEZ��M�B��T\�s%�e������Мe���A.j3�����:�D��=y%�`\[l-�ZM8J	�]�ȰP���0��P
�D_,8l&s��9����j�*�X�y��v��ڃ� �R���"(��+$j��e�vۚj}I1���C�ʵ�F;p�	 ��]E�3^����69t~{���m�z�MX}�J��'��x�j�$���%ګ�l[H�z�fQ�g7�h��n �6w��tʷ7cu!Q34�'��z����)�F߻w��״�/�Q��E%�[�}�ew a0�T�u��Հ���]��`����<��6�0y��g������}�Ѻp^|�FJ�ꮸ����?���O�g[g���y�O����3 ��(%�qj�E����=I���ڟخ��Z y�y!ϗ�B3r0�������%޻	��$캜�<!Ӌw'��Kg�,n��~)�P��ω,��u��|�YJ��S:l-�:�x~W�'5�C kN�4	��oy���<��][�����L'Z4�|�8A�&^��?���,ES�4�\���B�#O_��	J�����K����rTR�x>�K�Bt,����U|ʾM����u�S�H��"*V\;��T���S�� �v�Se+:Gΰ(X����9m�G���0RZ����Ϩ$&���N�
�j�fq(L: 4 �m���f
f5F;F���zcK���#��8v8R�A__��[.W�{?���<��] �.�Ѝ�I���<���'a�n��{�b��%��5�f��l�5o?�In�A�`/�X~]�5dP��P��=�<	S�2���p,�Ev�&�%`/\�@a��w�c�tS4/A"U���z�?P��T������RLY�<w�ݮw���ic8��z~�T Dl���ڲM9�����#�^�'2�޾��z�M�<�U~[�0%���!~6���,8�GD�,x��"l������.�g#��-o�1�+Ӟ�8|hssX&��1�5�V����}�'�{����>P��� |�G}�7v�l(����d���P!
�U�+�2�۸K �|z:Qݸ�����}_''*[�\���k|��IR�t�[M�f�s*��̇&:�Q��0�|W9�pC�Tbk��[(?�����1^� �����;f.>�Z�������W3���Q:ZD�z�7�E
����� ߣ5�10�0�R8&|rB2����s~��!w����D#��[�6�O�!0D�F����ĥ�a�=��Q�4�S�@
�}�,�r�-��D�"%�bG%3�D\gj$(J����t�t�]R>�r]}K98мs��DI�>*��7b��%�����p�#LIBe��9��D��]q�ɥ�����
i��tu!R͖}{ Ti�gU%"R۞�<|D��?�@7-�W�L��9v�F����Jv���"g�ȕąLl��w���L=	w��A�(�)4k/(���M�X�6�kJ&���,UpF*T41r�XƫK�����i��<�{�K��/���Mi����`T^t`Hk�#f���l+%���Ձ�h��-�ny���ok�t�f�<�O-叟�T����#�h s'��Ն�o`�![I����g��N�}f*=��<ZN�{Ɏ�}��X���a�
2ԉ�@*����!�ݦ�@Hx�p�G������6@>Ng6������˚��>���1C8qVw�N�-�,Qꪄ��D��*|��3=��e,8bW�M�\O������Ĺ�g��N���Yl��vb&;J:�P���.��T�_G%}p�-�.�&)��e��I�Ź�ߏ���i[z��#��:>�t{��M�B�d��5�h�3����<�Ӓ�b�\S/����� � iq�jcR-P��"�8�P���F�Go�+�<�c�<�_N���V\��m��fZJ��M�'�Z^L��p��u}�qރ�T����Vk����������w'aY�W���D��H�i�ߐ��I%��+��X��;J��i^0���O/���,���|����j8��m��|�U~a��O�FBDp��'q���W���	T�l��Z����~5���)Z�94㳴��w��{.t޺�q�f�3�x�����4��XP�&�`�����]��sowű����u�?���ND�M��P2����?����w�	;� [�/y�l,a�f�"KgSk2+_xkQ[IUX5�Q$Tv^x&+�k�X<+X�&�^w9҄�:ș?y������8�K�܊G�dF4o��phf{��H�E��2�>���x�� %��V�E����o"�R��Ɣ��2V֡���I�dH&��3����M���u���F�/Sx���fj������o_�n݊�OA��}#��7s�Y�d��5��`wV�3Z6���F�V:l�@��{_X\#��#�/��8�_��j=<�PH�pp��L���_L���-�ס)�sBB��!2f�W��N�ڟ^��ғ��^^ex����2)R�b'��x��?Vx"]� �A����58$��C�{�t�k/ wD	I>�u��0ɑ��Sf�����8��b�鸘ʯ��*=�����fZ~p�q)�X@�3�p�HH<Y�k(t����+4�2"��a��/'NE�}�j����j�e�T��͸;p�Z�lYV�-@�T��zV��qJi\��]@eR���'�գa��&���'�$�B��ī��u��kG����!HC�����[_nE��V�t��Е�њ=�ґ;��[�yq�����Y�9+åt"��"zͪ���8z
{i���q"�n�8|``��`�V��L����K:���m� x��p�j��Y�*i�q�fYIXUPJQƧݲ� ��Y��mn��i�Ǥ>�\�$"V��H�%������X%���WJt[ͪE]�P��Ѹ��-f�0)�V�x�	�����f;��#H'6�ge�W�ԩ����c�!�$�����\ōC
� ���.\ak��(��eR7�O�!�5^�(�"Z���SaO����O�V���Ґ䨩�mGjY3��ݸ���ٲ�8�Q׾@t<���]��h0��%�!������"�e��l��=�z��V2S��S}���#���i��O�5����4	\���,Ҷ���&\����qNՅ��(C�Ƿ��p�w<V'���˚{|{By�v�<��aw��;����4�O~�/�۫f�6yM�Ѣ���ih0Tc�
E���?�!���2t��l#lt���-����~iIp?���7�D׋P�3�۲.@#|
=�1ѸfI�@�� ���E�2��v�Ɯ��_ȝ��X� ;Ź����X�7:.����iD����`�1š�(
 ���K�NK[�����[���|�Q���T�L�-��n-ω�ud�>�W��]���[���Z��E��٪���ލ�SY��6�?{�=r����x�+Q��O[U��6��`"?Vj(	���>(�H֩\�����vmM|������`>	�-����e�������uH/60%��T�Z�Կ>z�M�������wS X��ci��oW��G�jY$�,�)�|%���b-���^�&�(ߖ:�`�fb����o�����dZ�E�ן~��7�}kt��U������:�Z�u���.�1�	��G����a��T�Z%})EJ��*�Ek/��,��G-o�e��1)�bMX�^AEhI~�q�O�M��#�����af������Wt�"��=��I�5��7�oF�L�z���Dc�*���3����p�N�BB����e��2w�,��E\���n��&}h���Tz5H :�t�/�A��r%.�2/���X���6^�5XSTp@�;��� w��J˓_ՙ9�Ν��?�ҧ��m��$G����|#�N �N"����)�3XHy�����z��m#!n�wlc$�VBGJ�/��e������Iz~��in�Kx��.�\�ܨ��N�L���v���h�}����qVcs��>�!/��|��Bl��
hh/q��f��QuK��@/�5��qT$��>�)Ū ;�cM�T��҅A�X��Jky�*G��~_�K�L��U~�c\�ΉP�P7�8���W�:G�L1zu(��F�nF(%�H'���&A� ~��Pb���Oa�吹��:����nO:Oy�$+���v?�pב9��f���3��������_���?�r���{��y��
R/��}���31��~R��LKr�ބ0T�k�7��K�K��Ξ����p���
J�6�\�!Z2m��o�$Z�VԴ�v�	�J�,�>��ɲ�S`9t��!��1Mט�sF�x[��sي����� ]@����c���
��r��]N2.�$?�(JdB����a=�$WDsH���i�jZ�ϐ�D��[�3��{ș
���ϲŹ�̞�H�?3�P�����;Yt�{�mF�p-v&���+���D,3�K�i0����Î!��t��;ag�Q_	3l�8S+��!��x�"�����_F�6j\~�|�v,,�-�����Ш�X�M�$~T���-��_͏��׫�m���)�:)����
� ���O�j�zu,��s0M���21�r|�:��*Xy�!����u�d���6�L��fHE_#���W��G�-�?7�	��fh��M'�$�������+`]fm_(�c7y\���?�e����o���_����8Z_/"n����{���z��lv��%�V%H�����2=aM�"c�c}
&U��pt4��:���@��$#2l�l��U1s9d4�Q(�e:�|8��/:��3�?�!Wfq�ŞQ��Z��x&,�4@�#�pa)�?��^���X��� �sC.���i`�>^ �B8v�l&�VȞL�#�TG�7��Z���I��!B�U|J��B��4ȁ��.��J"����v�SVeE�K�����=W���;����r�5���m���Ќ3�p,Ye�cj�F@k�� �6^��:>k���1(d�E�o���������ks&�^O&bD��%��h���>=i8IX�~���K�;�%�X�a�{�щ��`ΐ��r��@�޹h��v甲�P)��A�z����<Y_JO���4>��2�℥�@q�)o����$�zz�%Q���HU�������Ǆ��(�E�-��/Ϯ�">��J,�u�藕�zQ��6b�ȹ�yJs�$r/�����)1���=���+o���{h�o}T����ac�[��O\�V�>��]�Mx�9��A1>i�����.�iB����t�h?<g?vTőf�j�0��־����$ '��ء#�����4e��_��՝�L޳��d���"<[f�)#��l_��pK�e��7��)��+�=f��W�UD�l�̵�>�A��Q��eWhI�Yv���?���G�Kc��������Ώ�������ZB�@[L�wiDO8��.�l�1`�msF9�~v�.4�X��Gᰣ+�C�Зy֬<��:S.��6@���1C��ɒ.��cep� �s:z��Z��2]����\���o>��)?�uk4I[��p�B �a�����Ayu���c*�������6�� ۲�Dg��\�
 ���CW�.B�X��&~��o�-9�߻xA
���=5�KWʶ�@���������4~fr�
D�M�J�����f���W~!�NGԦ}7�m��`�L��� !RL4
!u�]-2?�1���Ԩ�x��C;Z �?a�t>��P�+R�,f(�����Ck
>���QAo78�[p�����?��â)���iz�Z7Ǟ9�m�0���F� ���O��`M(��Rv��U�C����S�ٺ��C=`��[4�5m�ϥ��̎�O���h�� !y��1������A-�ױG��_�T����nZ�0:Kd��ߙ{)y�͉6��	,��{�q��l����O\�-��H��em�ϙ�&KK+~(;�x^���=}o`�X���U&[8�I,{Ë%Z�D���rlfw�[.ܳ���ɨ�u�޷��N�K3�}AK�&-�CӈV"���M���g:��ٳg���D�<�f��i�b�h�p�p/���N�}�D�䠥Ⰵ��Lq��`_C��Q��1�I:�e��/�������|�J��͘])�4�Ux�M��
���x�m��$��˨ݬ@ T9Q� ��G�#Zhs��>Ρ�+ ���Ҙ
D�*�,�ZR��v,��G���F�q�0c�}���>߆% >:�s��7���a-�}��H���|ć���!�������:��9��@q־�'�<+�)p�=\|��fA�x���2wD�T�G���FM�`��N��$����6�� ޭW��HW@�Fbo�̂Q��a�Z�Z�
(��O��%
yj����S�U񆲔F�8��ͳHŶ:�+��.Ƒi_������ś�2��n�c���p4�^>Gg��I�D��Po ��p|�@8iϹ@:e�<u�Ɓெ�F��a�,�U.�8.��m���\�U��v��y��m��yj �C�(��mf�'�rt�P]��Π	.(1\b��Pק�O���>�\��6���_���v=�Og�f?@J*o�}C���aS*j��<�<�-�����n�y��/���3I�2��^�)�Y�S��V�(�o��$\�K�hP�lX��y]�J��|&�l'�ʹaA�v�uц�@�kE�Vh����i����!E�^Jmq�I��l������XT�ApK��݉#ʻd�}ɜs!rgG�vA[ݐz��� �%"��b��j�݊�T�ɯ��v��S/��z/����e�j8H���l����ה���ya�m��weji��:%W��1i���AY�N��W,�O7���������8�Is
��[f��"d�r�`��q��x�;*�6��c�K�f�k2�\�����3_̙�30�Ěm�u݉���Q{F��q�[mJ�I�l�2��] ��)}��^�6��l���r��2K1� ����gݤ��o؊�s�(O�GjP/�@S�C���ZZ���R��%��r��F�>=�	rՁ@=m���|I����YוK��<
Ơ�W0���E�#?IB�#�`��3�Ɵ�����E�:���kΫ�����Z�r��hY�zO�x�rq��k�m�Lv'\$͎&��^i���c=�B����a=���eHO�֗{d5����m0�[9��9�S#��.n��g���E�(HM�#=�O�R���襞ش��-F��W��� �)����(ׯ���#���Λ,�_0%t~">���꺪G��E<��H��}��,
��B4�L�
�qT�<,���|�j>�Z_�2q~�!T�̣֣J
~G����Y���J�z��~�n>��
�VP>X���@K�4��B��:a�b��/�\���Ð����>�p�`����z-�d^�zY��Dݘl��`حO�!�F�%�ߚ" %�)"UO����r6ec��:/77��}�X��J�ܨ:&��k �õg�`RS�Z�$"0��:(%�s3�7p8�,�p('/���b��4Z��|o�bj��d�����,BM�]�;�e[8�b��{tq�d���Q��?��[�5��G,�0 �gac�������A�c�i�V ���ڈk�YU���/�dW����x�C��&���@K�� D��gV�[��t5�x�ca�;V��bo��Wz��S*� ��x��=����� ʗ1�Y )��n+"���**�w��ć�w؇���X�:�h�D��tp��q]t��-�ӊ]�N�l��dL�8�p���@���61�d��t�)��΢��'�z���O�K�lv��B�O�����ՀHw(1�HKBέjƤ�ㄵdY$&��o��n%R��Eiu�1�-�/��|�\���p�,� ����"�_b�f���Hd>�nn�����S5m�󤲸�k)�e� >�����z��G�L�e�q������*�&
�6�I�h(��l�̛�=�����4�J�;2���= �!`Vuf�UcX7i+r�.�r�6�3{<�ب��{�f��Q���vxU�@j\���ԕ�g ��Uq؉��b��&�D����������Y����Q/�V�|�F�g�A�+��r|�ek&�e"�@�w��D�K�A�)F��t����W���i� \�݆]<����#�i� %�vy�rƎ��_ܪf0w���D"|��H��C䔏j��� T�F�k�\5�����*�A8�|�{H6ND�ׄ��&������sgj��,�ɶ�}�Yq�YC)��if�@�c�@�c-D�x��+9�
�0:7l�;#��Jr���i:���zc:#�5�+��4ߜTqT����7�x~��V���x��b,"W~'k�dxJ�2�9�2uAr�"���{����=��F���ՙ97yHT��X� �	��.����/,�h�ō��H�8{FLa�&�3����Lх��wZc��(R{�±U��T���������s2,��C�s F���r�3����8~��sY���y��=�DA�����j-��F� �9k/G�2�~��;�B���IhO�$�׎���nD��n����q�{pri����u�u
��Ҝ�ŝ�yNO��R�Pkˬ��@������Rߝu��وF����e�'�^�/�A�I���u�D�.�E��j��!��C6�6#��'�
{ t,d��^�14���֚����w�(�lLd}�B�,<�!���ɃH��B��;0��;.s�G�;E�?�%A���;嬰mU�I��4�Ų?�~^UjkH���Fn�3�?�a�SoI���y,�A��>���ג֨�a]#"6V���6��&	J)$Ǌ�G��Ѿ�6Q�J��-&Xq�߉A,h�������d����~u�vO�u�-M3�7V�b��ډ~�@�?��-��H�u���W�л�R��N�?�M"�#Y�C!#��t��I7�����oLkg�w5kj&Z��7ffNڮ��[�[+�G�X7�y�Ȧc���]�`ƷGuѰ�j2P�݊�׾��d0߃f!�h"<�(2���t�Kʐ\
��p�u��PEP\��z%ZԷ�gz��w�<��Ô�.@�w��ג�-��٥X�_I��zղI�A�y&vSb|���`�<�����0��Ih:vn[4�'*ƃ�\���sQ���m�S����]4��*J�t�MO���;J�֯C"F�X���i� ��Lb��tUiC�j �G�e]5�䟁�[O� �~(��1˞$������(}��s���Y�8C,s�y�9�k��V8^��bh�r'P��Vۭ* �u�p'CP"D�;�^0�w���Ri_d	=&Uٕ���su�]��K!�/뮃�CG�!h+��lͦ��20�Y����h�3T�3͞@���g�=Q�4އ}k��mk�0��c��]و����*#MS��/^d���ɹI�?�Tn,�[Y�R �(Dh����eZ�,.��q{�k	���F�� ������ Ar�$P�z}kӥ���
�Q0}E9�����A&��搫���C*��n:��Z N�x�MTkX���y���1�)Xqn>(����z�FzA�`�ʕ��:g������-��z�K*���vB��I5 sJ�l�aÚ{��Ջ��+ ����U�Ђ�ҙ�.�Y����6�U`f.�B8~�.����	T���_�3`��	_t|"�،���t�n"�ML�)��Q�f�;�o��Lm,2�R��Չ��nVZ(R�p�{]�^�Wmk�F
��z�����' ��xY|�&8�\8gZ�>�����n�F69��$���ߞ,W�s��c�T]�����	A4WT��D��7�P��D^Pp�K�)0�V��Ra�v:��Ԁr�0�Hܨ��8�IC����ab�J���3����;��w+���8W8>����Z)뙄*���YT!u��9#x[R?��8'kԴ�C���:@bT'4*3�I�jf��;�vxq��Q|��uF�U`�s�DJl��k�/�%��%�p��d5+�V3/p�3�{6�԰|^s\��f@VW'�p�w�����L@��u2�irp*��hQ�Ii����a��UkxN���)�R����*i{S�tQ�9�������� �0��IϞ2�ɦ|JWq��pqwJ�ñ��8��oY�7v�z /u�u�y�!�D�՟�i��s����iZ��|.U�D�� �GCGrx�����dy��L\,�
;i�c���&�nDT�[�,��璾���{o�!1�AC���Q`��R�+O�#��fm���m�P�T�1�i�� �HƠ�u"��E'ǧ[���u!O~.C}�T�]���4CSԭzYD5^w�}�D�}��t���
�M�A�B|�jmN��z�&ؿ'���Ti�]\,�9@2��0-�]�s%O\��9K�k��Uk�%Xk�B�Y�A�-�m·^ُ� �!�z(+n@���B�r&_�y�"U��5�,.q����ΰ3�L���0	�ʧ���(�w6ڷ>�e�G��y�Ln�J�Tb��'wK:W�3=E;�<k��K�r�e����J`R-�p��V�%X���`�!+�������q����ԭ��b���Z���"���Ժ���-;Ɣc[l�m|�t�\W��r�My't&�6I�4���Ug������/8��
^_�����0������T�i�S��]}���X,1FU�Fep�j�~��S���D���7i�Iej��q������J0*��<h0��4����.�f��\���f��RW�q�9��CrZ2ɶe+��t�%��ȯ,��TߤkU�+�M�1?�����_�YLXE��b�=��.؛�p	ͻ���ܿp��ϼ�`􌿟x�����ޑJf�)�P�z��KQ-�	4�R�0�C�:[�����<�v������@Bi���1֤qSyH�4p�1���k��e4�! i�=�2l��c6k���z�J�9U�4(ૼ	����)��d�ˮ�҉j�.�j��:�P��pe-���	���Q�q^�Q��$�i��F�[�.Dw�JF����%��d�ys�j�hn�����ƄX!V��aX�LibL��N�Rr�F���v�$�p�'�\BM�� "q�Q/P����zn�2�"+Թj��*���l���W$���'�go1�(�km3�����ٲ,�H��wp��U�J��f\%C?e0w�����
j��"n�N�ջ��1�W��u�i�i��w7�,��+�x��2�[�����<�948��o;�� �cmK��Z� P��Ũz�N����9%apJʒ������(���К��^��L�f�2΍Q�"uC�|�
��93���+�\�g���+%h�qs0\�},+��ٻ���{��{	Z�Q�(�X�?8E��5�{���/ؼ��2�G�|~� 3U�U���?��XU�����G�/�M�w8�HF�"��1*r`)j_�Z%�#s@�L��6�x��n�.Ӻq�a��餳�����W���W��ܔ���z���-Q� ��1�^�F7Q����F=ǸQ(����g��0]ks7��M��,<q2�l,�u���$��8�*֏�?�oc'�B6�������_9x��T��޷�N~�hXȨ�10E	�ػܻ��i��V�ME�a��2�+��F�]�cms����9~�F���E`�t������z���p�����ꥷX��,�|6�Z���K�\�I��,&����o쌟���g���W?r��1��n˧��SqL5�'��f�١�,���֝�����B�����,rV>g��ω|C0ӸT(�Jk(�L��"�"�	I[R���ΘDf�o��6���@l�B�L������r�j�v¬/6 ����=�< a�/�[����6O��Ή:�ݸ���G6L̟R�`HB@�5��ܦ��சx�r|f�XT�5���Vc{V�UFsL�
���6����ǌ �L|��� �TI� ��I��p]<��@�)�c��{j.R�;��k�>
8��?�M�>�w��z0^�T؟+I�Ta��c�B /�6���� �hIӯ2j�u� q`ͯZ���Lz�;g�@�~2OZ����
cę2#7�j�]|��R��ш}Y-c����R]?���L�1ġ�n(�*�b��P�9ħ/I[�h��^��N$�4[���4ܘ���D?x�����-!��BW&|��	I�9�e�о�x�f�8e��Bb�����ɴ����8=��0��.�L*X$�!���ل���v�����o���U��貏������c��GkOv��d�n��NnfPyM�3R�< g�l@}e1�2O�, xCDf��I�X$8_#��� 8b��M&�F�$p6re��{�hO�s�Pʃ�!�n�匀�u��mA���L,&=!�*̗�{Y����c/����
�N��2{J�i>��(�N
��~Dk��b��ďE���]0? Mf3A�Q0D"�+^9�D�t�1�����|�Ͻ>ac�R�
X���L�'}��}J���A9���z����'��%�v��Z�g;�]P���#����t�>AW�]k	U��Q_+(9}V�Tb|�ڙ��f��h��@��e��������BK6�\ſ\���&e7�'�_����ֿ�
ځG�@_��M� ã;�ß1�,?�C/��!�H�h�h��D�P���s'B"�5��K��7���9Iu�M�_A'b�h����p*�ӷA���Mf��������V%��B��m vJW��t�$�S?�A�.����=�Lf�a)�s^<��ӤXv���R��#cq�?��u\0փ�'[&_<�:6Q9<�6��.����b�F�^�?n� ��}�-�4�W�M��G0�݇6VB'?R�Ėԩ�,�8%5c�������u��L��b�6%�MXE�[��p6�La,��X�9���(�'>jH"�R	���p��i��m�\tpN)ZI�q� �����lf7�'���p�K�-��a\l�k������r�	�/�J���H���N+-����+l3옻k�<,�2���9�;Q]��`���82���I�B#p?ݡf�yp�Vs��mdG{��G�J�F�I76����r"�u$��V���Q`T�$��	.�5�	�S,��m������U��L�"�gkICMd�}	���׹��ɋ�+MR"�7����;K[�s�A]ܐχ��gy�~�q6����vw,��j�������S� �bK̛�j�*�քn>�32�X�'�`;G��T��](#L��ޙ�GR&������6���u�Җ�I�� �yԆv�#O<��;t����K��o�HAk(��>zU�����l�-
�T���:o��<�LƐG���/W��u=Գ�Tǥԭ����v�Cw�M�9�VS�YrF���A�f�e�ך����Y�VsO��	�>;Ë� ���;42�Eީ�z�Q�-��Y0��.��6���k�S�����餟�R��:�'%����>�Q/J(�?I�¥�#����o����E)���,�@
�rH��1� ��a���bwQ��R+��5���҃�H�$*�崾��P�k�3Hίc��w ݫȩ%�m�H�c�3W��̣���[H��)FG�S'�y���=*�z�0��{���G��	��2���Ą��w�`�V��N�����L&'t>�a@P�|Үb�Ɍ�F�ȭ�+aZ��4C+��%����basG�l�I��ռ�=��} �q��_��
c`9�?O~]�L������M�	�#�Ġ*p�x9��3if�p��z�fMNk[2U)U�.�`y�24z89�w�,�mѝox�S���<P�׺���WR����o#2�`��V���'�9�cu{ރ[^�>�9�V�Ry������bjb�r9i��8�����W��9�c�C"�REs.�Wp�e��܍TX��	m�h 9�I�m"�ɰK��a�\�y�0�.�F�[�O�4�ay`��b��`aC �:;]�(m������«@�pPv.l�N��Y����ԝ�,�N�����t������+��${�\��Ɣ��ї	���"䝱'�ѷ���^��/��3�j��1��Rig �	22��;,<F�A�"���ȅ�f��cp�!��4��	�v��s��Q�Ur��q��Ѱ��іہ���*o�U[=i�	�Ig�t�������J����ۦg��v�^����_�K	�5�&�ҿ&����E�s׈.֗4�З�Ea�x�ʦ�gX_]�бJz����em�AL���H� �R�C
�S������_�A�ʫ�$,�`ӂ*���Z��p�P'Ie��Nb�̀m�*2��& �3n�%��9�^�E�t�] ��ɱ�]l��䟦z�³�	�6)�HY���o׵>��T|������χ�-Z5�����1��m�結p�x��=bӧ(��ݖ �y�/}=+�k�W�KD�'���"��zO}Q���-\C��͟���P������pB0K�Y~?��nēg{9�mK�
ɬ��]�(fP���@�������qOt�u�� l��k	"y�W�"Q�'�u�����3���c�P�`�ځ����!}7j��۩&/ƥ4aoF��ћ�CD��h�CM}��J4�6.���&H#q=�z6ʕ�װ�Nk�M��2��6I�S�4VpUxH�Z���4R�w�⓴�i�9��w `W� "[X���
�[z����;2}��R�Z���OAk#v��Ye����ts����o�YIʽ� �W�c=%,|��#ʒ9M�7���LlP���Z��y�	�w��O5����y�챤4�@�E�9������5l2Ц�PM>l@bb`L����ǧ��"ႁI��pū���+�5d�b�@0�����p5�s/I15�.��,�\�78i����
�Ir����FX��VW}v���n�y���R
������ɓ�#f����H?���&ܢ�X����o!1��g�=�s��,&�_)���!�y�k`}. �Y�gG&�2ϊ����:�ы�7�x��-�C�qU#�� |I�^����5>�̞�잋�2r��:�&����<��t�N{v��Z�G�,M�V=d��$6��[��4���t���[5wC��,��u�4j���1��9/*k��2��*9VC͈QC���h׼$B��Q;�>'t���hp>��1�D@4 G\�'Z�G_f9�q:���ni�&��N�"����rM�ӂ�K7u�H�W$���L��P�g�vYp�J}��:��� Ey#( @Hop{�)Mk�6�ΩE3#���;[ �?��ә����ja]���D�O|qes+���p�h�x��h�����)!K�ć+���_mr�L��Ȑ�F���u�BmR���||��-��o�2��:}�r�����n}�j:{��"��"A7�.�[��+A�T"~�s��d1h��^% Fai��f.F1���d�����%V�P��%s�fY�W����[6u�(❀쑄0��S��2f��>���ߕUV{zy��M��躱����纴���v�%_�S�(i"��g�w��a(|�� /q�K�P�!K��]�4[D���Є�}c8��0����=��y�>h�Pf�&5���'Ma��mi���JΒ����޶�e6�G*����@7�-�����������B�SR���ͮ%��]2��/��l2+��dH�s� O�`0�ur���V���Lp*Eda)T������9>��ˉf�K!�~���I�㒔	��z.���0����q�	(4 $���*�sSѓoA�S�G:�<������ ��Yo��nˁ{�t��i�NU � �/����]<�t�z(w�
�%����I }vM���\��^�,��IC����!:�����I��OF�m��N�W��"�������:nA����~H��[���}w�[����Ҷ�
�����Aca���ӣq��{��r���:��@n��([�ڮ���S���f;{�p�P����Ȕq/R���A#o�ұS�~es�=Ĵ8�c���Y �#S��e�)J��R���x�Ŗ���*�@��q�v�Z�:ZY�N]�(����|²���ӄW�c6�
B� ���<H<�<�����4e:}�L~N�ˊ'3U���*_����K�h0'@���~�(�D����hbtv~�䀌���.�b�Pf��E��*Q���~�~e{x��f'ךi�����+L�E�A]���P������dCz4�!�6��6�a.�@AU�l�(�	�ԑ���/�'*˃�cq�j�]�?����J�iv��1Gg6��T͖����_��*dM�������4{9��rHM��u�#%�"�iN;�ȣ ��C@�!Q��h/k���c���r���%]� ��q�q�~�P�v��ׄC"9ٱ0���Î��֌��棸�p�E����m���k L����*:NH��]o�d��yq4�;�Jf�	�+�3��[dO  ���8S�l�Ua隩�EuD`ƫ^^dp�L�����o���u��Z8�0c��I����J��MKzq�a��y9���T0 t=-�cQ�2_m�C[D�Ģ�4K�ӒX~�&t��{y&Z��?@�V>�+]�y�&U5�3yuX�,ى��O�]����;��g�,R|�0�jA:�&�Ռ�덱��Jޢ�G]�G���k��ׁ�Nm���j�j�l��)��f��u?�DC;�A�E�r'9���ÆI5�pl,���頭����s���1)���S�ӷ 7I���A*�����ȑP���Q�؈�v��ʁ��)�]R�����"G��i����
b����.܋��9�w`f�V��N��;	v���Dgz�������3���G��D(R�P�
y�ᜬ���}1n�ɋ����pw��u�	8%@�$��T�H�e��j����S諨�܏D����֌u���z,���H�ݸڑ�,ƅ��X`@g�������R�;��Y��
;-�+m�h��I����#g,�;xi������0��_U�v��\cAX��|G�һ�,��������y�0��誒�s/���7h+)��?]��+�x��n�A.d�ld�C��KQ���g���d�Q�t�WM3�r���[2q����rޛH��x� (b�.�p^h����a�55�^{�7�>ڔ�Ҏj'��c��>i-9�s��כЧ�/gO��x�&��J�3D�h0)�=�a�O�v�η�:좥iƕ���nv
=�'/�v�X�TH+��������,���	�����C�A�66F�R(  �Uk��x�ܿ5	��h3C�;ɕ�O�ͧ��{������rsδ�/V#l������=�ASk������h=�2#at�/u܆FF5�kU�[Ǿ����$�X��R1���� (z;���/�-S)�P�^ل����E��8�ʇUk��8�}
�m�S��{�z�a'%]��|.۳3D�xv}^�$�$���J���Ѝ�>���m��r�|��~`s��~�Ҵ�+%>�GE�P�n�t
V�_SJr�TT!P�����ş
��	��-�y�K#r�g�:%/wm}6����D� ��}#���)j�EȔ��\U=B
x_�ƴH�'���}GJ{�@oչ���e%��鮡DW�'jRS�%�{���V�x�4��׀Ld6���gж���y��LZ��(�����ʬ<[��%B�a�3��IXR:��^H��Mΐ�;l).F�lE�x9�X�3n�R2-�@�����l%��Ԑ~IP��J&]��۠��ǎ�%
j���g��%8Y��"+c�G��8�^~F��? ׵*;k���ٍ�A@A�N�լ�$�@��p�QO9���d(8ŷ���Y�*����7���=|y��|;l.���]Y��`������f��
]R���3c�P�$�+�>�+��od�I�ٙ	��a���p���B���IN�]?!��n�f��q�9)�����{d��[�V+�AՔ��Asz����cOƌ�DPK�q?����#�i��'�D:�颵E�o��܎�SD,��T,�Cd���:�kҖU@Ç�ۣT	s�d˷B�z�n
�����<�$��f[�g���m�h&�d�(�U�%��|��X����b����
��+���I�{�m�j�"5+��!K���čN��T/+��둞��oH�W�S�� /߅�$SplM%2� `MJvt*�=��!��OлB�i���
��u/�ɡ\�����*M>�LY�����dS��{�`M�Y<�ͭ�`����^��U��h4�3X(���V�no�%����e�Jr�����ۓpH��ı��!,�IM���ϑ��
��X��#P�e3m�XI�RF�u6�Y�/��l�t\G�8�zģ��jӰb��CQ&O�+vEH���.���)�>Gwr_���W���PW��4O�h���'�~>�<k��EO�CAk��-H����2Y�RBN{��$�t�ߺ�[ac�|�TB�u.E`��v�@+R�M}e��A(�EU���:�_5w/f�ð�pk��@�?N�$�)�^B�J�.��ҁ��(��&��[�Pq���AN�g�W�a/!/&�{�/�Q^}��ߑ�}������]4��
@�w���S��,�`���XF�af���!;]��$�eq��3呵*J�f	Pv��\��y��.M57��`B��_"�=��Y�3��h�)ݫWJ��`���Q�R�.�՘̟p4<΀C"�� &QK�������N���ӢY�2��e���� ��X~P�\����@Ψk�[�����Ì=��^�-��y� �0���.HQ=J�E���rM�erQ�ϫ�N�u�Zv��m���q=.&�ӫ�|.�K�U�'	~�8P2y�Zq���&���:w�+ʞޟփ"S�\L���M��?�bA)�ix �
�w{]�]�����~���>�����o�BJV�a��!9*i�I����T�s�3U(�D��ކi�!�_<(R�o55+n,�n9M.ϋ�XwG��ʓm�1�Y1�o�Ӷ�SEz�.�����م�{4��G�#i7\�w4r�������hA���y����d�Jg�N[�To
��׼���Y;�8�h�~i��9�/�f=�N+>�E�����J'�`�j�e`[������}TZ$����l��0�6���t@��K�Q��Y��K`����N,��#�b����u����L��� �G;�}��s7sֵc�&|�P�+#��Ytlj:Ls���ٱJbg0�MJ�*�/	���ظ1?_z:l�@�����|�ȱ�e��<U�D�Ư*��CE�|֌@U�#��[��%4�⤲��ض샴��H���q{e��(;���([����<��fȕ��W������/Wui�8pY�!bH��<9sm^FX^i�o}=��,;�3,#�E��X�6C�4\"����^ÑG���ƒ��[1~aL8i�D.��]�u������
�	�瑳e�!�f����:���&B�33m]��"3��N~\L�GF��t����5�Z7�(��f���%Q���
X^U��@����$
�����:�znL�Lo�=����Ys��^t:��#��+^���8�җ6�1�b�f���DL��ѿ�ox�*���&w<)����v���L}KU�] 3�@���1�g3 �P�7�����Ϩ���.:��f� 8i�	�&	%ˑ�E�_G� ���Т�d��+r�P��)�d"�w���2��DAXyR=,ɑ�B/�f8E%`	�	'W�Msz d�u�+�p��3O�"k]�?���/��0r6�L�u�F�V�E�6U�3�#�T��:KR��a3��u4LEfH��lkhc�; �T/ʓ���e�/�vg��|�]*��0�	�
����wU�z"S6�[/"��.��)�s]D�OB1��ܣ�[��N^MD#�;����ǐ�����/��N��¾{? ��=e�n��X��0'V���=�z���m5�J�'S3������3$0��F�S��Q��$����A4����M���@=��T:��Mur%t&i	��ɕ�-�w�8�S3n���OW.z�(�w摓�q��9�ըf��SV�N5(q��c4��Ꮯ��S-%r8ٴ�A�2>c5S�J�Yw��@�?G�,JK&�<Y{��R"fi��������pOn�@	��tҀ2�ۍN�:7Z���J���T5���B��LK�0z)~
!�r��(�ޢG�J���
�E΁�[�l���'.B18�Q��ȉ쬺	�_<�ʀo:s��5�'D|��D#��Q @���R�^�f_��Pu([����+�K`)���w_�2��[�����0����v}����+`g��BYݲgN<�t��^J&s����3F��3�AuL�[/J���?X���c�������$���ݧ�T{�Z��a��rc)ⱕ�����wH���� ��tc��"=w�_8H
X;�HY��i��jK���Ojг�ݨsSySm��K���Y����O-T՞=�5k���>y���@8<,K���r��V~8�5]��W��
�wB+�@l������BD}���Kf�@|��b3RW�،;�V���z\⍞�ܑ�7��F��������*n>9ᔭx��)=:���i�I�/}\�h�V8K����:A�E����ţ
����2̮��U`}@*>뭂 B[s��b 0�_*K����D�=">����'!0�$m��sR�߳.��D�Ҧ{K�)����v��P��s�5 w�J�Ѝ��;_�����>�϶ʙ(��o��q�!��n@8d��ӑ�ｍl}^"j,�P������+�y����Q�<�c�@8��#-�7��)�L���&CIQ���V��It�G�G��b_,v�>5er�4�Ǐ1C2�1�|��v����_%��Ņ��e�B���>�8��"��v�Z���.d|s{TTL�`�2����z&qG�-0`��㾊H"~�h7U�����b��m��!���宱!䶖�.�EB���J�k,}/�M�����9P}+H,	j�>o���݆%!o�����R5x�TH��z�!(z_<rP����+۴УN_,�M�T^R���!	1~4x�z�%�+) ����Y��CH��5�0|��,i0v�a~�~;Ss���9K[����m=��|ή?� {+�h���>�h,ʬy�6������0�u����J�N�6�z�fQ�����Q���fw���P+.�}����S\6m�o}����|+s�O桐��t��^���{�{N����!��I���j��77o*���a�,;c�H&�H${2�1�	J�J���+E�s��/�7��8Ϳ^��̐-t_VL����;`�yW3;������X6Eϱx�{�.1>��ت?~}�أ�	DCv�dbcv��"�	�>v ��"W��?\^3_U<r��hB/,h���-���~GQP�F ue�yU*�R��/+�P�{���Pk�!�U�P�,i*K���}a,�e7�}Y�3�n�l�$�}͡E~��2�u�|����`���&{�s�ffrN�"+�+� �׼�?�^��%
�TOw�4�чb��҆΍ ��%i�TM�šm
��3ʽ�bW��^�}ŃI��%_0�d�~�.�!d)۔ϚPi��!��pkg�i�������ΛB��%��2�32m,VA_�{!t����W~�:��p`
�/��	 ��g7u��YCVSTɐ>߬��{�n�4�y�����c�v��8�Q��2l9�X��N)gT0i'%(��/���JZv2��_�k$�h�pц->Om/�*d_��Q���|��zc�����;N}���Ā_=�m��;Q�]�u���"E��
<8Tn�$ܾ���
�u�c��w�+������no���u����Ԣ�GN��^�MŪ
<*_���:X{�M�Fz蚾~��O')Y�!si]�j�|:^)�0�v�R1���m/��Y��ϵ[p)��d.���V"V����)�������gـ�Q��s�U)���N�^��ܤ���],h��_�^p�q���z�o��u�8S;��Ѯ�����:�j_�1�m^#���$@qY@)�cۙg�F��?D�vuT~�,��g��~E7vm+7�d	��50�l�x ��_T���/�l���Zd�wn�Ÿm@5
�� K�`�������)&g#� Hab�xTF��<2�&;���Q"�^8K$���xM�Z���>��R���cd�ׯEH�z�L��&L��ɼ�$�u��Х�6[$��2��\��Sdk����G ?�=��g��VZ����Z�0yug�x�#h�����o��k��=���<νĿ������
c�H�0�d�}�g�]&1�[@B��s��9[�ɥP���3qy�.e-��Ŧ�B�k��kH��ćw�N
խ�2�J�nH�-�Z���2*T̤��qn#B��C9 �X9�D�����[Mx,n
�/H�m�F�W-lɒ�,.!�c�&ZG�ˍ���;�U�a��\'�3��P���Nt���B��4>fi�-��}NF��Ay�Ie4T3�l�mn���N���'`?���].�����m��hOܓxzy_ڮ��R�<�F��!�C�[S�����+c�[=p�k�F�T5 �������`]�pXk�Z��w*��~]nt�sU��H~��I� _qC 7BX�"�W�U��K�}�W)+&ꐜ�F*|�ؚ�:G��
�ŧk襝�/"u0z���[='�3*��0F��0����"� �YV��x]� w�`U��L����fD������)�?��w���;��|KIs=��3�q�Exօ��0���.Y�/X!>z���W'c��K@��؀0��nF���d ��Oke���avQpZ%3�~t���B��J��Z���A̯�}R��k�a�RU�A*g�MBr`��D=BkW����A	av	�'#ΜX9��_<� ��pӌ���ڭ��������F�Z�E J|�u�a_٢��)H^�iT��ѻ �J�ƈ�zӏQrh���Д����%��Y�Ӓ��K�2�=9�JLy$VR҂�y�*v�T�m�(��?���)�v����.T���㧤�����ݜA,gʄb	�$��N�b��A��~����;�|�������/j�7��<����&)ƫr�����i:'\�ϟȏ*h\�*������Y�(�~�_��DRis�)�8�� �~��i9�Q��YB�d��7�L�zב�� ��U@(�<��B�+��:� ��zx�p
(k�>������yId�U�0c���d��aX�U^tc�C���2}V�eI�������j����sb�s]�Lf5Sl_F� ��H��i 7�r�c��-�O?\�L����)h��r=�|5{��n�}sW�u�Sn)R�Ǐ��'��Mb�d?��2�"�0l�˂1P?̬D���2��=� ��x_���jV������S�0;VK��H[���z��v�!�Qԟ'���;�-���Ď���[�`F{�閙g,��qu���N�W)���
<��]Z�Cv�0�ܫM���&J�H"�r�D�i�y��J)--(��B�*5�ۂ���6 ��f.�+�>]h��=�}�c7�唤������!̿øGm��o�GkqL����Hk_	��Z�ߒ��{�!�F�����ߗ6�0��k�h��[�0Rx����8F!m��mc�7'-�~=̧O���=nf� �T�F�ڟ����ps�4:�3e�������z��
��I�l�+)Ɓ��x����4�(s0��{�Z������B���z��W�Ģ��>����6$_Â�B�01o#x���>˕�����!���-�yż-�m5�d�˭��1�j2�⯨�a3��m�d�����|'4��e?OO;LP^S-����/�&H�\2���!}B����l����N�!�a�c~�i>�](��ɒ�B�/cV�Mu��x	�J0v��j����~�'D���7�Ј��)ZK5����6��!�8'�ǥ@ۼn{SG���(�#	$)щ�t.Qj7{U��H�B&�mx��0[ҝCf��qt������5��ǻ�#���N���9���7:6w	�m���jg��I��K侾nHｃ2֭$�j�&����xvC�b2 Ѡҹq\�\�Y�\k]8EE�w�"O�6���8$Sc|Xڛ�il�����H�5�1�M�$�پ����um/�BBJ<o� ��T�c�MK� �k��(�Q2�����I&�[��<1f�<@���9sؙ_��n�̗�f���rbNa����;�Y��Fo�WQ�op?��ږ�~�Mȿ�)CY{Ŷ糑��}��A
����MX��h�>=� ���`_Щ����~�ՔCֱ}�0�J������i�R1�?T�Y�K�f?L��k߮�����05w�s�`#�p?f��o��6X�S�	OH�¸t}3aNz3h��| �����Ȣ%�'a����2�"Q�G�:�\fZ�ߔ��%#إz�gf�%��T��{30���G��Q�S��Q�ޱu��GU
l.w(���������0>����[��r8h{O=n�?Y�_�o0�F(�B^���	��5��<�ە�c���ܨ��KA�)���V��s�p&�9�3=Z���C#�ԁ)]~�Aq��_U�{�ł5����
�+��p����&����o�֓���"D̙��[ s~~j'�?� e׳�(B�RN���8l�l���7�ɋ�r/>�l��Qx�������̇{.LW�J��ဪ��َ4R�����b>!fZ��=[����[i����w������]����x�z�(�NZ:V�aej�}��y���S�$ c��(�zT��tk����X�U,#v"�f�D�����̱Y������X����ɿ0���0�ݏjJ�[�pWj|�|\,�fDl-�8�ج�ȧ�E� g�C��XI��P��Q91e.��\�P+��4�l�p7���G.�N1��\�����p~���~�ȩ��v0z�T� ��ƹ�K��2���Is����0� ,5�/�[���'X��=�=����z|�S Q����)��֤�dR�����BU�_�w�+X��#��¨6�ʭ�<N&��(�����S荌{g��Əl>,s�bY=��K��7l�o����9�D
C�i4F���8�ϝ����s�A}�cU��}�+�j��6{��:�	�a�.�Glm�Γ��ۖ$%�x��s������(��4]_��s��T�ŷ�Y[辍���Nmtiv���H���
z?VK=�]>�#x��漢���}<)���Iv��]6�{��m�a��v:�n�D�q���[u���"����Y�;D˅)�^	�N}.8�}�G�,9���	��M��7�.ǿA��
���Y9�\D2���7IޣR�sia�UA(�3/���r��,l@N.8)�Bvo�4�`w����b,?U�>��.K}@��N�-��?HNP1.��V
��`U����r�Tz�)�m�[P6�%�Nb
�"C֘�X��ĉ�(~�	���h���K��v�n��K�$`[\�1�;�z)Y����n1-�+q.30�cp�P�g?�l�?&|��W%�f�����KZ�����0C���� �;��L��eۨ85��fǐ=zo±�R���& ����m������IJA�syWS?&�4�>c&Z�K	��x:���h~��@~5����.e��~�t�a�J�������{Y�%��ؽ��w�t`�P�+1CW��u�����Oم7,�Ȍ�^��P|��d��S�!��Og4���\��o'Z�6�D�?�s�$A���q`���x��.GDw�^��vl�}��*�*Y�~�f�YG���YB�U�U�1�]�� ��	|��&B���L��_��㖃�M��᥮�D�xK$r�B��wI}q����.�	dZӠp9W�4��e}�w�,y�R6��ve�a�@�Fe����%�z P�ݑ���S%v)�wf���]�{����hP�ᛍ�5��cR�Y(�<Y��[_-N$�A�yu�K�����\m�	sQ�{H��I�i�L?Hem���H��}�w�lT��|��o)��T�*�F�]�4Z�ܕ��Ӹ�0lX9҂rf��9A�������m# ��f���2���7��M�:lτh�3td Yʲj�H�Z����$��%e����V�a�"�oɫ��7k9��<�����-1N�.�R;%2���0&:�/��M9�Vu��g3�i{[26*�e�I4_�S�M���ݠ�}��)c,��-s9c�2����4��ڐ�u��.٘�L*i���w�ݎ�ı`��~1��*�S��/�F�-i�Rm�IpD�'p��^�<λ��4Q�f������EM�. ��!�h���F+��:�>W����jp�t8�|���
���F��2ȂO�J0�!���F*�I�k(n������m�P~���,�G�9=� [x�|Y�A��E����2���#)��!U%��Qy䧞)g8�
i��@�W%���Հ$��`�`6m�F�M�l��κ���G��4^wV�[J$����A����P�'{1x�2��'�^YG%����2S�0.\+��]/�D���H�ڄ�c\�İe}�mV�T � ��'TH�����j#��p�K`Q��=�<��6U�҄|���@�����t�{k�+";Ǿj��S�nqv������S�Z�/ՋA>1���kUn���vΎzYg�7҇���0��?�l�y�+@�|�xm&Y;rd6kM� `n�Svw��u��k�K�ƕDШA ��o�9i�p9m�ﻭ�fM���@�k{�V������H<���N�Y��$)}��^A�ÿ�I��@�����[����_���ߣ����@�G^$�k���0t��ɬ�_��1�]���vc��]lhk6��e���F�����h8P[���|�+�v�K\���W�,�a��)jGT����sci7���u|H��,�ńM�݉��z�!Oh.���->;�����I�y,U�LW�+T����E�㨌9k8e�����W2P6�����w'�Nt�	K�o#W�ȪG�/i���cc����4X�|Y�Yjs4}���2q����;hf(ԛ	�ԁ?ABȖw�ܙ7��,��kz�V�<i~\B�S7����������c�ءKdL�~�����m��]�Q��R�Z�{P�7>~�$��l@��[5��Hq�a�K��g�#�D���2o�څ򢠺zX��,fC ������3{絟�������If�B<,�h��u�-��~UY�d�ˀ����W}�<����Y����"����@ ��"U��y79/��ϻ�T1�&��9�����FR@~B����l�:����	�$d���:�yd�����{���5��/Y�����M� ���$7g��ގ��PD�DyVuS���+��a1Л�����a'P㽯�fvgJ�ۑA��-A�������6�u!{?m0h��$9�\�7Zی���
�hAztvvϜL�;�ܐ!��T����X�W_�i����-౔hc�G���H�iN£c�>0�'!�FuPQ���b��[F"[PcC�z^dz����;�ڂe���}�n���)�M�~Q,�Q�5䡅=�i(�Y��\�8ƪQ�ou�򵅙~!`ظ��[�80�[�V�"c�S�����W<� ��vFt�Y�G.����<bY*�	��uc �{t�@�3�!j��#�}����*N�a�f�$���&�3�V��b5��Ǻqbe0wh ����Q�:�%�F�����7�&�g}�z��	��Ֆ���i���+͊0��C6��C��m��Am�?�����[{i�M4� Z(lG��ƴ:�9>������c�S�k��IP�
��#P�FXՑ���~4�BЮ\{��v�xƆ����8PN�2��	o�6���N������K��mi�_���!,�a6��WT��I��/�J�#/OlOc�[\f�@|�ߒ���(V$�FqW>'Pv��m��Q�>�,�w����^���M��(+�����o��Bb_�}�#ѐ{U@d��C�im�-���U�mܫ��/�U
)�E��x���h3��R�dF3�%�c��3��
?�8>��S�}W�䣅�L��k�W�e'�r��C���v���댬����%��n�����;�P�F�}�&RS�캘v|����H��_���?�`�����Ŧ����@1�
6+;�c^>�&oye553	
R�{V�1����aĜQM�2�����3��H-�$�'�;�������m��d��'ҁE��K��]FV��"~|;!��!(9Rm�j����W�w���E�f�(��������vy�d�K����nD�h�U�I;-x�xn�Gi�����[�30�Hu2L^���WM
��-X|?��o� �����_n$v_��ۿ�i�N��MQ�v�}�)�[UG=g��]�>�j4Q8fk�ީ:�o(5�C���KA>�g:qt����v����E���+��xO�/`�u%�t;�|��K�������2�%�����X��Z/b�Eh�"
�pN���U�j���p(x�O�ΠЮ�6XSV�S��7����m��yA�t�3)T��bU���/�8��
:�z����q�� W�5`8d�n��e|�`�;q��jc�)tջ� (�">-uaId�����5Kl ����E�"��:�g�`|�B��]!�����	ҝ��S���Ә�~��C�����¤�x�9�u��}}'�y������++y��� P�7CX�|'�4'7�^z�/m�-�?�<���G��i4a���{����>�4¢k���@��(SF0J)��a�l�p�@P�A�:�ȓ��r�p#�ߒ�Z�Vh����=�M	����Q޶B\?��\�Q�#p)��j���-¤M��.�����H7x�}��d��gk_�u�8'�F��}�fe|�s����S���s��"�#u3�_��e����%8~"��і��*�i�)�@oբ��Y�_E��巆DՕo�g�^�0�J��"��.�5]:�7䐣W��*�����nx�.
��<�����Q��lVD��'�	�_�$1C��	c3M�^�ѹ=G,WѴ����ak3�s��A�Rgb�������[�FMU-ԧ�/&��᳠uN�odF
��+�o��Ƣ�Ft��p���,���]X$a��x���ԡ[?�.?�̠,��F8V�K��pz��-�����<]Cк�z�e6�*i�ORT�:W��qHLQi%�!PՊ4�lA�q�@� ���������4����~E�t�f����:Z�$���� 8�?�j�J��ZZ�����B��-'���ؿH�ҦQn�d6�;#�/������۔��|���_>�-XQe�"}	���!V�e1ݫ�ȟо�X� �����5�>�r�$��9���C��n4fؐ��c�,op��6S������.n�'��1w�E�-�8���x��֥�=ֈG��zRɁk�m���� �x }`k�4U8C'R,[0)��f��`�]��q�^�L���8���88N�
Nu�ȹ��dL;q����k�x~����y�tՕPg�07|�V�	'c���Y�%Β �Ў�nR��m��W4\�@��3�I+h.Z3��$R��%���h�s.�!]'"\��"�����Z�yN������f�)g�(�|UYC0�n�_YQ<Vd��ws�����hp��ݏ����0q�ڸڢc^��~�����歅C�c|�2p0`�8��*�i8��}�Z��^�W�Zxt&J��~�
�F��['��_~��dҒK,F˦��,���k��D��"2n~[>�5zae��?(gc���
�6?jqdKuw��!�ćV	���{v)L��kx��h�&`ȇ����$Q�Hq.~�i�l9��C��|���t�����ʓ�T��|�T*Ȑy|b�f�ؑ	i�?X_��� t}i�l���L& �OQo��w��3�)^�=+g�g䌢���-�O��;B?).8���U*�:2I�!۰�V+K�O��M�V'B�%k�ު6VA��V��u��.(_���l�?�I(���|1��5�,�1#/J��̤:�����o`S�d�dr�|�J�1�q6b��]I�$N��N�⸦��T��k����p�|�u����0��t"��U ����g^^.Q6rw2���x@��'��c3��H+LT���u����4J��H%�N�w��o�`�D�����5�V:���D���<=@,a����#���n�h�x��Ox�Lg�|}���$���#?~��\���Rظ�o�ݰ�p�'U%K��@�w�����>��墱����9�e���|Y,�N����sgȥZBhxe���bט-G�������өQ��3�/�x�ʍB�h�H��Z�w���:�'�2����� �6;9F�!55��.����|a}�QZ�;�^d�5Q�8�Y�?w��C8��
)P�F�a���ւ�$���Q]i�g�^��ֲUy�`>����̝�s&P� �Ԫ�bB4�Djɜ�c~B�����A��qT�I!�X�V$��7N���,�(@�����;?꾸�����l��KJTߖ�B3=vO7J{v���|Q 'z�:ᶍO�E�n�k���nK����q�����D��r�Xr�$YV:M`=��`��aW)�K�������$n��up����xZ���5���=��c�#�
��	Ι�K�^�;
�_/Y�N�C��Ѝ	PsDy��D'�?�]�y�Wѱ-B	���%���y�|՜c��C ��Z���t��uq\u�-�ͬM*D������h�?�gX���)�`���	@Gے�r�b�Ŀq�3����Z��kfF��f�:�m?y!�a!��b���0�.��:?#j�:�z��j���6:K/��!�Nt3�ȷA�9���N��8b<ݯ�ۓ�N���[���v�F�t��ӾL���\0�ك�{���=7�Ө?��L���E��t(mlO;�sjB��2����[+�K��#�ޭ���j����������gY�ys���	�a�{�f�������aP`m
����䭓�]Lm���\q����4��i'Rŝ�E�t����ŀG�/mG�o�a�|**L��?����OQ�:�\�)r��xU���
H�!�����f�G
z3�d��dۘ��|qn�FL8�;xZOǌ4�~X�n�[�s�� |2�a ���`�ƾ���Ð�-%#ea~��5��:�EEt�I{�w"�Y�<��)l�vɑ���}�k\�7xk�j ybnǕ)eF�If݈��l�nv��LQ��j��^&����3 %4�Ѯ\W^haJ����k����703�uj��*kJ5��gsE�2X/R������ӎ��ImSQ�6�o���woW0m�3J���园�z2�g��"��H����K��+>q��ւ��Q�(��:O�+l7߰����L�'�A�O��`���"��E5��O�6�9��A��R�ح��qr%)����ZQ&'6��X��~�##�4vFè������\S��=�$Cr"D�zPL��A�u#�tM���n��9Es��¸�̮�g��:]�������������$����9��6
�$Dn俋�����+�XB�-�9��ڄ���S�����6�t������ϧ�`A��6� X���o	\�r͗(�����E�[>߇8��5���l��LJo�,cZ�]�HPҕ�L?%8tC�G�O���d?�F2�fˣ[}�|�ާ�-��m��)"5ok�vf����<z5ޞ�J�i ��~�I8Ah3ja�W�4v�A�&�+����K���(�l�v!�2=J�? ��@�)bg?���ח�+�D����Or��C'��o��H�ͬ?��MY�EѺ&_=�)cK���3�TL/��iHf �>)b	,�yҲY�Z9��#�ƞC?κtT1'=�`L���tt;E�f���.\I�;����U{��E#!~��6��=չ���ut��$���q�"�t]cM	�iTm����~����\���X���t%���L9�=@��iy/	ٙ V�g��L�N��'D���#2s+ˡؠ����7�����kY���=�����u�������Ml�乮�3_�$˙�����>���X��s؝����Gg|�P�X����8R*W�j��ԗg��A+��ԍ����ڠ2��v�f��O0-l�1��$��6�I�$(�~x3��uDǂ	����Y��zf�8�����[������*m�w�nGC��9�f��\s�'<�X�.�ͦ����>��Lo��5ݧb���&	��{^�;�9�+7J	^���g�w_棫!�0֒yza7�|�l�E�M��W7�8/��|��+�r]�6������Q��a˃�?����R�g������8!&�7���S�P	6ε;�����'q�J����*�`ҋ�nm���&�}�[p����M�U��%z��}�.W���Zi{�{!G�'�k�R�V�8�QU�"���VQ�>��g)NoD����W�e��|��R�֫<A�v��4�~���;T��6}Us����;��$�K^0�?Tfh�^|������A3��V˷�̲]�6{�%ŗ�(���=�jX,_�	�b=�ʸk���J!�Xϯ�+�mӜ�� ,I�����/�(QWrk�Vq�)Z�7Gd��lɸ�-��U��l��i%���џ+x�̳08+����G���3�ecI�n��8g��rG@�ї� �Sh|���T8��H��ma�j;)6����9�F��ն�/�f��o�*�����TDn	GɷB>Lf�
)w�%�y[׶+�gJ��X~��/?n����e��2��8�RbVض߀�e����h����/D*�i���Μ��N����o�0����"1��c�&@��S?Z��'��h e�ZϿ��YhW`�i�G6r_�
�y2�&)�j���^ �Ľ7I\��Oôqo>�W]k��o�be��R�Dor�5�� �G!łj'�0�&��@�k�(L�
�-�t�K}dA�lJ� ��@�Y�b�t�Vw�]���U��&�M+���h@ռ�ɬ;|���75����S�߆�gc/�nQ�Р��h`��b�߁��s(��{�R�]݁�`��#-��Q*_ mzP�mb����zz��J�m��^���"�3S.h$�A��q輥�d+��Q�z_�@���ۮW����IR�:��e2JV������ >@(�{��O)�1 W{���x9:���_G#,p��YQ�_g�!@��9����.��(VV�Q�J�7m쨂BH��')�C.
�1��e��a,����B���xj��YdYf�w�)��NÓ��L5���2}�u����y����5dNu7�sߪ�z +��!,X�#�25�'p��p��9���C�O�r�%5G+��W��r�x̚o�d5��	f@�!-�J.���������4���tv'T����4��7T� z}�J�v=ǘN�S��#0)� ���O�k��cхRc�N�h���;��f98��І_t)��H�k��g$S����H���V� {<����2�᣻	��.�6h��@7�!�mV��>} ��5�6f�J�mZ�@v��!wA���&���$M&\�~2�`aF����7*[Αp�i��&�Z��p��yb"K�"��9�6t�H���3����O�1����5%�x�ɜ}�����i}t�����b�oM%�{s	�QFcR�Ր�\��E�@̎y�]���� �!>��kr;��X=�,�~*?s ]��@�ݴ1���(y2�����@�'v�00A�(�˸D�β����+�{�g]m�k�m�'�r��&��n�[ [p.�v�53�&P�k.�`%'��XB���=�įxe���c�I~�d�H�'��!��4���0�R9�&��*d�*ָ�������|��Zt���꾣aq�������OB��;HF�<܋�xG�.82P�� ƕ2�����eQ��GLɅ�#~3E��>��^s[�a�y:����aC3��/~�/��	`C��_�+�m��Qa6�0�Ko��J%mN���A0�
�c��Us���F�z��!iŵ=��A��^$:e'Jf�:��c�F�1���UH�8�e\Xǆ0��/yq��?傆�� wO�,�Ȥ��nJ���\y��î�+�ƴ���#�0���2U �l�e��!�i3�_l_�� U~s$������e�<|�;G��@�4���m�!S��5��D�K��ew��*
l���刱ۚ��x��ί��ւ��^A��8����k`%�!�΁�ah���9��eL����(��u⋃>��S����I� �9~�B��,PB^"N�*��-�j��ӳ�R)�1�W�<�e]�NuUK�K���·���nQ�U&��6E"�J��(Ǹ'X���#�l2���┙��B.Z��j�㙑2�P*��*y����`�h[�pxb8����h����q���[�� ���ر���y�sO
�|J2�l�nGԆ��@<�����3�B��FM�v�CC���wL��%u�ײq�l8�/��}]�Ȣ�cC�qdad��d�E&�OB�x'�����g�!�xM�yM(^�3�>�W�Ǘ�I�v������.�_8s�P-�g1S.���MV��N߭>	��%s��yZG�Q�xW#��&�Ht}>�l�W���C�Z�z���3����p(zE�{ ``�1~�h�i(�L�P���y=w,��jn`l������=9G���c:j��r\�d��o�{��7��57�fC�Ą}2�����B-�K+!��٬������j�ݣ�v��ǮUp�;b��/��\��h����*�r�-�� ���B���]m}:iC("�0�<�¯�ܶ�D��߳t�:��j����L}����_�����"J�P!"aŸhp|��p���Mb���:�o��ab�o{����/�q�)'�&k��A�N�Gap��+�Ȯbe7 �t�%T��0G�)�OQO��Põ��c؋�q� �S��f�hze��h�4��T��[�A�A���.��1��)����M�-�IVٳ�₷b�N'�L�*`ऱ���:�B�I�u�f�a�9�#�T�������f�9,�rZa��Iԭʹ��JI�~'���K���`W?k`^!���0p7�xe�����+K%\曅�F� ��cή8� ��P+ՆQ��Z���稼�K�A��"��f^�v���q�(���2�Z����cyR!��+gYa��.��*PT�.���H�V�%x�\�D}�����1��y�q\���ah��V�E.o���}�)�� �_zK��X�^\�2}�mAF�{9�zo��$M>YV"��5��h��H)n��cb٠|�>Z������I���������ڀ�����rz��ҝ:�)[i�D�s�52M���/�����.UJ��	�1��	�W�ˏm��`b�v(��:��pg \ЪEvH4M���RJֺ,��߬8���g��ZJ	w�=��Q��z�����>��h�~2@�Tւ\n#H��>���a���,&}�-,�q�y�%q�L�R�+���z6@A�c�e�n(�#(H�8����-?ǝ6s����
��Z����@�6R���V.J,};�DR�d��-�q�aw5�Мz��������w��t=g�5;	���8a��s��6�|�c EY�����9�����E���F���=��/J��p��� V�ni���q�h��4 ��lJ1@��Yg+e�d��RJb3�V�{��Q�c�n��ٱ�j���� �5*��ĦN�w�&)഼��>̵�/�7zNą���	>���`q7������o;`�u�ϝ(��e�2��x�Gw���HB��/J5
���;��T(�D��ǆ����G�\��?�ʔ�\	4<��v�ῠ�d�w�d�d0EȎ�7!�z
\|CW&zk��}��Tl�����>�x�pJ|A	ҫ�����}d}e'e�aV�;�o�4�\EF*v�3w}>�4���`F��4�CcqZ�T��@��%�:�8/�֭jт-�#���`�]g����lq �>�i\��8��4�f���<N