��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����F��':�ޜ�2̼ߵ2D�c�k	�?��lK���ګ�6�6K���}^��xF�u��hkp;���j�n���WVܫ� ����c������jɭ�L�5}��>��<L�=l{��	�Q�D�\V�d�s�囏���Qz��
2W6�ol��hX�| �/������¾7�z)�5���KUo$��bv̛�EQ��e������Q,L��d�tӬ�7���Y��]7�9�MD�vD��g:����rz}�|��x2��8R��X}&}R���)XGn��l���LUK�3�s��,<NqǬ�l�ٿ8D���qd]_�#�c){\�-�э�dK��N1����y�~�.�ߘ�c�� �]ئ��(�����Fq���-���F�e*9������
B��1���}ͳ[��y�?�,c����}��O�sW�Ɛ�ö�i K�lĪ��&ެz����Ò��$hP�?e�=���D���>+�`9��_Vs����͎�/'��I����_���s��A6#�3���h�<��J����v�F�8�2�Y�h�vhm(&��N��c`i�#��+�4�6'�q��0���	�x �Y��c?�g,�?���^3��HŬ���������o���5������x]�9�[���q��)Qp`�R,�ʳi����}�����Yz��r��ʉ�#\��-���l����g�CF����g�uLx��f�K�jk��Xs�ǽR0��Ub����� ;*C�ٲ��^�0�X^&I0O�8�h�V��M~q��J��(����4M�
�Qa"��`H˦���)�vtť��1��t��ʭ�F]��-�ƴ@�k!�o�ܞZi"ٵh��P[ę���t<7��Z̵+Kmߦ1��%#����M/դk� wp�V�*�~ZF禞g�-71&7���:8�e��z�8^0/~"e�`F��fBE8:���d��_!}�/����ݽ@o�Su���GJ|>�����kԵ�.��e�c�V ���� ���JH�I��g�l�D�y��v6�h��}Г�����y|=�MZwO�{�wI��O#�.㴤?��L��k��Pxx�4����E�=T�Ӂ|f{4���:�ܱ�?"��E���<,��[�]���t�tN��l�J�:�q��%!xg�C/�ݯ��b�~�w����%텟�WIQ��)dB�3��H�{#�~�*���j?��H��y@|J��۟"�r�R� ��>�r��*~}u��*�$�K�o�؛"�u戂u%��8d��*	'�u�u��&��?���)�NZd�in6(�P�+RQ�KVm�rN�G��3�sj8����^�H�
W{}iR��
4aE�F_�������\�%'�q{g|�F^lI�Za��W)
���10/��OAm.D�HB�+��V:�������޾F�C�	�Pyn�f�m����9Y%�ELː1C
*�F�~�"�<_�vR�ј����~?1����3*;���M^F�£��x����h[�E�'zJ��(��	�
)�P��N.���^MHԸ�ƛp ?>�p�8Ѩ��
meVHi��2l����~Pg����;:�����|!K�=F���F���b�GZK���塨��4lo>+e7J�Rx����񎉤ߒ��:Tݺ���i���ݍyY� ��؀H��m��)���q�ԢV�?��`{��	��c1�Fz�.z4���-N�q��]�, �'y�~�M���v��-�L(ۑ]��"o�=l|��Σ�G�j�	��Mn�0Ƈ�?r���x�\�Ƚ-��J�*��]Hlu�I�}�[�U��:y�X�O�ں���&�=g�,�6��X*�P�gy��=��˔�E[��\i���I����wR�pèAW."v�y�ءR��C�-������3������,��#��Ğ�32�q0��E,ܠ�[ �/���K�ݳ���2 *uk�O�'���"b=��c���<S�;.n��"�,:�{@g��?�pK�y�P�my�[&��=\%Kd�i8[�:�-��v�8����[�����t ex�c����D�N���Mr#���@��NzI�w��J�  ���ҰlLCM��d���]S[ӽq�k�H����ܦ��y��`�z����j��3�ȭ;R��q��&\!J,B��X��k��|M����\t#��RN�\3�J�~AA����
�/�ňy�zɾ;8%#��0S+@x0nҴ��T^鷙�g��fVGd��"�O�8V���Ih�#f����+z 7������W������9K�*��U��;���.�b�|fv�++lr���CY�,GV�:~�pF����%߮LmX�[�[<VQ�:�&<3�F.�����!��W��Q� ��2\_H���r�2!�JNY)����T��T�IJ�����9��?�J��'?�G�# A���&�-u;(�a{=��V�<u���ELf������ϗ��T8w�J�����;.��q���b^mT^Q1��m�W5VlG�^˯�v�.��\#~Y�����&b? �dHY����`⯛`�>	I��88	f�.u�
�l`�d��n����s"�@�r�����h˻Ά/����	��YAI������2I�~�� �P���Q@9�҇��!K��@͏�%L��6�DNr�j+��+m�_$8r���v+Ewr	��?�Q�j�$&�ۨ�>X~��Y�TS�C�tO���\7{�2���E�$��)��6#a��&�l����cNLU;3�s�I���HD/��uG!��u���9h��1V��;�3!���
�?���o#98t�`�)�����9�r�ج�R�ꖛ���,Q+���w��.���(�"�vAK��a���H��϶�7�0B �7al��p"Y�m#�*M�Wc���}j�nD��e�7�U%ã\Z���� n��
��%��Ĭ�.��ئ�{0	D芎�b �KlׁE4w�e\�p��9@����ޫ�ZP&I�'�z�UQ��-��/u��m��O�}�p�-�6p��Jh�A�kk!����(�� �Ҟ��>�$�Wʟ
q�__��6Y9���4ʩ[���+������1�Y�Eϖ&� �~��Ճ)�)��qU�y��
�K٨AQ�F�{��rl[+H�5kڃ�3ť�Dv�ø�4'�@��fr	���}/�3�0>�?�Qx�.6�Ab�W��#F��m�5�%���!�=Ӧ	�z0���-��!��f]0��ѰI�`������[2���)�_*{�_����78w�=Yŋ���be��>�$��)��n�} A�Q{����f9��^-PBS95�Ț���xh����Z�#���K���T����pᙞ�	�J���$�-4��KEw �����kټ0���i�*-�/�K�;lh�u�WF��ghj���PM4�Sx�������69J�����B�m��ErsG�
��t���BA���"{Q�wW�SI��D��4��QP�4��)!B��|
���z#���u�r�U�A!VT���W�ݜ�fCP��o��*z�\�5򒑬f��E̫ 	�����yMz5��_�����&�-�ޓ�);.Z7���� �����%I�u[h�Nd�K깧^)�6m��E�������$���eïx>9�Ai��jF�w�}�׿���3s�a�T����;V�	:Ց�w-4:
g��w�Y
�5V�W��"���vG�s����',��T��8j�$��u<ɴ��Yj\��.��܍�m/��F#z�\�{f#�@���������׻��Dl��� !w�%=H�	�(L�Ж��4�p�k��@�Ƿiw��2q>'����m��o�]�E�Wղ��3�Ab��901q-
h��f_e_pE�zF�v� ��9h(��Z"g�4*�%����&@,�\
��OhX��7�]U|pT(��lw@���Y����Ÿs�瀂��q��O^ J}\6eV"�����~h��g����95����x�ca��lBV����d!���7��t�r��+\wwosቆ��f�jO]囄B��i����6��m2��_.CC|�UE�e]������1x�7���d ��R��JF����/0'	�#�����YG%��%�)l�Yo2E��˯�F�<�9D/k�&zP���g�1�F����+��ɗ�X�V�)R	n�����: T\Z��d�� q�j�qF��v�4e�.���i�kg���5:"����Y���a}�OQ�<32������X>��Ɣɲ����Xk��G�h����4<��=��Ɨ~���*����>��_��6�Ma�����{	ja����<~����LW�I?2�� nl�Q��E���	�C��E�[�P�_Y��[�o�1�ԡ& ��;k�z�O�U�r#����f�W��f��NV�G0�L�ᮊ��u�͒<�l�@�I��p��j���m2�Q��i��|,����R����,�0S���F�\[��jxd%�*y�CFK���O�䫇tSh������_�N&^�1m�ۣ����E�%,{�Su��,�<��Z���qi�qN��Xq���.�DJs�q�����f�Um�+��Һw	e���[c��'�9� �)�(�-�4�k���7�場pBv'�2s`G��5��͸W�j2�)� T2���%J�(�������4)N��w�eJ:ɥ|f�1�/*cn�2��"���5����xy��Y� 'cD�r���-��%��9=��(�M�A�É(/��@�n�Ϋ�fƀ�W���.�r8�J(�&eƨ�y08E0���ݛ�M��$P?��o���<�r��@���@f*�	8�$�
=W��zUD�!>�޸�&���{�B�2pTj��1�#B�S���]lw��t��т8�a�ÁH
 �  +��C)4
�s��djO:�9#,,Ո�vP8㭦670t!N<rU�=�P�B��kc"�3cL�Ad+�U>��>�Kta��o(e��G$fk���G��4���eG0�J�C*��BZ��iKG�@0E霵@�$cR t#��=z1m�o�ҝ���U<��%��R�
��TR_���x���'F s'�&��l���f�uuEHz��TGO�ⴈ]�AP�U�fcV��ã�7?Z}�����@e5���$��tmYäuo�Kؕ �߁Y��ч�j{��dw�%OsrS�Z�ˤ�#�W�ǲ�|H&�ȻV�.F�.�(��8���D8:�%� 0��N�I�'�&�6�m/F�p�m~��gW�W�O��홯XvXu�"~��R��Y,|*��r��7 ��l'/o@���wy���[��^9/�S^�HP�=�1�Z��H�ڍw�qǮg�ҝw��^����5��S�`�
��|#� �K���L��=F���/��pYb�^�v(j� �U�~btx�M�g �Նm�b����VP��8�k_)R�W���� tD\c��k@<���>��Y?A1�X�p�jZy}�xЗ�XȜTr����kt\r������ʰ'S5Մ�-�D �a�e򧦌+���aF�>��
�+B�WG�u
yY$�]��6��^�O���^��Uk�+c��������)T��ٿA�z����F���>����1��0�*�"�.��a��=Ȏ�����c��E��"8�`
��'M�ћ��'�GG�L!l����H��i�M���`:���Q�&�g߀�[�[�����`�y+���=�]���Q�J$KA��`����2+:���&�w�{Ԡ��t��귔��Q�h��|'.]V�M�A@l�����U(9�e�kG��:a���X�N��;}�����k�R��$���:<�A����� Ut4]�����/������K\۲�~���fo<�4�����Ok�����o�ȕ�u똧F�jv�" �ө�$��ċGOaՙ��X������|�H�� Q����+�����rI��*�49���X*�iJţ��+�-��E������"ϔ�)1YH_Mډ�9���	#p�ΆS��Oj�+��_A�&��GɌJ��Oú	����~�;��u� s�f�#�m�E�PTL7�#�B�0j�"9���Mʳan��	��{�%ӕ�����r�SVn�:�o�V6g�q��(���Wy� й�/�,G�!���� �,2�q5'1��gK,�r�v�=L4�'s���`H� �q���w�~7!� f>g��I����>���s���wny�U7�f���5�2�1�Y��Ȭ��k��ʷ�/���Y��͜ Eb|�+�)�B�ٮ�c�.����`r�s0��i�|��צM��md����!]��u��SR�� teQJ��v�s��)^��Y�ތӇ����rdEWw���j>��g���'B���k�S3SZ�e�0:���%�.����ܕ˙:ח�C�v��9��D�!Ww�o���߂c�\B�ml���Z��� cBx��cZ�������.�N*�	�ͯ����ֱ��p<�Q��o��i[��[<����a�#��:�?��Ϯ���ǖc��t@:��q�Wf&J)9��gE��y"�uIX+픎;y����J�䐄 Q1�HCsz�ԍ�O�����Ae �x%�[�%$p� Ix�����N�v��W��Ӎ�<'Coou�Ӕo�x~e���Ҁ�-C+Ac����(L?}�=ÆU"E���!_�u�j9,��%*c�F�%�/��\C[8��l��)*��=��ː׼�ő����/͌��f�"��E�ԝŨ��g���j�i����Xт}�!����4ϼXr|c��y��M���yl'��l�g]+(��Y�^�b������S�B�,_E�҄A�Z1o�j���J���7OK�n�]�I��Y?�@ƴ��V�x]��+PH�����u���I�Y��č�E��>GW���v����῝�>����u���c���f翗���"^�qX�mIbH�D�ma���"3UJ�`O�<�C�ne;�y4�<�ѻ�I���iW�Wr�X�9�KP��lE��j%���>�ܥϱsc
x��X˾���΍-y�H�`۩2�ctBU�b!� ͮ�(]���!ߞ��-�-S�e{8�~@�Q{�{�x��� �H��h��gET�||��z�2��)�o���N��,�:�y�g"4�bߠ��`Gta�#%��vpCq^�������Wo��O ^���鰡y5�;�?./��g��R�E��:ݍbk��aya�ͼ�n��&�9����i��D3BE�{������`�E��o�R�~�����~���wN�;nJk����u�'E�-���qz��!b��Q6�8��=�A��w�lFػ��m����]�~����Z��3���`�E�.�R�`�ǵJ���oE�/.��Ќb���	��C�o�K����`E:=]��/J�~y/�DpGv��=�: Έk��A]��6�����PjYr�!kKH��H��Kx̉��qZ���N����cyP�m���T�$T]֙�'�+#�6	�:%�8�!�t�c�XM+&����r4W2{߄,��0�yѯj�D�o5����^V���!\�� (��	O��5��&_���93&���n�C���ʕ���*/�]��"C��}���{]s7u�,�O���b�[g��a�%�U3�=\�D��>&���ysn�,�Hd�wov∐���m�l���|F��n[6�JG�KQ�c��
|�F�N�E�o��a��u(V��|��'�WV��o([�m���8M��a������CQ	���z^o?4A��q?�@�4��ZX-�{d���ݎ�b�(��U�2�sx����еM�{���T���fw�ƿ`�z�^�_��	̹dB�b�?
x�G�"c�����J�����!�j���[�6'O�@V��ͧ�r��#��8���{������{���O8ݭ���"\f)��ȒK���*p��7<�x5 �2�9���� a�n0L����`hHƱ�1����#��r�q����w!:��<��'1��#!e)C\�e�{m��e�Q~�1����:�I-3����b}����%�R�r�M��g��ຜ80� �}��/�f3�dc4����Wm@�*��3X�����
@�o����-<�㟸��������%9:�Qdq��-���j3�%l�>��O!1��GS9����A�����k?z!��g��7�{�h��+�\�G��ݛL�+0��.�z���稢��҉3�����F�`ը�R�(�'I�{lV:��H=7:^�f����u.h���x���f����X����#��w��R�\'�b�ĬY�A��1��G�]��]uyy2��p�*K��N��jG��	v-!�c�s-&0� P~��p��L�F���*���M��h�V�᳼�<G�\���^��M��\��i�U�ɩH��%�L��B�&��,;��C�"v�Y_���i�\\�K��}�iw���K��e�8���Z(!n�`�b2w��|� 
x���+5_��Y�m�,Ȁ�a��Rɯ��������ݣ��ݖV��ͳ���� ����ut<x>i��#�8�)_A-���m;̔󨯫S�>@=O>9�Z�6@\8~C������:���R	����u{�*�ko���Yo$m��z�߁�*0�.�*u �ٛ~0���=���SNM�(?��Ƥe�R�0���������dvNp���4e����M�m޵l'��[tx�ѕ	x�8��Y/�����F�6�'m������%ب�N͹6�M[@�	�p������Qx�?J�#G��]�^Vt�	H����ο��T�FN�E����N��6�Z����/k�y�^"���i�ϣ�?�a�̝���'R`La������=�_t�D��@�鯄?�b����z���V()�g �b�ߵ��d�:��wi<"4���Z�(�&�!S�K\ �\s�� a�l;`4A�R�V�ۀ+nf��KKaۛ��%ptg�>
{*���&�_�$���Z��������oN�2��6��p�+�(0�s��Sk�S��g�D�m�y�?����2���S�ԱU9y��Z[�ڔ�]l@�'�������W��'f�{�m�"������*Cy;���"{��e!����� z�q�JH7ɉm&#�2DSx�專�2;�a�{�ާNm���WRM$Na�o0hA��q�(@����w����"�a�|���Gu���_{�o͵JV�j8�W����76��S"� մ`{�y���l�ƿ�whm����`�$�
6D�_����W��xp.�#�)�H�f11U�z�~l:�ܦ1�%�q��3Gb�)Vw 3�'ȯ��QN��RE�*���e46�lO��(��2�I��d��(X @j!��u�ƫ�tvpe����|iE���zl�'	dwS�m#�P3�~�i޹O�"q��״�_�@��1���3%�Z�1g��)(�C�J!��t�%��*�~(�c����Hͷ�A�_�h���w�fA7���
o��\��0��0�x�5 P@pB��5E�"9u�sU7tcȻkʌ��c��z�]�5}X�X�W�%2��?N��D�e�񔣮��0��YL�ѥ eT�+=�i���Ql��h��
���5�Q"�������ae�K�h�nwȎe+n9K����.�mX���#������~P�+
|,<��@xμƌ�Y酙��T_�!E�֤w���ëm�ŀ8��)����.|s�=�	�M��;]��X�0@#F|���KO�X�׭�tE�f#r�/!�q�	/��ߝ�l��%e��X�;� 0WJ�Q��bӲ�'�#U��5����w҄��7�s�r+��0�����?bOՠٚ�OX�_��{�gAssDX\�>U����Q�0-1�/����*B��?���ѥ�U����
-��ڍw�%�y�'7�ћ��	�����B�GMdٺW�/�Ӆ�Ⱦ"@�|@��M�6���^��$�����! +�����k[S��*.���3������v^��f>���=��R L�E��o	��bvu�� N|m��5�k�?qA��m(�ID�����#(�������s���8�:i�h����� �X&� �ʹ����ُl�%:�7V����T�{���]�9y�O�!���b��%�.UŔ�S��M���zq���;�k޿.�@VB<Ŕ܋Z��������z����z�hGy���PwBb.��}�J��<"h����-Q���^�Mk�1�,w��:SXƿ�lK�6՗W�N����� k�v�/�ZI�b��#��J�]���������KD_]P����Z��U,�m���X�QO��`t�`e:E��>}�Ҵ�×��?�Wq�hO�{�ۻ�_9��R� wS��&�|��z2�<�λ[�^���D��:�m�&���"����y`��h��'9f4)���]
�1���C�O��ۿ�#ZD>��*�7]}#�s�}��?ѷ	G��8~v��ig�;���V� /T����Mt��X|�d�S)���qk��=b���3Eʭy�M��r%��Sn����G�	�j����#��x�tѲB��_'��d�_;V���R�dQ؟�w��
��"��?0���p��7�3���T�Ad��Q�]���k��k�6�A��E˻�{���f��!� ]���0�5h�9ނ��HhI!M�eć����	��*�x�$�/�$�p�+�a[F���W�>L��a�/�|s�zَ^��D�iw	�d�%��]���/�P�?���i���k�ٞ/�A+��ʪ|b	����Z2��{�ԠhWkZ���h왤\l'����<��k���yI'����Y�[�F� {f���sg3j���e̱$QE�y��
��m�ǯ��w���Q����ů�������������R�JC�v�x��PYsH}Qu��a+Yd+]	i���8K�I��A?��čͼ_.w=�]m;�i�C��������.D��������[��[!	c��!��L	�~Q�#M0��۸:�(q�&��H9,�p�I��-��k#s}ܽj1r£x�yŠ]{&B�\���'�i�~|��lǪ�[�e'�|I�Su�Ħ{��SMS���O��ϔL�&f���n�چ���:u�.3o@�W[T9���idq�L)Y_6�:�qpt��-j�ȥ.���ІjUQ`�W��C"X��c��=JV՘�\׆���Eel��}޲��f���sbE�ۦ�t�tP�W�~�!Y�-��c�\p��oA{w�S��MAt�B9�Wh��t���sT!�g@�s�e���S��m5\���ۮ|B��Q�Gv�U<#�~�3_ʒ���6��㴍sl�dۻ��Öɦ��w��QOfd�{����9�NҜ�Zr^�Ey
��/�%�8�nL*$�=۔ƹ�q��s��B^o��kڬ�V�V����>:��ޅsSs|?P��<��[(J{����]!("���vG�4��q���`���.L���G�IÁXHO��ތ$�!�0�ֻ:+�#�`�N����:��/<iG~o7_���].��-s7�NOL�}Ä��m��&�X��;��-g�;O|Pz�#M��T����'O����~h���������:��J	��T�@׊C��ٷ�qA7~��:� �Z��)����h�p#c�(�����Ϋ4�j���Y�?�$�p�+�yfp2G��:G�~L쑉fֹ�'��ϰ�P��e-�ȒD� �VIs3��XH����{FE�Go�'��t!��C i���j?��lc��i�I����X��u;�k!ljyi�3�|�C����l���"�+P�SW[�Oт7�����}��:�[�gj\�w����H��%� ��S^o ��St�܄��G�F�)ó��E�0O��n�fZ�- H,׳�PXU���ho_c�a�3]�����E��9��E�s��s���rqY�i��T���f+��X�好��0������#�{%��6�@�4�җ��舒� 8����t.�k�=އ2{��N��O ��q�]��Y����#�TMUw����qmQ�4�A9_�4�j�^*<�r�I\4�v�o�-110,'<��]U��P18�+���֖]�����?�N�;��Jr�V"���T���0�>� xa���H��Ž(�}q��*h���N:E�y���l8\�7�VmU��o��G�-�Y����3���C�Gh�R��7�m���(-�Q����2lr�D����^<��*�L��M&#���i��@m���L49�y�ܱKAw������m�_�B��c����K��i�U�}��f�+]� �RE߱Ю����=ĩ�j�������I��8x���!|+|��5cI1�9�3$�7nB�6~�|���X�ID;���U�P�_�@w���@��C��{f�և���h����2�X����/��T����X/Z8^����$1\e�,뿽�J
݀�<�j�1j鏿w�s�٩�Xv���H������&��I��n��@�|���a4pE@�"%�,�qY�?�.���+
��.YǨ4>9��!z�:I�s�msS�x�>��O��%��MC	��yf8F�>��u��ļ��C�I'�w��5m$�m=���4J��r!��oY�`��K׀�c!�ڎ��������lV��>z#2��%��w�!�3�Y͕(g���$�]
C��Aާ�	lc4�M��G롡>��ΰe.�A����-Չ���D�@
�Ɛ�ٜ������\�b+��{o��ua�O��ψ����9̬�'�z��o��*p�����KoM���e��8[�=�*6\�{0J����ϺʉI��@�@�Q��Q�q���X�ʷ��^���o��������o���s�*Ag�X�˜9�����Ǿ����A�v�p���u�$�?��rPm~��LmU>S�5T��XR����I��T��@�aI�PO�/��dkm�!7��t֢#W����,=\Fz�-�&����B1�]��J=2�M�:�BH������� �)�D[��xq�������5�j�N�g��{�����=�y>i�k�|�Ǉ+=�.��j�BT��y��&���%U={�d�~�(\�o;��`MF�>
�9�6��e�'���0�b�%�rK��%�i����mc��d>/�Z�|U�,���/���
�2V/(XnĴ��x�1�&��`Fw>S��'�{�
8^G��0D,5a�}p'�ڧdᭃܷ�� �n,u]Jp7��{���=i�Җ)v���/ۊ�m� �����|�5\R|�H:�ʖ�����^r�jj�K�{l>�G2��K��AI"�@���^��3���;�25$�y̵��b2�EI/���J�P�v_#]�&��6�B�'�x8XE][��X�'��g�[WB`�>�_�/x�J�%���1�=4��MXnI`�r�y4T�)�-"5N�f96����Ń�`�hO5��z�������)9_8�%�X��C	�8��)�
j�M�j)D:�\Eo���i����F�\�l� �œ�h侸B�NY�	�f�LNMw^�<�$i�8���w~lqͱ�3duȅB�޸�Qq<��A<����[B���$Z �#&������!���h�|��+�����6�&u�{PlT���f�����BKI6\h�M���WJO���\J ����N�h���~�O�5lDʿ�����ݰkS�3c!G�f#{�������C��{��q�I�תx��6S�9���K�́�O�8����4�D����y�Q�Q
ڌ�y5~��qt��@��xaxF|q�*)ŝ��Y�{So�c��r�W|�&yT��FaxIk���3=��&�d������J���Zto$��6{9x�sB�%lR��I�5>3�'�1E�ߧ{=r����h��0?�
�0��٠��t��{k�N3���|�=��6�`����/��nK(��d�@�-���;~|>y��|�m��6jb(>�i@�C[ܤ��������><���쯨@�ǐ���S�(u�[A#�T]-�I��t���`W������f`�U�6��ݝ��-���TM<$�kI���Z"�$�{�抂���H�PE7�@����	�S�9� �&/d�$��mZW��n��v8t�YA�:��o�t�ǋֆ�#��Ѻ�m#=��T鉮��x%;& ߬�M����)7,�g�1��z;��i�p�b1�,H]�4��~d���Y'�(�27o�.T�LԜ�D��y��d��	%
+j=�H��a%���T�]h	ʼ�
a�M�^��W�}���GYJ������I����RU�8��z�*���~F��BӬ4������@���z�L�Wƅ��.�%�K���	�lYIQ�9��5Y�k
���-�����p�~�������Ź��.��o���n��,�rz)Թ-�؝�вHU(���߿��14Fw�[�q 3�\���|�������
 0�ZB1�����/^Ѣ�U����c��*��R)�x�JD�t��"4b�QwxE��8��3������&Qz�lJ�72��bLlL�Bj�c��%��_OA���ަAY۠{^��.�1;��a���0O?\ّ�thɥ����ve�N_��x�f�CcI�瀳^ͯ��j�y��G���Qt[%��E���{ڲW����a~�/��e�𾔎��q�����A����*���S �>�����2�?��:ujز�'��OU�oa�R<��=י�W�C��Lq4�G�{eЄ��pe~>Dp������d�f��0��ͨx�k*x�\ݙu��Ԇ����M)#�:X9R��
է�U.(P+ݨ!qS��^����e�@V/��5�\ A��S�=��F�藌	�w3�[��[t���E.
9���6���^�����]��j�T�:/490�
�����a�Ee/�����t9U�^'9�h��!Q~Z+혔��l<kv#�b{����^�2�#d)�a���f�֡�f���
}y'3MA|.��`��N�*B�����!��7Tŉ���#������]�J��� q��?���]1؎�^�J�x-V��>��x��B$c��Y�LM�v�����u�ф�X�o)����"�������f�;�$+6��M@�����bMX���d"U������O�ů�2�������G%���~�	�	�lc�{��w:��n_��#����94<x�F��|H���;������q
rK\s�<��eE�H�z�$ �j��� ��z�֘y�a��e�.	^����[��93;֡��Y/�bp�a���ދ��_��u=�֠��F��_cC����������,�����k�4ꀏ<+�Z�#j�>8w�ըI�M�d��������-�����)�OF��3!���g���qWġ���#�K䲍�qL�$U��ՋG�	eT�t1����=�͎���]��h���G:��<E^��E��4��r.����.�r
X�h:� KtY�,�&	�{#�Z�'H\�Ǥ��[ͫK�X�������-����?�4�}-z���v�R�Q�������N�� k֙z����ٰ ��͌�С�mD,E������#S���DQ�В8��ǯj@��C�b���sۦ��%X8	g��9sz�g����խ%m��7k�M��T��J2�"_��#��ضCحg�O��!B��?�q$'�jIŽ5�[?�h�@m��D�#��݂�U*����N������D�k&f���C�#��ld�G�Q����6���Bs�+���2�_�]��=n5c�2��j	�2˸�:z
��F�cޢ]� ��ߵҽ� A����R�d*�E^ei��D;��g�e�pl+� �-;���L��ԁ�\2?C>`P���*�3����[y�i���HȊGO!��7㆟�8]��<6�4�Er6�����7��1U`6���E�"��FQ,Rx�]X���k�(%���9K��D�n�U��#f��a�U����O+�x�Jd�s?ꤚ��U����V���?J����y�݆�eU�99S���Փ%�|��*p�(�}<�]�hi��U	 ��J�8��S����N�Ak@�ĸ����yx�����8���O� �r�jc_	D�W''R��'�awؐZ�r8"}������]v�q������h!bcV�q�ջV��Ϳ��j�"�`{C;�b�b;O5���}8�0�m؍�{�GT�yre��l �B;�s,j�7s^Ƣh�	�jҖd�T����흌t
����e�q��F5h��r���O� ���C!S�KZ�R�(�[���)n��Wv���"�eT�%)6���ڧ��ta�׶�4��O'g��W��F�/A���aUO���2�_�2qp4���(�M����+�	�!�Z�LZ>V�]����[H<��(H���%�Ŏ��dZj�ܼ�.t��2}���&��R譢<� BW`��/�� �����qm89� +�9Pٙ[
]�������6KC��(��Z��l��z�*�S��.zՊ��r�����5A: 6�}�j ��5�� ��V��=(f&}bή�X@P@��������h���!:�9M�H���>�e���?��1"��đ.��{ݍ���1a"8�:�1b`�jF��E<�5��S ;]��W�}�
�ms�^��u�V]������"@P!�ǼV�׵��p���q'M�%�5�F����]��dqm���zJvQ,�eY\^��!ٲ�����c�ŭ^u�6R�e�3-^+�b�K֍wR�H��E���}�Ѯ�^[QRx=�y�2;7�I���+'�I�),�D�r�f�,�pU8�������C@a�?v�EV!�b�f���k�?E٘ٮ;� KY�L�kT�Z���
C�7��������5#|L���,�.8��j��r�Z	e�5ɾm�DL�����+OKz���1�מI��Y�|Zc�N��6
Z ~B�$����9Q}>Y7#⚑���n�qFY`�i�|�����$�P��-�ftD�릹Y��%MgG4�(X;�\��,��%3X�����*�ʷ`�%��b��;@)�	��K�HX�����m�8�4]�[�U� �w��W���_�������ڻ$��>���<����τ4I�S��t׌�\���}�pؙĚjDt�1��������`Q�1d�%s��YmQ �B(�l�Z��Bʳ��ߨ"耾�vV��>@3.)e�ni�Q�C-՛ѫC��t��(h�WtY���AINi���R�8�p�#���~Q����.�/Y��=�rQ�/�	\�|�ԓ1�J���A,����,�fF�i�6%B\DҚ��ZE���+3؛��D^�c���.T8Bdk%\�߄�u�:&�@}? K#h��d!&6@�$O�ʊ*��68��~e��*�����䂶���b�MH��-$����7���H^CDgUku���}���-�!͛L7:���H���=���qLt��[C��\a��)Н�O��|q*��� ��f���k+P�3j��T�ζB���v�� <���a��u��>ڵ+P���x���qQ��+��%���u��o�;�I*��b�-���v~Rƪ嫹�;FE��ӬN����g�BvC^��ɝU���Qg�s���u�
t\Y�懑���E���$�!�+�G,3w[�D"๦
�~�NŵW�{�A�l�=����[�E���'~���شBGx6:���P�aӭ�=���Ҵ!ϕ�)ҳFv=�3�ߤwv��|�=π(KPf[���˝�B���E��!S��v`��)�V�nxk��G�Y^&��2|����o�J4u�S�fՍ��͆�)�`|��&m������O�����UfR^��e"�U f��ܵf�Z�a0��^� ]c�Uȴ4�oe&����|㪄_Wf�+��pG95�Ր@e�U)5�4�e35��5����R�M�1P��mZ}�L���f�J��h'�DT���u��vz��j	�t;��C#N�F�5>*|�(���z�Ӱ��:�)�"�Ƀ����٘���-�I�;�\W3�hd�tUX�-�V3�D��\���($A��T�+?VGꞐv��ve���&ǎ�'�1�j�U��X����1}:����Χ�
���S���.G\+W��u?U���t���d��v,��A�B�{�`���T�r�2	�����3_�����8���%vUw��L��,Z�x�5v�v���?���[I R6G� �H�M�o�I�$����2Fr7 ���%X����"�,����p��[(ѡԣe�oTDߒ ��z�p4EbJm������D@���(o��p��D-�J}�ٲ�M�����C;�����L���;����Fp�_z6�9�fJT+�(��؅��ְ��B�]d�_��N���"��>�W�e6ӰR�z��v���zC�z��ȞUX�$e�������tV%�H��XV�'�[w<�H�/K �u%f� mX�C_�뱿���>��}�����(��tP���y	�}�`4�X D�z���)4��Zv�ˇ����I��Knb������*�PI� 
�I'u�O;��ɿ�	�ۜ��m}�����M�Z�$I�V���lWD�:']1#{�5���x��*�cId�tmYJ�c?2�*����gT�ޡ/�4tI^V�q��B�aq�+�qp9^�u��u�}?5�Q����7���-�/e�����,-Q$�3w.O"�-%Y;1H�����"�G(�� c�|�E�-l��x��2���F���PMn�ӵ������z����Ƙ���~��?3/�o<�*�j�ͺ4荣�dY��ޮ覅o5��7�����}�{j�$��d �#<�@�>�f�`2d=D	��#NF3�yUh�����e�/ӗ��e�����=6��;-��o�Y`l�L�X?���KuG��ѻ �MuO��Nm��@�F7����.�d'񡄈ɖ�"HÙlI�S��N�F~�zD#a8$�������d�	Rr%�]���j.����VK�_W�y�Z�ak4����R��M��m�V�B���L�Y�[�_�N>;۫���Z��L���<V��(�3�Zt��{a�R�h���eGt]f֬���	i<(�c��0hn��(LR��=�[����U漃s�x��RX��\/ZZ��85�r�p�Wb��9y�O�ʄE����|�mt�������D!(�.��'������ �T�X��+E��l�ѐ�:�h_�,�A�������YZ��.�0���1� ��~~�e�]���b�yʖ�����X#8�r��D�;��j�vH^�*;rStI�<@�!�[S'0T�Zy�Vo;��ЇŖ0���0��y=j2�x���
�X��VF�oD���/�ｹ{�'
W
_EB�G�y��ưfY�`�s/x
e�x���Ò���7��¿�qUSa�j�p�c�~��$:0#�*�ޱL�A^Z��L��7�C�(Dd&�A�C�AO0p����f/I{��g0!���Q/����W�di"����j��N���2��̮咰i���5���ˊnx���md��a,>�ip���W2���y����3u��J���=�@��p��^�3�U���W���Q�m���Yǚ��@B�"�O�IW1n�����S��cO�7�|Y�,3���Ruy�A@1�����"\(�Ə9q�;�~��$���EK��M�z����1[y���� �Ox�wtlP҉dX��m?x~̓��+����'�
M���W%UX�щ`���~+M�4p>�~��
!N|��:��R�`��d�����lksl<c�.*��wX�F&�6`��Uh���W�xہ����1�%r�O�� 7�pO��V�p�dhW�Y3�&$��������=�0���<^��y�|g4��њ؋��Kf�6L��}��Ͼ���3r@��%|.}�6���t��י��#;Ĭ�ZD�k'T�e����<���