��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�d!z��� �vD�����?�gIp7��P 8���%)=:ϣddǝj����.�����{�`o0A�~�L&�{����`��6e:���W��ӥ����5/M�^��+ϵ��^��%^�F�6*v�����u*���b��`d��-l�Ņ��M�?���n��۔��z���;�������rl��׭���G�e�#�.�xx/��،���Ԝ�qқ_����8S8�A��<���T�Hw�>�ũ����p��x�i�<0�����J�:G�8�4��^�	������t0�@���Y��(���B��	䎒�\Q��OF�űC�/��닁�|]��%2�VCp'2�./C�`����M��x���y���437���H��'��nE�T���c��!�b<D��r������ϗ��C��=����v�7'(���,'i 
ȯ�� ei��V˼�4�z$� J�#/C�a���YNfb袵�v�OtJJ���%�GKgD[G�/Dm��Xf���=�4*k�Ќ�*5���1XV�K��R�_��\ʧy�V�oi���IK����V
&,�Z��uYy׬�Ź�wiG5�d>Ѽ�&H�CW�����Eu�����N3&�65MB�!�_1�,�U(��R<#%Orva��V��̵�� N^h1@tšt4o�Ed�J��wu��+D������Lq�A��9�^S�R��U�����$@�@4J��d�o,��^�`��Ϸ����n�P��M��訧q�q",5K����6)7d_�m��R�GU���VlSD�����Q5hĕ�J�8��� ��i4�dps����µC��!6�����E`DVOv�i�7��,�����/cS�\� Z�C:�n:Mt%�<�� !�vE(��l4�}�H��HZ��l�G7���wZ�"�z��WU
���J�?R}3�>\>�G���Ѯ�xBLӍ⃂�rE����#�K3}a;2*��x�-ޚ/Oc3TG�ۂ]Ӭ�s=t�j)��V�X���|�(�,滔.�ˎO]����)U����i�}ဋ�ꓻ�;�U�y����%��D���K�\Il����,wa	6Xy�MJ/�_����Q�n�  ��K�����JB��ˡ���H���$����\�-�͞O��A���rr�\���f�A��S�r&���kU����B��0����Z�j�+�@���&�0@/PC>P�>Z�D��'�Ҋ�4�jQ��&G�x>B��}����A������2VUV�h�ŵ/��ʾ����3M����*��'�� ��}ԣ�����Y������ ��J��J��� _zi���Vz�f)"�s�>�~������wc��H��K���l2))[�Զps�b<�أ-a��ދ_�G��r�b��KJV�u�"w�ʌ'�j��!��iy���� ���<:j�!�<!Yd����f[��z���z�3V���������q���sރ������=�Ț�t��*G��da��Ũg�`�� ���EKf����`��� �����cZ&���������Kס+ڢ��s`ڍ.��A-S"�F2��ϳ�ɪ.�uڕ�WwFTq�*���Jh�w�M-�t��b�j�X����X����U��9�0PDa_�!���~F�;y5/c7���ZcK���aV_���Pw�x�/Τ�xb�"-�U��<*m �]�\��Nṅ��P�)'{B�u�#ǬhJ��8��A ��@v��a����z�&{�S��eWs,���QW�@Qej�FP�l��l����tPH���̴r�c8�m2a7:��쵬"�݉t�S�h�yvuq�����Ă�W4bX9Q2�'*�e��B�
n�]da��s���*�L?�Gd����dDZB
�f�L�I�e�"je�����H\~���,�__���^{���K)ޞqF�>:�ik\��e��]8Pi�S��tR�rhZ4�"X�~a
�ٓAB��o�%n�NF���� ���2�+�A��2�÷1�����t�SF��yV~+Z
.��q� ����,5	׶�kY��?���a{4z|4�1f1�a��Py��U3�����(^ڲ80���<	��ݰo^W�S�D����"n����,!� �|��:�>D���� ���ktI1�:�vEk�_l�{�&���c����;�P�u��&Z�;$B�r�1ӻ�t�՘x���ʍ�}�����<���v{����{e���u�t�ȴQ�WE+�V�)�8`F�
L{B�h�g m�O4e��cJ{��U��j���S닥�y�~0%�)���Ck8{�ب٪[GT%�/z��`�TƠ�%OM�l�qXq+k�G����N0�=S�g�x=IޓA1M]2���p'�U[+�id�M�\�w�C�bOk䄟� RN�(/��C�ě!i��Q��"�<l���Z����v$
��
��ɝ��/5��H�GJc�?�xb8s�לn�8H���=�Fs��{E�`L�/b���:do@���,�.�s̔�'ic�>00Bܱ	�=�uVk�������KSFq�|���ЂO��V�~�O��1M�.��nd��޶H��k[�
m��B�g��R��2��Ei ���M��;�R���PpYG=ޥ��[�0z=�Ao����� Z��j�4�P\�b�3G� ث���v/<�[�H�R"\���{�	�6�x���_���}�a��A}+��G��Q�e�?HnU��>j<FK�V�#�DȘ�Ǜ�u��{.K�~2� l�xm�.U�W���~Ro E��C���I�����S�,�3�O���_�Er�P�W��o�M|�p�hf/7h	J8�I��}Fn�-�X�\���%%���Z�W�c���lX�뱿Β������D�0V��y�]��2�Bb2R3�����o�$:c�	"�r#l�I�d~���I-�GL���d�\��\W��L:��؎�zx������䈄�:J��5t���$��?���مX~*�z���tN�<:+�S�k��ܙ�@)��y��;�ڡ���)uGu�Ƣ��1�
W���]l�_�H���SW����B��S�н�Z���ߣZ�X�7���껵�K��Qt$�o�͜&��}��w�:�Y��wj0��.���df��~���'�̛,�����`̚��������6U�	�1M:���uF�����4󖼼z׻@�1\:gq/�J|�GN2p��,���IĪ�X�&���pş�+����Ϻ��c�a����?�y<��Ջ|R�:gm/�=�u[�"��P���^���|�TΪ���g�F% �l�hY,��6?;Z�;ݏ���W���X�&�H���g�cJ7bK��N*�Lq��?Y�=tM�D��"�U��uMԭ%�x�Ϊ��^?�#��,^�1m$G�6CDPN��6g�rF�5x|�rŮ�<d�f4��Ի��k�xÓ��j�u[��_��k����.c���.=���s��>�߈ù^�>l�����?�,���`0Y�N���꜖D �M
�/P&�0P������p��KTX5!���'p�:%��VF�_�i�N�N$<�J7aj�	��b�sY!�J�����F�0Ǎ$�VJg>�q���m�23��;�K������c��ȶ�6�����!X�[�2���ƺRTwf���da�����V>{C�<�R��?G#&�06����ۥ����/� ��$��,�q[����~v�C�#(�m���]S���D���R�	;�8�Yc\b��Njy@��}�Â�Q�w��g�8,����G|�ܦWt	{l{�\�Ӣ�r�˱��U�EܠM�^�p0!o��o$�+�WPEQ޲�x����WZ�i�:�s}���.�Y�6�wP7A/�D�J��7 �+���=��QK���Bc�3��%���N�JYn�\�X�^�E�����d��J�:ώ���ű�w�<Vǋ��s�\q��\��^��*'��)�A�c�6ZL����˦C��?aS5�"Š�;�����4Mum}��
�c���o�;.��@��U	w+�@�K[<�F��y�+V�t�� u�r.���ܣ����1��@r�_jI�������m4�,�, g��"mN]���$����ջa;�l6j��r�)��b�S+�Ԝ�������*�T�]W����T2cd9���y\`y�bI�.���3�n�Z?���ZL�e#_��'�W��&�f��U
um��aŰ�*��j%Yς�q����~]�ɳMX�y�O�=[�T�$�y껺0W���gn��|d3��0C�s'pյ��6h1_�imo�i�ŭT0�Y���$�+�kZ��=^JD�l��(�.|Pd�P���������@�.��s$�
lC�p�K�]4�d�hs�8�Emu�����|)(i$�����pxF;������n��'�
lDc��iJQ��d��/6�y:���-Z �2Ǵ�aЖ0h��#����GJ��L�E���әi�	�����E��I!���&4��f�Ֆ�i,�KZ�w���~�
���@�����=��"����iE�3W�U(?ٺSa�$ �=�(D!hSm���� ����O�$ׅ���
n�9X���F�ua�9|��,uŲ�	���G�<L�m�(����,�f!�Ewb���h��"����=�������g�?R1\hA�����r��1`�n�X��2I�`����N�� Ga�}�V��i��M8�h:�-���$BPsopJ�_F"�/��{�|p���&Ù��`���ƍ��Z�f�l >�^��T�����b��ky}���:��2����֭��Ȱ�-����|�b�Z�l�Rs�B_sӐ�QY}.���=�W��@𸪎c�½���]��I�&OE6_�᯼�B�9&L�\a��ظg�q0�!�w"J��v�尶��_�A�T��܉�!��B��x-�2Y���� 
���o����N��ꯖ�����tQ�x@=�Q�K��@ӷǇ��t�.?y�@jcB'��@Μ�{�Wگ���cZ�b�>`�>�=j[�F��D'mTm���j�;�$9[�ʕ7�ޟر�OAE��!��i�w	6����޻��.v?���i�q�V�	rMF���.����`RY��%$J.��CT>_��e��;����c�zq��L1�U�8H7&>VJ���5#�����	��� iyh�5���/���ٔ[�X]O�:��!˽���µP^DdE��O$���slj�Q.L���Ӛ��:u?�һ����#