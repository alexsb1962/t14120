��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&�����6u��%�R�l���ɒ�[������ e��4t{O*&�z"iM���z�� _��)X;�g�(������<W�;1�g� ĄY�;�MI�u\�Ĥ�P�њ��P�8��ڙzd��<�<�\(�*wfn2N�
�{QG��I��"��6G���ꪗ��� ������M�`��_�5ThZ.�8,��ND����X�Y�Z��p�c�U�q����
���z���а*{��Z=Q�?%y��aDIp�M�:��^�*>[�ǯ�r��a�IUIW�u�w�[W�c�]у��FDG��ܾWm�􄗐���O}PĜ��(ӄ�r��k�	�;�n-��>�Ƀ(�ԞМ��!*��й4�e�U�ܷPM���	��Y�pA᤭��GQ�E����յp0���?d��t��p$���Bx��tk����n6��H�(�(�:��)�n��H��%��������h�:��h�X5T~%����HH�����4���=D<���n��2ʾf���ġ2���<q��f��2<��a"�R,+�V�|.�qHޢv�Y�C���H�C��@R��hDۦ�#ۡ�����:>�i�E�K�:�v�gmY������M,5�I[�w�im[ Z�mg��8g���~y�G��x|uJ_���2:����'k�����y���$m�����Зkj��{�iT�M��M�b�b�;>,HM�X�Tѿv�bt����}㽩m��,���*�6eď�>B�8l��Sl�jr	�I'7�*9�gT�c�a��b�D�e�u�9��=[h%%i����ʘ��`;d�	�������
��R���H�S?�����%Z���b��؏��I��]{�߂��ow'����M�$-��&q�~��V#A��.���>l���g}�bg�F,���$jh�Ч�L�*�Gќ�8��`��G�ٷjS�Msş�:��9��S�4D2i�M�b^ȴ(�c��k���_�O.�8���>uJ��B�xwy"xe3�[�s�y�g1(%_���a�Xk5���X��ţ	�vj��%è�$��ca�z0�����]�q�0�oe�J��ʉg�#&�gZ��h����h�Γ��2�q��y�r8-ܺ#	��Z_��[=���De����ȬA���k��'u�@��k9ϖ-NI���)�UMX<�`��P�;v1�ߎ8��;��:Q����ꏪG��C�c��*v��t84��O���ZěQ.��C>5,��W�]����?��Ӟ+,� �īB8��6�T�LXl���QHʓaM^��C:p�˔\���`Ws"z\����g��Ţkg<xZ|܋���2I�m�V����*9-�(��"�n�y���!C��y?�eV�W�!sO>�7@�s��ÆJ&q�(�4~fP�팖�Z<��?��x�G�c�d��]���T@�jS
yI�Pr*����4�JCNt������E�rA8/�fV%��$��<k���GV�y�~��6߆H�X�Q��2����:�����$�S����M��I�<܄�5�}�t�1���5���� rf�?%��&�`��is+Ʋ��z�$i~
�H�4���>�t�z�|���p��ihD?\�K�D��{�{����p7�,?YYv�ԮT���چF�6�(���𹄯�H?�&u˺��]�MG%�}Y�Ƿ� �~�����½ͭ��(��0l%^X���wW=�~�1���Q!)�J�-����/7�J~�n.�ƥ�`th�n�����-D�!\��e����X!D�Tw��r`�h'mW�����|�:Ny�m،�3�+p�����W��Y�Z���ur�LD�G������A����w+wZ���qhu�z����Q(���s��dUƊ��c,�6i����#*6���m9����t��;�O`&Q��ܺ���>�������j˓��_��yʖ�9j����i�61�i��m�z�00�mO�,��oy!O�=�\�ݬ�R��X]������B�|���^ 8��	�K3u��|LS5�F�5�]�ۿ4C�'��[�W�^ii���j�ʑ)4�o1Eh����i�FXJ�>u���|7u�s�0�N�K`�yjd�*���5:�}C��9ؿ)�ֹ�	�ަ����R�Fȩ[�Wω����5��%�R˃���&�c�C48Z�����*�w�O�t�cX��N~�x�*r~@�i��:�0Y
�Q�7�iXjƑ���q���}<dV��z����<���3��A�[�~��h+�	�r�obZ���o�7��\�� �	*Pɩ��Q¤b��3r_[��%�#�<�ɰ�&�ȗh���zق��1���cL�dQ8y&a9s�%�2? E��Q���A�J�U�a;p�R���7�$
�g�Ը��:�YG�����C�/�q��S�����'�SS�Bwf�3q��;�@7�˶�,��ݟ����X�qxd�R~֚��[�ރF&"�ԅ�Ƹ�sH���KUI�j$���7q������!Wp
�q�|���s�uJ{���3���b�[�!��>-��o��<zN��px3S�.w ��8	Ӓ�{�_T�r��<L�%��3R]nXf�N�n<������K�E�(�Qg�E-�D�ߞ�����Df�ŉ|^Ҿ@qf)xR����q8����X6���k���/_w�~3P���	j�����wz_������K��T�`f
	�A��
~�
�\�`�y/���L��a�GX�V%IJ��pw�b�x�Č����`��v��>g��?؈��D��Z�_�ˢ����V��y������uN�.�
��I -^�oOJ�e}�X��Lx�9�V5�9cC������8�5Ps�v>/�RC� x��Ƀ������u��>�
h�������&C��7��¾���F�Yw�byb&e���yf�4���-`���5�c��H�ay=NU�1�X
�'��!���;U{��Fv�����M����F��k$�%�jj:���ft�_ZA��qYԶQ�=?�c�>�p�;�w���"��Z�< 7��H��� �aՂGk�b�kg��S���-^S +?��v��%�[ZD�␎��_���D&S*�����(�����q+#���q7�A/J�H,V� 7	�����h>#|(��ªı�����D�ifW� ��)u[@�7���@X1��ebQ{��\Ue��D���5,���e��N� ��F�Y6 ?��7���+4�!X��
�-��&�YLB��>�w�F�5���h忕�\K;�Wާ��a���h�&C�p7�e�~̕��hS�%Q��#�rd9�ӈN�IXђ5T�NF�����N|�LI����!��] #w/I��LwZ���z�i�g�ٷ'S,Vg�o�a��;"&M�?���E���b�M��T��jO�?vsM!+KYXT7r�k#N2*U�U���ݭ�!�K�	��#ҙ�6燴@��s���6��H��9c�L�(\���f)4�;	=g�i�H���ŭ���3X����5C�%�E��3VB���e;�޲�v�"�)�Ӑy�F�&�7x���4���gY[Ԫ'�`��֕��1�+��Op�e�=�Q��$���X�$k�_Q�Np��G�����3���C����Y�"Z]��Z�uG�'�^Yz��T�x��|?�[d�
qk;nⳬ{�X;8�ۣ`�Q��6���z0��Dd)z�G�n3�dK%�lh�B7=��E��$��q=?�&-H�S�Mo�������VI˶����:��Ky�����F̫�&����ν�xvn!��ȏ��U��7֎��E�z��ֻ���9k� �O�_-}�1�_�z�Ӹ`�<����$A�#���0r�[N�肬$k<�S�Q���K��k��Fg��	�6��ń�����V�/���=�O��z-	�9)x��缟敂mG�jJ�D�����:p52�������X;���b�"�I��7�:�����m+�!|�	���g+!�Њ��(����x���bk��s��q�23uۏ�m�%���Xֺ 	����]ψ�d�=)�fMz3-@����0R�M�+����r���3��l}��-߱'}���p��C�S��C��.�A�xP�+�E�n�{�m_S����/"�DV`^�.�z�ٯ�R�y�i3,��+&TR��f��K*ce{�I -���w�+޺�b�uv���@dt���f��ً#Z����+��:�.�)YD���� �K`��X�',��:�?A B�E�O��t��\?hY���g���P(��d�Q |��%�Q7����3=���!���xLP..v]�A�yŽ=�SO��2�:�dG��؊�2Y[�0걘�Q�ˏ�w�,
�֏�9B M��˾�u|� �0¦.k������u	�Z�CD����S�)�j�V�#>
㑩�ޓY�>/�{0�A�5h�>���WKF
��A���b�a���O��ڦЛb�:���  2��V"wtĸ �e5������\����4��(���TytId���ݕ��(�ʸX�xeG��S
O��yX~}=־!�P��?fV�Uut�'�I�$���"btG`#�q��~kP?2���bu	���M�~-��� �n�= �vr�l?����a�+?����&a=�ψ�ߕW�h�g!x7��˜ũc_6���̗{g\������e���b �㑛 ي��sĂ������2�쿟�;�0c�ޥ�M.���ܖ~Q>���I�˱o����3��1sa qQ�'��n-�T(�?ɍ�җ%'{o����e�?�u�!/ԎG�*4��G]�8�W��,[�Y������T}Qk�� 
u�h�|L�\�:�)u��UR�-�]$�s�]�������e
*�%E���=y9��fI�1͌L`q-������8(���ӿŰc=S1OZ�4�)�����c����&��bE�)�ގ������� ��>��!��I��y�%�Z��BZ�C7�dA �U*�-ɤ0g&��U�7���m͐��R��`�^�ԎE������A6����2��'��1�JZ������,�^�sA��3��D�hG���G{׍��WN�5�BH�~Z�Ks��\�!�1L*�(]`�k��\o}��e�0��o_F��z��;D�i�B�0�@�@ \^����J�+�;�l��c�'���޹o*,�\��һ�LĠ�4����^(fR}��|�q����&��P1zzL����fA��E��|�~ �U6S���U�J�+��F휮���"���B�O�nؿ�����"Q|ɴq�H�}�P�O�ߑo�aU�F�����n�e%r����МdL�-/�2�v8���S�y8�|1?n�h��	�jp:U�)0H~9�AQ�o���N�C�4*�X��	�i6ވ����� �.
�ߝ��{%v��9�u�$U�6����/%�@���X��Oe�#e-־6���\��=	����I�Y
�.��{��W'Q9;�����L>��̏v��;$PGC
:�v潁A'@Ho�9�yW� �H�`{
zd��y��Pt�+b�Hj��0�'�saiz���@���RV���,��h���z]�g�Ϛ�2,?+`����P���A��t��s�l��G��L,zL���0��7.���ۢ�[�X����0X@+����kg��kQ ��!�����.��i�]%�|ܯ`u���p��'�˰�`�Q���q$���ڄ�(�%=N]�s`;�4.�N�#���iv���>c�TT�`f��QU��Z���k�j���cF*Bs��ԙΡ�������YM5�m��s��}F�f^ ��S#�l(V�u#�6��¬iv!v��,c�K|�����J�� �{�?|	���5���'%��!���ܢ��3\��"���b3h��!�����M����U�2���( �]SP�L���/"�yZK<�CV��EA�Yp]T<�c9v����_����Nް�M���aH��	�KN�ϛ�.U�I�g����Q������I�GK��q���PTT�I"���rc}׉��Ki�������EW���	�k�Q���4]
b��a�&�¦� ͔�S���9��3���Xr�D��-(���.�6��6s�X������@}���3p�WAP] X���%�T������ ��SQ�Z�#����g|g����x���?�M/�=����8wGԷq�X�K�	6{(��8ޤ� �߉4�����_��H`"1ߑ��kn/���*k��n�6٣�t�[�8�d��3�(C	c���:JR0x�V�jd��f��c�*u����s�)�_�敺�@h��駷=���_�b��e�O8|�=C~����A��}x_w��҄��M�Jݤ(cdD���+�]e9o�M�k��6o�a��X�:��L'_.���;o��%�-�PF���E�
W���ڕ�+����l4�g�W罿�n����<#U鵬�ի�V�l&�=g�C-n��Ue��^<x�lP k�S�\�ϤK	�G�8�W��6n�}�W4�l�Hr9�G�����/�����ꧩ���3bS:����`��82�V�����C�nW�U��|z6���:�>4��Q6��
+��f�iZ ��j��~$�;��rN�@^&���]S����=��s�f���Ӱ"�3#[Ձ`���Yu5˖G�Y�����c� ��h휯�L~t{��A�s1'
��J7���J�c�:06���o�L�Ϝ�*�CY���|�l@�Lf��EW� �f#]��Řie�)�I��X yv0�r�\]Bʷ��Q�����g�U��]�g���7�� ^06����	�~5X�?��.i䊎Ô?�m�s �����������H�><,O.�K����?���<I/Z�  !a�0��O��e�K��5�+,��f{�0C#�e�(�F=�XAz�,�Q�]+�Xb��_�Ŕ'r�E5���]�>�4�#�(ҏ�z!o�OcڋR�
I��k'�H���=� �V��nv+V/"�¢�Q;Rw����!���oҺyYY�P�5�c��@ւ�r�J��-:��u��l��[t��?�>��MGQ���M��E�t��D����jh�_<8>tX�(��K�=h��8������S�x��dq0�p����ͺ���{��`�ǵ՜�v֗�(X��7���e��@M�pj\�J�<%
�$ԙ
dW�s�EGz1��`�&C�������F��F�`��,� dւ�?{����9?Ȧ5�8�D�����.���$:��g�,��Q�0�Wq�wq1A�/�d�������_=��C@�fTc��r�7��@�s0R�&m919���<�'2d��ǰǶ!7�ʏ^���!��t�G��O�d�y�o_���y�An����P����6.��`i[r�OB�������������OҙP�J�s7�����wBP��,��F`�9�c��/�<A��3SUॣ���m�������xɋ�'���;z���V���ˏ_�z*�3����D
��̛u�N��.��j�}m�b�f��'��p�V'��{��BMr`Y�П���9���">� �ƪ=Da�NN�s���Μ�d"L����Y v���rD��?�QeG�ۡ�6b�5ge�\����H�H� b�g��|_u~󇷒,�p�z�� :@(ؚaT��x�ҕ�5�����AWU�8��^�B��r�k����F�vc?�*g�oe�;%5�b��ւ��q5���L��n��'�7V���D����=��e����Ap�Nk����p5C��?rK�=�𡝉V�N0;���y�4O�hH�}Ww�^���]�IG�
����[��ak?��iRj�J-�CT!���-;f��{����F�Kj�Vz*l:Uk����c,�и}q�"�X	]���4���M�����{��"�<���y��8*?@�ژEKJ--fr泦�.�Ԋrx��µ�Cn�ǽ��t��迓�u��!����y�G��q8(&�'�Tg����Ƙ�%g$?6E}l����4����)ܟc�t1���P�Uzauc,��2M��y�ڇ�1ҕ���8t_F��6�"�vQ=H��g_a"-�P�^�q����P�\�]T����^,>z�x;�x��ԓ�A�:TnCM��y.�� ������m7hv�����  薯x^�d���{��W���'_�/�lx��XoAz}�����\�нƳBZ�>ؑ�:��(���9b�8X��;�5��N�P��.g�*f���b$4ٻ=}�<-��5����=�k�;1�
L͊�D;��u�@o�@-�a]W��>ĴR��b=7��$��P�+�"^����NÕr�CD?�6ۦ]�_6�h���@2��?l_3h�e���r)������rW0���a#X��f��^�sy��v���ğ	 ��-�H��Ћ�U(DEI�0�QB9�m@��p��m�l������{��rH�d���cٳo�Q#Z!w��K�Z�ݎ�4C����l�1 Fy�+��7�G�dlO�o�1s=���U�R
GcU�7�$��=$
�� ��HGh|�D���8-o&�t620�Nc'��!�R�H�:���*���QO#
���|Ud�.�v�L��]�����+�N�O�f��� %��M}�in��v����0�n���2@M`�.J��W�f�ϮDLEA����򌝭�������Px*�ItO2�)��<%)C�^�7�T��'{��hS�1%������{-�/�T�,�=�y{E�ؒ��	�$���bS<��)QnjF�Q|�/�c����0x���ԡ��-OF�U�	+���}p������f�t�b�*Q��z�uK�dw%vVه�8�JR�`y�铍@���]�������PL��e^H�@W���-#F��2�%.�%?��F��_w,���$���G��z}:X{O(�G��ꦉe<�ǆ���?��x �}��0�V��ؤ�g��t=!R�mf˔����5Q�@����?):N+�7��.A�=��rWȼ[��p�3�����M�{�.��$V��99>���$b�M�ޤ�l8y�N �S>Xu�6FkX�_�j�֌�,�<�;��	����٢|s$W�>�`f�Ğ'Ғ����&��
@F�ԈD�PJ�Af�J�W�.�=�����"M�0��j.O�{����񶟢����bmΤiP�S�}-&�R�'&��mbZ��=�*�]��Y��"��g	)�ty����ޅ{�<�	g��+94����EXmj]x���^D �{xHp����u������IѬ��'�e�Vqs�BQs�zU��3���:d𙷍�W�	������!�ݺM���!Tн������/�8��^�qߠ�w��"��U�_eJ�ހ�f�i}�T�&a�@�z�G��b��-����<�[LDYr}e��a͉"P9yDڕg^�=5g��>�b�Yz¡��j�]���mJ.7�PY`	�� ���ɫb�틩�[�]��i�%��Tו3�����SqƗ$a�y
�{��xM�ֽdh�;YHg���.0�o%~83's�g{:ab{|��v�`.��׋]���y��[@� �=9�	�.2���%����*Q�f5��&Iu�n�
pŧ����)���6f#��Bl-<	]�m�{|`5q5�Ъv�կy��FAs(dN�3�b��(�ښ�U[P�aH �c��ʨ'gT<7��j4��^��c�x� k����^M���SݟS���7�0Y~�w&X��z�FN�סJ�X�O|��`D��9�^�h�	Υ���8�g�d�ZF���ԁ��*6�_�?c�
�e�UGE�ղ�Y������N�M=��'���מc�KQI�,5(�Q�����Q����U>ۧ-�<jհGt-����Ԭ�U�����=P��fT�L�o��`r�����z|���l;��H�6�����P,J��k��J,�nƀm�6��4,]��0P680��f�����<i������WM�v��<息�����еw��S�I��5�E�'.�d���d�Ήࢭ�a��r�?�"��7:%nD���~{C����T�����[/����rI�Jp�g*ut���|��	z�B��6��_kA�څWݳ�#�m\�vq;Y!#v�s/�,�	b� �Vf�����s3=��2��fQ��!���S�`^�g
, ݑ��D)?����f�4�N�q)T�B�vu�3��>|�����Nf'��\�7�Gܪ|�����|>�ߚ�&���1H:�IS�A�f�����C�k!�ظ Zo�<K�&��(��0 e"ڵ&˃w�,7�>6��㮞C�T7ͻ������d!O]N�Qj������Ջ#J��/��QD���E��q���Bw�e��a r��l��x���~�?^PCq$w�g�)Q>!'��F��T����6��c�As8&�]�gJp������v�M��Ưw�.�� ��U���m�K�HI�~�ѹm�>f�����+�F�g��u$�N��o%#�E6�>�}t��7�2�SL�W�(��|�q~w6>עn�83*N�*�g$Ӥ����t\�t1���-g5�t�w�l�`{U������e���(>���!��=��"�r���1����H��SH`�X���������Rr�9��7K��gG@Uɕ�V����̦;j�����|�4��8ұ����K�6U�UDv�n�VLʧ���e �	����`)G�Y���e��%�'¦9�2�cZ�Ŵ�7 ������%�/y&��v�i۲ho`xF�?���N�R_�UMs����e�J36`w�͆��L6��o�u�{Y�7-���9D7��"�O����N�|}V� �L�/1����I����b?���b3S����,�0���$�#��S����RܨL�z ��d`�E�,�5 �N����vT��Q�����]����!��H\F	����5��N��{�!mj��T�ꈽd !��#���4�ˏ�'8�-����QI��R�x"�˼��Ȝ~͐�ЁzΈ_n�'҉�VI߆N���uˁ=)0��Q2I�mEǕ[�
�� a2��J`1��,�5�3�Hٜ�l�"�!��^B@���B]��px`�23	��1oݠ�5�u0��{�Sx��߯o�b��.�앁�U�����9�G�R��X�lLwk6�cN�5@~3	����-�hߗ��c�f&.!�p�7"YJ�f��QBs*��d�S�[���mU�W �]9�z��UOܾ�g�A$E9�Lp��o(���r�.�cQ	��w�1���
?��%� ��Y��%���1�6>Z�n����2�1z���L������
DVd+�W�*���
�d*�~d�ŋ���QW�'�Wp }�F^��V�b�u�]�|b���L��_u��A���(���X����TX��l˯Z����a�e�����K@��s�%g�tZc��I�8�L�F.y(Ș����ŋ��8<}֯�����x5V�?|O4bvzɒ�J�de3p{�-��c֤�
ܪr4I"��(���v@*T����(>'�����=�=U���N%�5���|>O��]>��LW�7G���=�M�<���]��0�	�K��e���P�zz�@��<����"�����������蝭��z8����f��G�����$��r�)0�:�{71�����t��Aۙ�cH�[�V/��"S�[���.�*`u:�ـ�j03s�b���@L���fB�������*�|��k�P���H��w��y�(�H�0k���n�7�j+����z�ﾻs;�M\�嘔t���5E��k�FE��k�n�8���0_�Z��di�|�	���&dtf����8�T1�E��}��巗~����	N*٫0c:��/2�R��Q��	*��@2e�'@$�bع]�#�q3d`�_:jʇ�z{�Q�2�ب�6Q.� wi��V�\|ν\h�˻܀�	3��L�~��SϦn!�Sl���D�zն�H��&@14�ň�w�Jx���sv3�ػ�xHb�C<g�;˨�u8�}����j ���
���������ɀto��޺�,Š6�쓢 l���@�E��-,���L^�]��� ��4������~m�P^Z*��0��U3&�.�"�zDg�oG�菨�${�{��yu��xq�w���"g�9�7�3�R�E��]����~yZk��2��x?%�La��#�Z
�Ęu*�ƿ0�lSa�o]5����,f~�H0}$R��9ś��`o#V�#�2#�3������`Vه�hL���`Yj@*ƛ�a��Zi�LVٕ��Nz�r3��Zd��㙙t�2閎Y��5M����q�WS�ۚ[C�&ţ4|ݨ��_�V�}#���m�<vPL���{��Y�+;ija�$��3��{0�>�PIdn9_|�z���N �}�ę�=Ϲ���ΨD�h�b���{ƫL~H Ex4h��E��[��S��b(�gb}���1���,��f�;u�@�?�3=P�q��f�`�@w�����ȍ<`��"T�2]�\D_�b�n���l�%9@������W4�%�Ah��8��뙥9'Oc�U܆���������3e�
P��$�^��3f�X�IH�Y��6��u`��H�Pw�X�1�AT�L A����A6�dϪ�Fs��k!~�q5�|�4�lZ~��MMJ馵���&�͑xc� dh�g@��:����b^Ը�o�=)~�HC��`��a	��mB�2�̃�h��j�(<�td>�p����z���&��v������Â~���N�n�`HG�U�,X�G�Q���
�Y-\,9�30���2l�I�kc�|_��\gW�d���H��� �A�~+	|5��� 植��aZ�2�)���]�:1Ҟa�|�������v�mQ����M� T����j���&�/e�?�l�A�-�]3�y��
���KM�~�;�? �H����\Æ��{��b��[�0��BD���f*`���pR>M;���
�����D'ۨ�{E�e�2Oɢ�m�Sm�Uk��¿c?���Z��s�?�S�m6x�-��a�d(�ͩg�陨��c��9?�?�3�֎�)�
� �u�=?���|�g�������kt"���\��z�h~����;�ڛ­��z�"w4G�TS9�v�uR>�
7 �4b�'���HS���R��U���> �Jס�M����{%3�}���$m Ѵ,��o4�zL��9yb�(h������H-*���y/;� +�6"�� �s�����<�1$�4��$U>"0*�8.G��ۇ���#�#�Ēi�w�l��
���|վ������TC�*�M�!���,�:���v?���a@}�!����&��LL�ɉOVcFV�'`���^%�^�Q]���UK����O�$cs��B�N l�T)u9�O�+?]r��(x騑�3�.x�ӭ&;�k��Jv;k�_����)�|)�g�M��2�6�E���U.�q�Cʍi�ُ+�;�,�-qz1�VoU(�v'�W�Ȑ�Elѩ��2܌nPEkM��ǰ�7Ѧ�ܼvI����!N\��誮RCeM�d^2s��x��ܢ^%�=���� v�G^u�-#N�ή�ud��i'�Io����6�������>����#���x��e"�i�{_�k��Ƣ*��F�
?l�0���΂������}Ք� ����*��9~Z���H��&���F=�r~Ve�_��������C�/R<5��L�a�MVC����Ό�A�4d�m��"��WC����Qˁ�(�kr��V�iw���6��s�߀x �ר�Ѽ�����w�5!#��) $�B���G�4�qN� |��Ч�`Bzw��?V��t���ws��)M�o������>�<����L�I�S
8��.�i0�֚��BT�R!�۩�<n����v�;9�`d	� ���|��0�N6���i��'��֣�Ü!�w��<���=� �G��D;�p�֍������Öf������vy$��͕�'�B��ڝ�Y��G��i��*��n���~������9~[�il���ϸl<��)�z�CG���P�[��b_��Z���RfZ�=#k��"e<P���>a�0f�;�R�@�E���j2癿�o��M�����cs8z�8֔''2 ��vyF되�>�h`M�7�z���	쮭���""�Z]}
�yb�3���P�=W�l�����#���a���B�3����p�g�dK ���VxM���4����!���[Pf�¸0�BjvA�����<��1h�N�ƺ�01�e�'�"���ڰī�� ��a��N�w=9�&݃���"Ī�N�L��]($�nJ�1Y�����(�J�G���)�R����v�(F{�O���9WN�ې~��=v���N��t�G��w�C���(J�डm����Peb	r�����lD�Ke�8�]��X�w��(�S��J$�M�U��]�Ř(�,�9,��G7�.�J[���RA�䋡�XhKr���f�NEK:=k��BG�O���.��{7�[U�'�c+���)V��;�O���n��Y�.ak9�261��G�u~���V�q��^=�GqWj5�b?AR������O�K�^=Ze�{s�ET�&E'�t��F��%KϹL�tN����q�F��h�2+k�<ükϘ(R��y���EʣUQRF-�;y�����H��A(Sd�)��r�N�U�ߖ�!q�~.�W@�=E�[���u�`ć1N���o���R��0ގ�%�,�5������fWX��c��I�^�+d��0y��|�NM