��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����~�m}:�)O��`:�5S�_��d�ߙ�$�#� w<����?�^� �S�Лv�"5K@Dz�������N!�A�u�����i.o����i�+a�|C`bW�s�i{p�3T��M�NlWZУ��B��ftDS��zq@P�ձ8h$�+}�}*�xX��JG��0ṷ������}�Xv(X�+Tr�,��^�
|5Dq�!F��@kN����2��ԉ�d=J���Hyz�o�B�8��oA����%�s�5Jk�a@���{��@��U.�^��j�h#|Ms�tE�I��t$��U��6��Y��-���k��Od1,r4�?
��n�͞��Zam���I�!�N�)���O�h���hU�$/VD{�~���"2����tv�0ͼu	�>K�^<�d�<�>�S�}w����Mt:y-G�]�S�͵�hz\4�hĸ���[�k��Ȼ�WC+�7n�nFAtQ�I���5��$�y����6�q]e��F��Gp�0�������RwѸ���ߎ�(�guv�X.}	�I�^d��d��ui��9�(Z�@>v%�!|Z����������i�[���H�9���}+ͺIaEG���%ZS8lՔ7�nx39��N_�a�[A3N���T\��X��$��x !��[�;9kT@�3��8y����y�J��㖇��+��o�;_3[����F�Z�gX��ͷ���EQu22e�-�o��1>@���� ��\.4�a.����m�J������L�����H��hŔ^���ᓇ��|�8�a�ۚ��%#S���n����5��+��:G��&�K��%�<��]5�Il<yK���2��~�@J �5��������>���5󾚚��fb<��q�i?Y1��3ii]������R�`���f+�әf�����4aU�Y����L��gp�g�I��K@Sj��ġ�C�i�����Zz�]\�y��_h�	'�ߍ�Q��#�L�騢����\��v�L|�0�D��v_��Hh��@>iy{�
��+����3x���8�O>)��(��s2��"�qP%��ؖi��Ebj���G�WM;ڷ>pyH�\%m�w�k*����~O7fg�K_Յ���fR�Ͽ>�˜eJ.�T�	�κ�W�풴� ��}���6x_T,JH�&�8�Y�/�
������X��F=�@�q���ׯ#]���o�Q��-Bp�Jۛf����8�JO���yH����2�R�Yp6$t%m�ќB�$6���O�qw	\��)�2X%��)�}¦��=�"��8�5]�1r��Z<��[ާ�xx�S����۹��kil� ���).ڄy��'__�߅�I��/~'eёN�BM�� <�ϧ�����nM{��]Kð��(�L*AA�  '��	z�϶
��i�8�k���oTffIoAb��U�noc(�SF�f�r\�/�&Aa����O a��)���<^;�?1�	9�14�ԝrd����EKӔ�F+�ש��N�K}�5�;�U��@c��^��oKM����Q�d��La��M�3-��Vd��^�
����=��0+*6Kp	e�U��>�7ҥ�Ǹ�#ʗ����xu��Ҵ	u�[
�X����Ѧ���Z�!:w�+T=5��7_Rn�I��på���"�3F��L��^�4�ȋS��r�:�{��|���v�B6%Q������JR���JQ5͓��_F�e>I���;@�&�*n�A�j�k~�[�<e��vl$")Gr���`8��(l]y��� 0��
�A���0���Rm���0p5�~���N�^:s�і�.Q\H^�A���Ip{��C�]h�%v�2L�H�eD�s�)�_��gT����m�58+*����{���9�e�E�
���>�1}2Q�� �s6�(����$�O��$qN���'���J���DUc�:�Q(�'y(�;d\������e�D�W��{Ζ���u������H��㏟�gX i=�¿�I{{�"7+�,߻:��D|K~�����h���Iŀ� }���l��#�S8<U�f.�A3-$�OG;.X�Ĕ��z1E��ӆ{�T��� tN�Yj]�*���i���r���
}u�U��/-gH-��"J��dO��S�2�k�������Ǘ��7��:O�π*
���y��\.�$���� �4[�d����6U/X��`�d:��h#������	�G��0L�{��׊����*f� !1��2��ct����*��i�
u*ي�'��$�
 !��f�y�k�o^پ�.bh�4&�V�3\t}U'c#y��\
i#l�
�HF�
��%����$�/eS�J+��=�?��ζy��i��H��̰���d1�� 5�A�e0�=.�x8C=�_t)pu5lzgK34T���v{�ȥ<N�j�IQIh��)dakV~(�=N6��ّ'{�Ҫ��0V�&��'�K�*���^������R��)��� ��(�+�&�N5���g��ŎR3ЦHeZ3?G���Q�Ʃ|·0��F�l1
����A6*6���� �Έ�౛k#�ɾ�D]ޅ?X���b�R�pB���Eؒ1<�d�p��Cϔ�'Eo�v$�b�r(����s��j�z3 �9�u���\����}���é�;e<G|\�1�=����O�����9�얂~�L4T��&5�t�A1� �=��^:Q!!@q�o�e6�E�m��[���$]�	�����1�®W�}���s8�75�	&�z�5$���8��a~@C�}II���Lw�ń<�E���Q�^D����4o��\�B_�� .��F-�M�=���?�<v3I�D��]n�epG
�J%�o���c�D��!���E*́�lA�R:���a�AH�.1㙙�I���ģ��A8�s�Dd�2ZM
��	1��gT��b��d\���}����,$�9>���|D���M���T�惎n!�3]���r�	u7���������o��A�ޖV��rў-��T���M�J�����ޛ��dϨ#2=��̬�G�9�����͟w�������j��ڪU��Tfϗ���	� ��dXF(t�?Y�=ze��$gc��U�ѐ����I84}�_h�ֵ�k3,��M���ܦ��_x��O�f��n�B ���m�Z+G�l�tnѝ�4�Kq.c�)�����%�
hm�تg���=c������;���]��ݰ�υ��+!M�L�����gzX�{.�����+H߉ � O���^(�if�C��{Q�q��P�G�p>��6;��w���ZS�V�� ə<��rBrZ����5IW�tN�N����=�A��˨9%j9E�Dd,U���6��-*\�ݮ+u���ͨ��f�������)<WxR�?Tgo2[C�}��&խ�#�M�s����a"�vL�N�s��b����?���`�(����Am���1��o���l~o�+ �<S.�@[�jĦ),++��mǈ�߮�$|kJf�`6�d���՟)�hui3(�dy)�~>=�5o^��B�k���8p�1UL֍
��C�Y[�{ڝ�i�T��c��i��1>Aϫ~e�p���� ҈��&�>�P���%ݽ�qu�q2��c��8��Rx`�*�ʩZRC�+EK6|�6 Qn��T���(��s?�?�͐�)i�0WU@!00|(l���pQ/Z��2|�\=���?�;ALָ�F�Q�8M)����^*qO�J5�T`��nϑ >�W�c�!E MA0�p��x��	��bN���ja޺|�����僴�lf��)|��A����	B�\����m� ��`�Sp����I��a���h~��lzaiѝ�uaQUg��T�JT](*>48|@�~W�
�Ub��� �.��X��;Z��ҽv��X����$��I�]�W~��������N=�]�R���sK�-���U�u9��pV�A��\���ӽ	�U��g�{�t�P�[�9D�	t0_4����x`��9�ސC�s�\S, </��6:q�6��/���'�v#���g���2�!�1��(M�����*ǻ�de'�gp���qdM�UQ��2muK5J(�18� ��ܛ5)F��+.!,S`fph&tW4p���EȬ�����p���1�}�Hn�݈eH��P?��&����C������5�YC�y�;7N�(B�<ދ����aV��umL�?tw�t'�v=������fI%� 	-0���Y��{]U;�?���_�q���}��|��ϥ2�,+�D����Y��E���7����d�y`�[�un�����'銠؍WA9��k�����1K+�ÑQ�I�.7���J7n1�%��]E���¯����J�l]��97?u��g㥣���p+Um<Z�-w�a�v؀[�]���_�qJ9��j�}A�[ܲn�L��:�а��:'��[p�EpV�fQ3�.�u{�ۘ��(�g�78O�/��,�x@�C���������1��}���D��,��Mb]�$�h�AS��;i?MOY���&Tx�ĈB�K�V�$���9x��P�^�smUa��"�Ţ�[�kG#."��X�R�^_E�o��>;�=���O֨l(V9s�8��x���u`u����4���}����T�PR�gnRnѳgZ�J�O�ƽd���oO��n���B�d�ZS�s�l�/�~��o~���R�1n���Z]�C��Rm��W0{Q��6utK��c�:ɇ3C�rd�zL�P0$wvڏ�F���Pn7f��x�Q�{�FAh��r�lZ��e�o|#�@����*��}M���W��f,���ty�m ���S+ɦ�Y+k��L�R�+�LrF\ɗ�$]���yO|��`K7wc���������T�pI�Z�bW���_O� �1I	��6�����N�s'����7��X�)������j�}�lm3��G¹��t+��j4�5���}`��_Ǆ�ΟɆI2��F�7olad�`ق��jR�&+ZH{�S)�|��kcǈ���a��>֒����\��$��7 /��H��g�ο �4C�j�&N������.q��\��,�l�X������X ��W�P��/پC�����1�$�o���]ƕK����'1ܾ�7��x-0�3�x����O!}�mݸ�w�W*r��X\�R&�I4I�K;��'�G������}#����:��� (|=���\�lR�Wd�`�8�~t��͚���ܠ}���ނB�z)}�M�:k�O�RFL���c�y����M�fH���f�?�,,c+)�}>j9�f��v�p}��Ӿ#W'��K�~�mb�þ_�"aN�;�S�WVk]Rx������fP!=��rY���S?��]6����%�\��j]�4�Xc����z����`���<V6���1��+��	�b�vn��Q��@��7��0�#�$%��ԶD&��l��g�}��O�)ƕ~�mƥ�;��B�&^<<�i3����>�㨊�������و��MY��Ꮽ�����/;��z���)6�!�aot:h!�c1��O�簉F|y3(�]䭲hT��Y���ʿF$�xH
|��i�_+�ISN�[GVd:U�jx��4+�%���:阈9�U`������T+-@T�6id`������ޅL_�=o>�������/�-��x?�B�;v���O�s�w����w ���"6B竮ev�������\�hP��V(Ei��c��Q��Q��W�8�����j�\�R]۶p�P�1;8O�����w"��BIqF�c5���֊�-eZ���=�s� �z"#��j��!|nmy�h�f��H!9��GdTK���I�HXwP׏@$\y�W�5I�gh���r@s�����堦�\�#W"y����0l2\�Q�T��#<�Άun����'{!dm/�y��Cg�b�+l��;a�1�|إ����d+��߉/��a�f��c��%u�zI ג�����U�@@/M
��؟.G�u����0m�/0�0>����6;��@���!���*�������|c]*@����Ĵ���7t�<�n'�@�?�PA!���_G�2M�h��O���F��yM^�Z�A>�1�Q�����"��I��"	A����2t �+���#޸DDH����"kN�)�R�� �s�2D����Y�JB�H���]e�gw�f�$H�GZ	�k`���fM���+$��̊!���8q�m�%K������
'�PS���5�S��M.� kc��"�yd�R�	��[g#�ѻtl���'�?��5���N=�,�+�}�5g�l�ه�]�����;�h��2�d�Z3w���m��"�
 ��]��]�2,��z�7�3��gh����zΫ^��)d���S�k��IX}Xr�q�����V�p7a�M���Q&wf@��Uv]y�+�����x<9�����V�:�c�n�Z9�\��#�jn&"���x6�%��>Fњ�5�`�X�Ɂ�F�� rpn#iʓ�����Ð����)$��(t��7渺RF1c�w}���r��"�#�p,��b�H�'���<Y��˺�|�C	���Q]f�+/�n��%�~��E�L6Q4��4����0���~#��	<�G{+?E"����Q4�g$�g�LVH9�<�A�K232BZAs�'N�[�Ioϔ�������+������\*>���@+��; ���[V�m���(G��Bp�K��%{�GZ�R�"�& d��X� ��;a�&�*|�մ����-����P6Nj�ݲ<��U �.E֟t����P��J���m�,Rb� ��H�D�����J�ܾ
X,l�����$�:���5�m!H�giDu���-��X�S��{���7}��� ١s��Ֆ7��_�
V� ������kP�i@���j���� ��ܢ
@>�9�����?�5 ƻ�Ss��Ou��xJ�0o���K���a��ɭ�u*�O7
��b@;�68\�h�C���&`����>~�/&�˓miO@j�m�5h&�GΓp�y��cÆ���L�2M�q��b�ڥ��H�Ă�e��$�F=��>��e����Xh�/d�b�'��w�ƃH잏�%��ԭ�p-�� �F	.�I�o��=��t-֮�*a�^5L��,���1߄u&�w��_���J�߽����
Ҕ6���
��;?��>�&��biN4e��Pe�!,�K@H�z��V�[!�g|\��l��ҍ�۷�
�MhG[�آ���ゾ,��7��KF@!<��M����aw�����D�?��̢UT��(�)������Pa|o����#����\>�@|j� ފYKA`�kF�DE��0O���'�AR���lT��_|O=l�|ڙW	�Vx�0ֆ~��^���(,�/5�l�A�!����'ɴ|��+���=����_�4h�I�F"������3ѝ* 'I�'�H��b�eHc��U���	ɿ=�dV�[h� 0��C���n��4�zŧ8�'�#�	Ԩ3"�^@�!hȓ�ùM���؃2A��r~u�C aCC�)�ۃ��R�t��6�%u=}��dŊ��++Es���z�M7{��ڃCQ��kܾ��t���S%u������K�@�����75�N���>|�����|�|>S�f��P2`��m#1N$�}[�)\<�m2�{m�� '�B/Ŵ%tɵ��K ���^tCJk���0�6�V��?p��)��kj�4lTt��	��G��Lܽݘ����<y�u���L.����;�<Q"�W��h���5����m��խ�|��i��)$��_,�5hQ�&|�1���7B�~9?�*�F����w6�/���d��ͳ�Ű̑*���NÐ<�e�)���Х���Qy�-Q�{���O#����J�kB,Cp5��2 ���Ԕ�|w�������{s�&2J�~��%���=]K���I¶R�(�&.�(�~A�:�MU/���������y��jd9�sf9'���;����Q���1i����%����S�2S�>	t�ė�Ӵ�ࠜ�[�7�!t���wӶg��;����D�^3'4�Y��_@г"������y������`Ψ�>$P1������cԵV�_�u3���qM;����4�w�m�5\��ס�q��X��'�&��+���%i.
,{��t{��*�vVp�ﶩ\u�o�^&YEބtf�"��6��F��8���.��g�F���=�.#r#|��*��7��A�U6��Ri�5��ӢiN�ObOV��;�ߍE���p>�F�X1?N�>/�)�<Թt3_Ћ���)r��2=�#$m�K��QB�F���o����Y��\�B�6��r	2���[���1sW�u���)�.��U��0�R�i�A {����~Է�Gi�"�D��z6�a�4A�d��4gI6����~�OK�Lh%H���Q����1���uћU��}�����6t�d0�$I�_z�`C�IJ�G�ͣ���W��)Usf��@��g|/[��uVa��R���Tz��D}�l���h�;�tj�<8<N��bH[��3b�y`��]�A���5�1���R)���4G�4���9�<��N9 ����@LL��YU��P�K�mĄ���8ы��DU�RTj�������'����lG��T��U�js&�B�~Ec�`�=��8-����s���Z�6A�Ñ�/9R��3�J�T\c�}�NoPM^Ηt�0�bhXA�}�L��j٦Y�8s�>O,K�.��T� T��R�TR4��y��;hvU[2$��+I;cF75��(��i��rJE;��{ Q�L�\�	��C�q�%|CإGg�~p@��9K��l2����R�R�?2�Rɇ�3pDf�����j�p�jd��u���^�@�s��\S��jQ94 d{�G��%�	g� e �z;�Dn}�%�#��}vb�}�7��`2���.�X�d#$_� �ɔMG�ǩ�}U����0%�Z�Ҍ����BKZ�&�t(�3�n�{'�ֈ#KЫ�\��Tk��dI�H����Md󀇈��e�8'�Tp1�>���S[�:[�.Z�̿�dVm3�v<��=A��ji�h�U:�E�=��gE��Gm��3t�u��[�b��g��2Sk]�B��*�qvR	��z_�`laV��񧕲�^�J����U�z��S�%"�J�7��b���p`8�!�	Y� �tFo�Ej�Z�-��������7>��X����O� ���cNQ�7j�nl6k�"L��t�C���YIvc��ctKfT���K�zc' "��j�z�>fqw�$���"r]�q�F����B�Må ��Ԏ�B�{_�qk{�������5������ȟj�;mN���}4oH���^��؜7]�7�+�`�e���}������Gl�9SD\������c�r>:����СDԦ�{�=k����&�k�L`&�5;rRc�k���{^Q�0lR���WM��}�7)�W���z`U����Y������+t���>�g���4�a2A~��!��S��amO�.|h�=��A�T��  zvxPou�g���(8�d�£�����b�`>5�F ,�ل���H�/�PI#��o�Z�O�ucހ�˨'��^��!�TW��/�1;'�����%�(�G
M��F�C�ο�v;G?tϦ>�#C���%��u�)�-���w�4f�@<LT���A���I��6	m֠c��W���֣�z��� ��ke��e�xN��O�%bpl����Q&_�jy}9��c��9��#{��=g�Ҁ�rCG��bS궰�.�oJ��迉O����ɉQ5C ���!dRN��cp�Z�N�˙OuB6G��7Z�k�.y5}�&�����jW#R�����)}$d�BaU����J@��T[��4���Pl�+r���"D6:��v�&�3�%͌'`	�xF�ރ�����\z��M6��i�Pg�q<�����vh�	��J����T+�m7��w�Ԩ�<O�K�r�\��)GC�J[d��38"���s�C��N�2��.J���\�����"��՚���V���c�;�h�6Yf�QA$9�e��O�K��( ? ��Z3�q��{v�<�2�A�lU��}��)e��^�{�|�<���~�2'�5[�ҁd��ˣHf(Ls�)?�l�G���-+�`h<1�p�{ߨ2�=����x�/��I4<x!�ϕE=#��c׸)�)�BT`���"X�I�ЇT�)�=쀇2=���G |K���05� +r�w"&�T���憍��c���9�C$��$L���>�A}EǛĞ����W8p��Q����Ȗp�Hw��sݟ�c�'�F��Z��=wo#�L1<d��'`�)6"�P�j1ݰ�	c�y�t��ME�I;�oKg��CI1�5'�lc��:U���|���?�o�����b(���j�ȟ.�b�#[�
\���w�j؈q���2��&n��U��V�M��Ϋ1*c]�>�@�YN�l6(������� ����-��6C��RI3 �k�6PKX>������3T�X��.�Ϡq��m ��[wCt5@�BPh�i��s���󱀡Xhb�D�o�����9&��/�B�/a��j��BCZ��⩴��4��f_M��K�m�r3��ZH&�]R%��Ӡk�|�m}�C��b���W���V=�h��vM���H��_�Ȍ��o��$�?:�����h��wv.�ص�G���ϑnR���%䮖6�`��7��+��	(���*�b"��zX�|��!x�̕�ѣ�t��6Uҝ%y6��8Yل��y0H��a�g�s �-��u�������\��n�c�3��BUl��ֺ�V]+pT+��#]���3܃nƌ1�J����ɜb{��T;*���*�y�ƨ�3x�+�0��4dl��M�˚,6x�j����뫊�G�˰�����Sx�vo>T��sŭ)q�#�qFɺ	�M�h� �x���-�إ�:�hy�T�NTT>�QK�m���k��0cy?
����k�`e��p�����|��b;��˱�����A�`\1����:$�� �y�O[t��f���r?ؠ�8�����W�u�}�`,�G%��m��A�a&�� �6t$~86��)��`���'ԍp��	k}�C�Y�4[�'�/g��[�� ^��_�Y�>^KW$y�x%|�%>��K�9��� 	*
��pܗ��@����˒���y~��y�[A��%���3��ʶ{�H	;;�����V�Fk��"��}^���NR�Ft��J��{�JR)P��#zK&�W������]�$Z���;���������'J)�ă�4���Yh}�� �l��X�iұ;���	rK�^�t�n�m���V��6��3-���8��kc-��)~����u�����'�gT��[�}�׾3�|�D�`�����
h�Լ��X��+W��86�N�pL��2�KԵ�H�_ֹer�_=��V�f���CHN��}k-V��;��S����G7��|����Wd�����4�}��^ĺ�`Q�H��t���}s� S_�yy���Z�N<�{��vd5��ʢ������q�SrM�A�a����/Qv�>b��"��X8_��5� �����4P'^!�_nnn�¶��R'�����P@1�����Z&�2���
\UҞ�^^�4np�Ƚ��g�#��/�����E#�sx�R�����5���DA|�Ƃ�8� ���i�'OS=;1�9�ꊤ����!S8�_&az&4����A�=�-�a����K���c��7��1��  vV��*�/-�4�b��((P��'��㘇\�/T��8��|O����W�y��͡Z�gR5���%��c:4��e�� �~EP�?3��Z� �S���A��34� ��|}U_姌/S�����.ꌋ�R��h�$��į��-��+�|%��U5#V�y����������>S��*���6v�F^���zU��b�5H@��m�vg��mr���	-|^j(oM��������Y��C��\2�)]C�y|���8 lJڔ-�a��0�9õ��J�^�@ֹ�0�k��k�o��꿼`��ƻ�B�vD*,C���.�
�$�4D���D��DX����ţ��ǳ!GZ@�b�L�~^�4g�ImL�}'���O�s�]d^	�6>��f���/P��W?���۾���0x�Ɗ�x/��l���{��v� �H�.�~�}B\���WY�ߎ3
����s����V���:�f=8#	4E���*S���.S3!�r@�T2OTG���w����E��c�騻o���Z��ig��JI;�z�"��u��ǋ�f/�t�W���Fg��#Qsy���'Lܴ&��*v�1M�d���{�d���B�O���J'@�t���;�l}�~q���j݄��h�������:�PN��� 8��3C~d��a���4��� �Y3��@�'�>���g�m�tT�mQ&��[L�Jf��l� ԯC��2�+վ'�ŗ�b'�/��GMW�|-�8����jf���y(zcf��-8">�O����1iL���M��O�,��>�S�/���Z���/��"�*��f^t�aTV�\hw@Hu�AE"V�%�'2��>���/��({�B�H�Wz0NHO�,�g`�Eͳ�-m����	�iRt��y:��������Ag��jd�G���m�r�=LA�%�x��D=c���S_p��E!TIG�KS�s�,�ܻ�g��^[�D�?�#���jm�{��ar,�M�q���=�u��w��I5ֿ�0R'�E-b����
xT�C����;k�o�)l�X�E������J�.;@z_���9Zp�Z�wQq�c��f���xP�ċ�>L��?��RaY�)e)��%]`1�t����'/{��Q��nN_�|2�}�[��E����2����/�2�j3϶9X�XO���7F���S�g����b�nSB���[Ǚy�Z��DDOƅ ���%{�r��
�+�w,T_D_�P�0:$Baw���+���J"W[�slޝ~�$G�-����z/����}��� V� k)c�{��� �����K�6}�3d�Ƅ;�ޅ��rM��I��Ϣ�]w��"E�-��y�f���y�,�7���K����]��F�y/.��W��7���!��i��	���G^<�#Jc��$�b?��G�z��e|3���:�5ﳇh��܅�\�V�_�t�EE&�`��q��NMiƓ��{-��j�#��e��M���~�2Rٓ�_E)t�Ig��>�%��&|����bW�| d���T�v�<"�Z�(Q;/�:Q����9C�&�w�4�oL՛���j��g���av�z�����cp��&��]ט�|�@ҜY@��ϓ_����;2,�K���.�����қ�#�D7:�V*
�G��QyU	�_1t	ڢ͘�y<�p��cdv7wN?1�Nٜ}��H����p�M�\�=��uRl5QM���9�
�%�!�Z����o|8Q[@[\�*J
#IN�s\���}%�~O���4^JL����W2�)�t�����$(Ц$0�BV�~�]7�Q���Q�z�QL��}%I���H��8���w����A,5V\�HV�O�.����ɦQcI����:>�;H���
g�r�v��}d��X���_GO�Iq���t��^�.5�X��t��cNv�\��>y'�Af��nd�j�!۾J�G�����N��[׃gAøMg�B ��ɡ.|��tD�,����\Z���kn�s%�&��\½1�)��v!�vǒ�K��X��� �dE��/�3&A+ZoZޙ���Z�:��1�S�j��Ř(rl��<�6X�$��Kb�D�SV��H���� ��J��5'��C�1H�W|����g���g8�rʜ(���g��~��k���k��W�WX��)x��4MEX���j�(v��J�-;s1����)�\){b5-5��k�jw�#�]�I��;;ǩl�5�/Wa��.�3pȌ���vF��q�±0h�Y�;X�v�}�8h?���{i9�>Ok�ɫU����@�
������n��NV�t91k_��9�SH9�)��^��	I�D=,p脴�6[j����5Z��H�i��^<�΋�Z�k��:]qdԾ�5���P��ͫJ��r�@8V{��'>٬���V���@զg�Vr�L�B���3���y�*����V���呸���Һ�lj� ���]<[q�܍�]�]�]��,�$b(�;P�֩vb�uJ�VD":��[J#eZ!��-�8;<�Q��_,�gY�8T����ՇX�]@��w��#I\u����c�J�� ,ˀ\�z�M����ȁ��0M�N��x^a���fI7ͼ
9��o,ݶ�$�Q�wF��i ��2Ah�
2%��}���>z"�'j�l| ��-�s�~��Si���]�a2].VQU� j�O� ���٬�Uhu!1|�A��֞�)xyc�`\+�����{��vC��?x�|��`���π	K��V��s���a��2�?�˚ڠQ1�����_�ț���l˴TYʰ��7��(%"��?���2sM����A�p�Wp_:���֜Wk�LU��^.��u��ܥV6��|���ٙ�,�G1W�~|ɍ�p>��x�D�2�I���HÈѕAi��G���4���+`M�܎��ڦ��?3bcǅKo�A�-F��Z��]��a��F�	�{�>�zf��}B�W�(�}i��J��ss����C�=��8�=�����+j�@q���"�U�;冨L+�����(
�W��c� o��w:7X���a/4�:|JO��{�ƤFcRq"�D)�V�U����t����[�����W$�;�c0�Z���k Kh���b?�n|.}IVP�������¨\$6�n�����e<D6V˾��;QAfe��j���6�En�����,-�߯k�{�3Q�ݖW�?(��ѳ�㓲��$�����k乹fI�2��ʧ��a�I�_�����qkH�����[{����U�r2U���QM�f�9�q�]�(eG5�hN�!��H{���de�#��ǚ�x��\�v�|Z7�JQ��彲��6Џ��s{�t�C�oTx�ş����l@�]:�,�.�a�C�,�ӗ���^23#7f>ȫf�}
I���c�ܸ6����,y=G��£�L�E��#Z,GI�����{�� 9� �Ο��CõO1)����k�E�$AU�z����t�n�钵��C��F�,����ڃ����V�s��l��P��Hv9R�y�I��l��^��;χ�O�q���J���y;�|Ć���u(M��u9)��U����o~�>l�2��)1S�L8��0�����+l��x�@|��T���U���\Z�/�����]-�j�\������ܶ�c��s����Rd��ݏ�9���i^`���%zc�v�Rb����ϧ_��l]���-�XY7����<<��˛�1e�F��a�J>m|=��IE�=�+�o�ZX@o5
J��֣'+Sm�B��v�8*�7�� ��r'��n�b���u:킜T�g���i�v��v'Y>�f��ܡ��4�F@p�j?'��v�I��%���ܒ��ے�󂢻-�f��MRR�\�ބ@��H�O���Xotѧ���:�ٱk�����>��Z�n�/���?��h�q͜��!1%��iۻ�W.KwT�8��0u�KH�x�cD��k�b�JZ=0E�׷ϡõ���`�nmu
N��Ή�z�/�8�Ippq����ċ\!̠��q�̃�.>���^=�����	( T�|�T��:'m��y����˼�!��x=0��b
<��иW*`��Ö��ˏXM�pi��t�HBL3�E�f�q�c[őE��/Ƨ>G��M�e�R����0��!�8w�0W�Ӝ|/�jr�����:Üþk�|(�޵FϺtx�XA@Q�z�i���r�S�X@���r��.�5�]���B_V�˹v�J��	���.�?�X��8(���?K̹;��Z���I����bVC��8��[���m�
~̘�9I��]�o\2Wu3[HiD�(��X����j-neB�g}�l% ��A�h�\�Q��j��k�"M�q����H]-��?Y9�\<sҢ��㊕W���9��b9p�>���M͍4����J���A�s�K0&jY-c�]],�)J��W�`��>�/�'�z�W��h��a�Y�JČ�Z��g�I�a z?�|��1�^4���&��L��O���dy�+u�����Q�sf�z���i���ȯ�\^�p��2Q1�V�A��MٛacVw��r_�����w�C�Lt��;��t�
��b���kݖ�]:;�y�ع�f	�ЏY�y�ʦ��r������J���D<�h`�kY��������/�}W�Ǟ_�gm�������=�PcR��nU�\u[ٖi�|��晝��&V�o`!���2��s�[��jM�U�D�c��C�{
)��1^�+v�|`e��U�k����!����h��乹&��Y�k�JJ����-q�o��M]��/8��Y�֟�M�ָ#f�z�����˚��0Y���>�_	W��X�P�9�v~��[����fn���恵Jw>��h��'f�яݢ�\?�hf�C�)�z����5׃�\ť�C�����A0��	�k��WҚL'��)�%O�� i�T�7q�.�;'W�M�3�|^���G���}g����I�X�QTn�Vj��U�u֧�8�?z��� ]��6�܎���� ր�8h��M�w	�>��1��[J%��g����Iܵ�5�Ĕ]��/%�%p(�'���Y��p�1m���Eb���Y�s�,�"��w��|}8 Յn�{��e�a�p�n�p�,U�D����vލ��*�QͰ��Y�[ؗ����ѡaw.��r��PB�DK���  �ʾWM2;;��ʹ� ��Һ���$��C�y��~*��/���i�v����uG`��)�����5��kB1�ą�8U;�}&�T�"K��=S��"������Än�eZ	�_����AhE�9����%g\B7���8���ߕI٫�H�����^e�n���\���#�@��j�!5\���:��d���f��"��=�-ڧ��E%Ud4�k�JS˵�4��&��ƹ��y�8���3x�����t��[5T%��ψ���$������Z_����ל�)�e_�5�`/�gAz�(�%ANtU�q'.ӑ�]:C2�H�2M�>���cȜ��J�Mq	Ά�O3o '�ԋEwq�&ת
�o�Џ��,3��d��d�Fw�C�s<{|�d�by~���� �b:��=T{�n�i-E���̷�>����DTd���#�ÅMO��3d�W	��{�/P��pY��݄U���jbO&�)�z�I����=)m2�z�t�o�d�]���1=\�v���Yo�[�l�\���ҹ!cI���{*�T�@�;�ڳ����9�S���b��p�[����k�TB��B��/���i2�:�sy>����eػ�~(������ry�kы˽E���
�|9#�;������-¹��>�8���
��϶��^�$GF���6�E< m4�~���}\f��f��ݺ~�z������t1sr�V{VZ&��.��)�|]�]k��I6������x�ã�K0<����k̤Q}Gl$�Y��W��N�>�j�]R�� �vS��LI,n���g��m��0j�'c⣐���'�[��iB���8h�o��u+�e�7(�+�'���뇡�W�
NU�J�J���/��<v�ȓ���R�H��+��U�ۥp�ZCa��%�k���fP:�I�#�Ν|ĝ;��X�u��c��4R2qc��~�#��Xk¾R=�BIx�5VZC<�1����-��J�3kg�Y!����%F�uz��xC��$r�`����B*��)�7!�,�_=��{x	�ïڰ�b!�ѥ"��Qh�l���
���G*7�u��+9�P�R�r��D=S���K��Ҽ�3���TI��!H�B��C�c*=�m���U��ׂ]x30a0���C�T`��L�2&�ϳ�0�� v�[w~9A�l%�f�u����"�o]���s�YJk�Ѡ���T�)ʦ;ؾ��'j������L��(^��U�F �B�t�x��maa�I,�J�u�̥��}n@/�~�晹�E8�E>
PK�=I�`e�5���'�{r]g_`�H�� -���gr��#��N@� ��2.�~0fe��]�Z�8���v�3�w+����d����H��
�]����RM'&�����|�-��Z�P��d��Jp�bK��%I��w��//>��ü�ଧ��y�B��Q�q\�S�q�h�c����#��aL�M���m��H�1w��p|�����S�*��E4.9��?�� �! >vZ<���(�垃\�#�t&"o�7?��������̩�#��ou߼w*2�7X�938�4|�As��V/T9\�^��y�<��.3�ƙ�$L���8m+ùþkѣ�k��T��۱hy��վ�V4ö$د�FH�T��/�6�4�s6�g�D��6�x��	������]1:)m#�
�� Ο���:��kyH�*��P�l> s�\��8HvgƙF�aS���ZQ.�z P1ZSh��ϡWLP����&�5�湑ꇻSwbf)[��<�U@�J�uL�9����+_���mR|�	?2�Hvh���{7��^4�>����@4�~�)	z�}�a.f��>2cu�K�څb����x͐��[�臨5��P��L:���f��`�#�4�1�_�
��1�́ŘԪ�����C�p���hMO�gd7wz�!=�ak�Q��_BW�G�0/G>n�s�m��Oɧ���n!/���:OH�unگ�}���tǥ��Ǘ���-�Ibݽ�R����MOj�8�l5� =ȋ�J�`3���~ld����e���9�F�G=N�!%�/���6;(�V,!<��r���_���páXVx���_6�"�3���u �|��,���0��1���"R#���l�����D_�L�oݵ}����I�6�S�.����o��Ȇ�-d�e�m�P�6HpK&��k�Z�o��|C��UO$Y>=���ɪD7�Q3t;J�*�	n�Sy>|=iQ�b�Y�*���cz9�����u(�<����O��~�n���yi�2�qT�:qG�� ]��B�:H��]�^lJ���Y_��\��Y��>N��;5�-�%(�7��Uki*S�+��y��tc���WL�>�	���Ν}�*��o�껗˄������d��q�FS�4�>������ebC3��m�Z�~��Z����z���񄧥���/�����_}��?�ᦂ}n2)V?��
%��˹�� ~��4Θ���I�/o=I��<�9�7U&@�y7�d� �⧰ZS���}p� �"΄����؜��r���Rm�.'9~TA���L�tK*�>T6RA}�-��EC�'���'u�G̦>e�&nK��98,�� �,���>������L��k��lb����`�a��*V�&��V d�*A^��)�?BkH�!������t �ڙ���`�ȳC� {B��~/�#�He�c�I���!���\_Ӱ�@�>�F�{g�1�[��o�~���b�����te�̉-���q*tq�=�� �]>z�cp)���HA��b6�]�5�-�@>��G޽�	��7vu�D��G+��ݲ���jS���Kd($���!e��b<���YX�w8e��/$�G��]y�A��L��X#6"[��ynWR�a`��D�a�Y�o��:�h�? ��˒V���ؖġ���2b��f�W	@�w�Z��=��.���0�/%O���N9�c�m^|�]DC]��s�&09��?w���� z+͜��������wYZD,zJQ�|̤<�aú w�� 1���p�;9�P�ƌa�����{�s�H��J��	��o@��@vz����Rj!�*7|$��<}�5��ZVr��[�C�(�͖rX8λ<��~{	J�1��]�BV<(	/�c�=�#9	�+�_�q��8��՜�o�!�o��*��Ĝ�:��&AB���t��S!Ë埐첲F_Ȃ��"�)m�R�r��-�-��$F-��^�'Ў6%��]S��kFOC��j�,�A����#ߑ��6>됯���=Tj�u[h�k���b��� ٴz�_�6�7D��|������2Z�=ϻ����9��K��ߎ2���0�V����M��ul��";�u(�w�7�Pӱ�e	�gl�{��m�w&>���@�x��IL��z���p�Ұn�*΅0��Hya�_�I�VJDy,J}������{��V"�H`� 
�e�oY<��/�7/v�Ǎ�*�H���IRK�N���3���U���sۃ;�3��HvbXmD篲�.!��K$����Nq�x��[d�d��IY��,@ҏKP@��|D�"�ow~W �!FGXn9ɸ��Y�b���7�]|ذNRG�Fl5�"ǋTG��>C���$6��u<n��޴ o(�W)d�#�-���n�ՠ��p��A�X��3"��f����g���R��jX9c��&�Ps���NI�'�xi�R����P��E��B�.v4����8+�H>�miG�-��$��.m%7m��~L��@�h��7�xqZ��\ϖ�{�$�6v�s�^�'�x̒�Y]�7��^�l���茚�2��VЉ�0	��p�Ȋ���C=ߨ���v���~a%�C��	π�ZX��)���,��j�/+���[u&bK�a |ݎ/^
n1�jY'>;f䚴E��<�Mr�O�
ԝm>���?2��Ah�%�m����{���bn����E�ـ���bzAv@E�YT#��P�lO����D8�L;F�%Җ����N�đ�<ئ�z5���א���Qʭt|<Gs9��%��Y-��w�n+����I�wZ�㨤X�S��x������H�|� �8!@^q@&?)��µ��xO���t��1�]�%�޴r�W:�/)ބ�P+{<�ɮ�P� �m��a�a<)Le덀���ٴ�,8�?O�`=�턶��:�ÚT$��_U��+�r���ZLJ�s�A�T�� �l�\w��H v����
�m�����Yd��r���X7��N���D�DI�|�Q6���%��qTunX@rq�}����V����A= �C ��Z�H�I�[��h�A2�}u���[U�ĸ��>��T^�xl|��/U���|#���Q�p�.>�My'Mܡ��o�Ӑ��}�V�Hu��;���`-��6�t��c�T[���(r�oZ��J�~ǽ^R���c��i	Vߡ͂�m�I @������\a+��M��)X����h�zZ��5lE�3S���Ƃ�1��κ�Oi�r���f�W�)��D�����Um7��?�w5d7'�;a̙i�~4���~�&Vvp���O9�U�F���2�)��5���+�A��0ZK�y��b�܁�l�o03���K1ѾT't��;w�܆T���J������GS@:k 2��t{ߒj˙���tm�����^�(��6Y�)Ks��it��`��O�]6�����I&�y��G���LD���t�*�L9��uu�C4����\x�4��Hd\'�szf�R���J�T��������"\	�V>qr5��E�Bu,G'�"-�;��W�?$B�������J��Lȼ��aV@�?ϣo�]; Lg~��Y��$� ���L�ὒ�`A��b:|�1`*y���3C烚1t+���h[g�w4j�_-w�����	�~E�kJ�=��Ź�h�a��m�?y����"�v����͵�����3$�7��z�i�(�A���;CDz�1A��mKy�m�C���r����~�XE�X�騄�.,��C�ZZ5??��_Q�%�w�(m=ԑ~��#c��L�X�}��v��}G�vo��ԡw�2�.w��3�D�D�9d����]4�<��7���3��,+�Y,
�X���=�Ģԏ��p�.J�)\.���J���eF� �N�h��v�7�c���Gqd+'�wi6��ʬL/�R�=����eύ��P�6�%���U�K�b�+�1��SW�V&��6C�I�H�'���Y˕C�rѥ��:N���.
�i�p�2�� �Qz#Ffz'�[����;�Rc�W`��rD���|��	t�֙�v��sq�(���t�K��E���������̝Z�~����rj�ACv��/��M������_T�6�g�u�[$��U�a�g�3�/;Κ3G�i�'���b�ZEfy���D�d"`t$=L
�&SZi�̺$iV��%#��P)���ԝ��&�fc���!�����b642E��R�̛5�C�
!��Su�(��2��t �[#@윻�R�գp#���P��8+����*7��� w��������L��mى��w#�'�(�2ژv}�	�f\¡��l�f��M���/C��p�S�=�bN\-�>��������ۆ�;�EZ�`���
$�1R}v��5�2{�������6��o�_yH������`��&`���.��*"@���Չ�"��E�h��)Ma\9��-�2��L�K5��+oR��ER�y��q47���U�(�hˢ�jV�;O�ba���g�qK�s^������o���-���l��=L� ёv#�>�*��.��֪6y��V�v�Q�oE"�e�$=I��ET�1L��s5}���48��U)�O�[9nf�[�(�x��&K�H �J�RWX��b����zb��L5�4��!V�ɛ&�&���	=*�>=|��͔���]�3`�,�g�I�?���%K���e$d��-�
A����a6<8ۻܮHi6C�Ub]/�F|�ى!�P7��x�m�	�$R��]�G�DE��^�l���G7����h2ٟ��.�T��L�҇���.�ծљs@a�!����f_#q��(MxHh���}k^��s�1;��o=��gZ��5��5�a+�Ɉk�!�M�8N�J�.�}���0-F%��M��?i�,(�)�HʩTb�}�=i r���{�f
�y�"Wqr}����ꊉ�ɭ乺���UR���٘�<4��I�같�e9��[+܀�GR��Bެ�#��{��j�v2�˧r�V��;vg˹���iu����.�'��Y�Hx��$w���@�B�T��F�CB�S}oP����+����j�3X,��)�v6@F�ؙ�[
�7!E�x��� 0���n������������]>�S������)�I��Vv]��:�~�4-9�4�[մ2>���r��eE,�eD�H4�>l�-J��d�m���{D�K���ȝ�@�K���9fU1�Ó����~4��V��ȅ��Ǆ1f��	:$�2����x�i4b���j�B�վ;��(�p�a?>Q�g���(��3Y)�!ѺV�U������HE�7,D�b���d@�}ܘȟ����=���'Xy�����W==b*��ӸS3�3>���u��5�z���R�I�q3��/Z3	�Ym�0�/�n���X�rl}�7�)�o`&�k�����M�G��G��n�uΙ*��W#�Rr�{�����-}��������c1�-?,@��[�.�Ŗ���U�#�&�[|V�D���b��_�'����'����&��  8�!�.dQ��t(����Vh���C�+��^&9�;�J�B͒�
m|�cR��O�/:�A<�!��s_��@ߙ�.�uf�H>�R�9�O�[0��-!�k��y��d�X� 6p˔������/�=��O�f�&9��1==�9 U	s����R;��7�!�k�q!b�+^���穅�	%pOӋ:�+�*[�Z/	�����y���C�S�|���B��tBsBs]�
����'��g��O�@�_��{=�	�M)⏜*vS"+����|M-]%�:fIK�)h�J���&���`���Cn~��K����pӏ/�[ƾ��э�.Љ�?�hB%n1������]h+; 7|Ю�?[���ba��TS��ubi�TM�̉W�=`u�b�n�7�%@�}͝�r���W1����V�a��,u���sʯ��^Fn{?VzR !p��P	H�?E$���B/�!�Y՟�@�K�`4�]X��,N�^/�ײ��_͙�%��0m��b�a����.�^�Ƀ�y��t��M�gpy)Dy�W�҇ڲ)˄Ъ���������9'�r2{���k�~��'�6�E2v׆���ԢX���塋C�h��(V����[?�w���L~_�� o�v��7��S���3��d���>N�l����땪�˭'4A�p��v}HS��?o�Tp��4�ʬb���F���t�D}�0�ϣ��@�RY	��)>Ϊ����{�?���C�l�z����lb�V�ơ�/t�N�U�>���/�r��z��Y����dn�)21e�+h?J��,�b-N�H��zNJ|V��y���t���b��d}���(�3�7u��G\��k�o��7$�P ���(�B-_>��;�1Q�X��+���?
LU����DR�7�EBt �O���	��)��ڕ�)�#��=2m+��PsY�K�B��	A�>���9�iH<w�Z^4̃Mfm�yX� 8�dx!�׀�?��Լ��#"��S��߄\���&��{��NߺC�O���a������7��Wr�6P���iƷ��{�E` �Zay�`�������r�ig�&rL�b	�Y#�zMe����=�y��K|_׍O��5�_\m[&~Lq\�@Ж���s���4�os�?���G�'n�O�"4,�}�f������e���g z��)��8>e ֆƌH�7=~�S� s�س�/W���3��y◌8���P��u9���6�� ���\H�!�Zs;�����x�6���Ⱥ,����v��z.� 4�\otS��Q �g0(xȩ���_I�X)����^�$�Q��/��R���Ʋ�w}���,�����A1�[U��� ���
2+� ����K�b&�9��g?��/�"�v�H��iP�
�5"@4��k(F����*[F�>��R(�hJ�!z��y��'/׺�}�\M�e$%�p_w4�U���do�0z���,xY���p�%o;�6���{���;|8����~�I�c���S����@�L������o��)ϲP���9�� B�Pv4,
��Am�Y�;��tK>���BoiB�j���O6w�_S��I��t���%��)S�Ze3�m^ ��4f	B��rL�ϓ`ͷ�w�~D����Y�m�ٗbq��;��&U�҉΃0x��z��ZC�w��\�,5�"ek���NK묭��{�����K`�/�0���7�3�v#E*ڧV�$�-;?x¸=IN������C���i���T���SKB�^�2ʃip��c����W"3_G���M��'w�In3����7���ݩב�����<�*Dv2�{ȈuѾ�m!g��*�o�Z>ͽ(�{����\�^U��ً<�EP<�^��qI*�4�0]Bc�T���勒��ƹ �ʟ�tj���	�s����w�����O���r���H�������
�]u��7������Q(���6�.�;�NX
��6�8[j�C&���=ܛW�f<��O7ɜ�h����r)_$�ȵ�w�?�̒��0|�����Ք��ňb|���8����lGtS�1���c��gݓԂ��m����k�V���ʗ��]�*�qB�������� ���G���`��H3X.[׷�:<-�砕���!q3���Zx$9��1m��aʨV���М�5��wJ� .2$�-�dw��WQ��;��?�$�%�xr\��L�5��&�SBw�Ɂ3 z<����MGO/ምv�����x�K���rx4���&����O�/�"�-�Gm#�^p�ɥ��9&� Y	O R��>��1M�qBμ���Y4UG䗫^�H ��60H��/��sˊ�b�dV(�w�LԆd��'Q����X��h���?_�$�	������75��m"��}ל�1�����I@�o�ֶv�}�(���	^axg��45�EZ��V�8%����[a؃��*���JDyq��br6x��"bT`=�eZaז��y7vԕ��B�����mWO��/-Tz}�N�"\}^4�֥*d9f�́a��Ć^��+�A� $)��>UN,%ޜ|��G�\0H�Egw��e2�,�/DD�l��ɜDA��CӘ��c>9�J�ݺ��`x�(+��t+Y�+-8q�$�<y>��\�T��� p�����z�ǎ��Q�P%ܓ�#�fo�S����/�?]��H�f�KP�![h<�
�<vE��
j�xAwuM}���,1���X)4��KM�D[��ɀ9&��8#BO�9E
����G�=��6le�""oyE��hg(����J��&��-	����!��ߦՀDG;��@N�;Z:P΢�z���}���q��q������u�5)���*#R�Qn�����LP��)i�%3��.����+*M	K�e�L� �>|;s��;�����ih��.��w!�DQ|䕍�X�i��Vf�i�qʥSm>5���-]���C�����DLX�*.����:���[+�L�bǟ�q��/;͘�ókW\�����P~/�t�V�ڌ��>���7�����k��<](9�EUO���\�짽V>(e;���oU��o�.]KN��Z(�O�Rl�T�c�k�}I�G���62@��k��W��;!�+	�AK �8=z "��TQYQ�%VԸ��+�LB�r(�q�G`ˍ���J�n��a��(������1	_ia�'z-�U��'��|���y^E ���!�r��[Bw-�}[6�W�}~����?�<6жN���R�����(���۽26pOp�CesY����Ǹ;�T�Pc��W&��;�ץ�L���B*. �1�M�׹����1!�u���J�����"�v���k��Wǳw$e�~��X��ew|	�]����^>:�c�����%���D�Y��5u}�x�Lk�!�0"��9����E�B�e�>�+���SG�0a��K���/)h\���C��H{JԳr�H��F��3@?��*�#�W�Cj�Y��jwz֏#;�	���Bv>�%�42��#x�S��h3���t��k���r�hT8�~rꍔ��ɑ:�b�-��.B0M���YL�d�߸x9���䕐��3�E�a�q�L�<�x���4�2�O�|窴���)9��1�b���-�
Gp��B3N��́�iRpV���4��|YeQ��g���)t���"���<ɱ�E��@�zvd����Wc�V(3��T�(r��
�"�9r�~*_8�;��g�����q� e�� ���t�-５�3R��X��#��ʙ��_X�_�H�y���	�X�ǆ�\�K�?~�P��6٠8��j���C,��o�X�,���]c���ϐ2�P���-ꠥ&=�*.[_�M,��-"��>���-)�{�!\EѬ��,�>n'�>�+9����M�3o��I��l������*�N�����}:�d(��\2a�`y
����Lɀa�X/ߤ�MS��݉+
G9GK�mIpt*;ڪ����O�U�է��B�,��JXRU�&(����U����$���d2c��?�PuHq��5ȋ�(��|��ɹ���_�׌҇�F�ZlJ���Nq���N���������v�;"Y���G!��(�\�i)0��g�+�>��(�U�Es�9��9���/߭N�RA�No�G62C���<wx衭��/�v"�(i��5���H34�Ԍ�wo��gh��~��#1b�N 7�eEf?����k�є��L�S�9��}�k����F��q�Q?�Q�4��tiIu��;Sc8U��d�3�?�N*4�ͧ�9}(�'�2)����{�ְWUS.���'��Ffl�7��e��a����	#��_ &k�;������C���.�������L%�ǧ��Y��U���>e ���̢4s����נ2��*�r<.�ӓc q�z��&I�P�{�A���7rǏ��W�ǭ����kwUYoe��ب�EC�+�0�|g@h�Bs_ۯ��oʈe�t�wVy/�33�p5�1��G_0Gz��g;ou��9�־(��w�*��Wz*Hق���������ym�2��>��^�3�i��\�&5$o� w�ʯH�:( �&� �i��~��(�+��R�*��>	ֺ��\M����&D���pR�P��X���9����<5t^��4��J�gn����7��(���,4��xB�8=��`�P�Q�&־1v�"�,Y�6�!i�OP@��R�����[֯��„�> ��z��'.���K� ���i^�\�{��� ��v���[�)^|����S؅�����gq����z�`U��tD����#�!bQr<?$+~6^�N�ȷ�ZT\�m˴���c3��ە.��%�|�Z�Gi��GS���tB�D�ܙ��Yᓕ�T�o���<S��E� '��O�S��U�I�F��/�i��'й	7�����m��iN�;Ugr�ܵZ ��W�"�9=�������Y��|��,ț3���v��}X��˦2'OA�Q�Gh���U��`���~�}
��^7�i���ր�Baw7��լ�P�=)��p��8�Y��zľힴW����=pG�"��H8��~?��9�R'K���B���sH��ovB��Iŵ޿��vѲ.r�Inz~yH{۷���A�"��܎$^� �N_q��t��٬f4˥'9,w���vN0?�̙���;͸�mDl@��3Θ�
���إ������z����y�$���,d����ڶ��!W-����,O���X�5wp�&��ѷϯ��@�U��u�#x�A�e"��婺&����W<�U*�qM�
�Q����	=z߳�0�����?�[^%љ��70-�����Wǡ3�G�3�pY�R�Ѓ�=,���IR*�u�&)U� omY*|�n1v�q�w ��v�ֲ��E$�kJ�ߤ;~��X`���Z|A�8���2���Lʓ�ř���QP�t�G�.J���)��t�ZA½� �Y͋~���I�·�<NC5l��$0���4$�GD~ޭ�d
�f���UN1�$��y@��MW�|�o�h��;�6ݢ�qu���uU�-j���>t�ED���z�R5�s�pㄸ�c������aQ�\�,QT ^�B����V��+��:�jK�N7{���	]�9R����THu(��|<Ȣ�x�� u}���]�ۤI���A�XΟ�G��Y�hɌv��b��M1�I����L7%EP��X�il��AeW&���/@5Sf �zi��B��p�|��[����K�K!dIŞ�P䯠1�5���$�xbE~V¼����2�ƞ�xn���
 2t�!ip^-r�:�J^���.O�s�K塵q�x�����upSbj��[�n������{��>.Z��?s���m�i�-�W$E�
��
m����Z�U$Tޅ�/�+W>�X1
�����oUOd�L�!tf�z�{@�#�}O�E^���5̀Te��DT2Œu�ӄ�F��}w۞d�9�\T�� ��R�5%��Ik��f��G*�J��-�-�/Ǉ|z*�eTSI2��!��f�J�Q����*�/�R�T9Lե[D֠j�
W�/?A�Μb��=�}��US��t�s�k�⨸�kM������}4;U��/���[��*�X�:5/(o������2F�R���b�w�(���O ����r��Xn�'���y�v�(M��6��⃋��
n�@L��F��z)�h�����={�&�j�_t"�x��}������b�ԟG.��S�P)έ�Y��Wy�ί�ѓ�c��c�e���dB/��I���F �Rq�9�u؍V�xS�2?��[��ݘ%��Lpݳ��-)�5>�w��꼃M�\������>h�?���N3]U�!⒑�u�W�@%�)O��Z�5̦�7������k���@��|+����)g	ZA>���|�?�ف���)E�`G�W�C��d^l��8���Z����ݔ(���N�i.��c��q�,P�JP �ųr��B%!�xc���-k��$��6@Uu��aO!|�C���X��JϽ�ޮ�(>�@�`�ڛ�\�]��3�Q��a�H�#���(�^��+&�d>�E\�ԗ����rY�O��'�pM��S˗��88F�f�;����?h+ �+�Eƿ��|�����B%-�|>��<%����]�E���z�Z	
��aE6*i����q���������LBadk�# EH��{�"��co;�rʱ�:���(2�g��8�����R^�j(�-��>�I�����O�� ���E���2��fꍮM�t���D�����x`Hi�O�I)cv&
G�˴%m�w�H�����ɸ0 �[�?�$�#E�Ѕ�R�i?����XDY�o9I�S�M�9�99p'����9���4���
�!����J`�K���\��8�Z7��V�l��uU�8gA%���|� D�k7�C�z���'�\��[\��U�����}�Xuw̓��l>�|�(�E�U�`L����z���GH�b�pw-����b�]�z��87S^gJ�#Ҁ�%D!�m���E��g�T�\�E��U�� �3oI��V�Ī�53�X��f����#	� ��`�7tZ�h��=s�&�L���Dd��p���!�q��6��CjU6S��Y���;���|Bw�Vi ݉Ur�!' �Shh<����&2�&�˨�0f�c���٦}I���'��%^Y=� Rr������ͪ2�d�W�+�w�R�c^eq���S"�A��;�Vg�a�ok"��E��٠�o�Y˰�	9�@#^���M {�SI�bw�� �.�V�Y�k��9W+b��v����f&��S9u�ٕ���%�i3����6p�:8-V��l�7�(I�!�0x��}�S����eBS;�ל��@�!��������@�4�7h�Wr��l����
Mfqx�>�9�  �̊W3u^�v�F?��9Ȟ>�Ho@q?
�l�kx�7�Jz���y��x�a����>�6g#D�kԤi�i;ڳ;	��1!NO�;�Nv�q%�5h��nZN6[n��l�#O�j����6z�m��2���q�y������7���TRK���q�8k(ǵȨ7w�4�
͓RP\
y����zB����yA2vb�,�q�+��O��ߙ/���Է,��K:�ӤF&p�48r���)��RB��6$�4�I�^-3
�.�gk�~��6�+E�9�L6U�B�w��- �������P�U� v��vu&�V�S,�s�}� 9|��\�}R�<V'���l�:D
��06C��&L���o��o=ڻ*Lc?R��mD��Q�̫�?w)@�ůC�X>}���ҡ&�[{�R���T�� ��C�bT��T�;'�Ly-Լ(�XH#���gp�'d-@���#�i,�_��r�A�2a�d���l�P}*k�����I*6^$�ˁ�:�Z��;���{�W�n����H�b�@�7`�IV��x���CZXNWW��<G�4��D���|��./`�nPD�+~C��ڤ>T`�ك�V5�@��E�+K���ί�Xb/y�d6��#F�2~���2o���F�vҳ)�F���Al�"���I��	sp�P%�h(9�����żz�_V�K�x��L��5ޜ�oZ~]��0o�i���l�庿����m�c{�
A�t���5�^A��0I����=����h��M��گ�q�S���N<T[�P�.��@]�"�]?H���	�ܦ�5����.؉�ok�@���t���� Q:�Hyo 1��3F��+E�t���~�-|ŝ-o���>=�]�TY4`�N Mo�M+�3��`Y�B4��O �}ɭ)�������@u�H!]42hm��K7����z�5�E�A���^�;�̱_rD��y����:��ϩ�"�3��Ľ�=��/s��sD^��JFẈd�v�!�����!"D���j�6:�?UH�Y��EOi�o{W"��Dɨ��O.?�fY��RGA�42�xe�҅4,Bt����2U�X��s��Ab�UZ�ѡr+F��$t��td�P�4���*��Ȝ�i?{ewW�3�rͩ\�LΥ���Rڳo���E�}#kX�,}("��dC�D�Bw�+��D6�Szj�k�nY���e�X�FES+m&p�\n���:���5�p�%���!=���Xu�����3�F�nd^����O�]u�ճ���H;Ȑ�L/Q"G4��u�
��q�O�cf~?����4��	�oW��5��y����F������]�̔Q]�Q��͸c}�B��3p���d͗vD�e3dQq�Aj���p����!���t�xH���v$�C��z�L�p��$S��Պ�R	���CN��>�W�RR�]]�V�V�g���২2���D1��G��c�jy�V�
�]��_��\�(��$��(3E?�d+0��
��r�߇2��q��8�δ�&	��l�p���kI8�[����Xdj���1-yG�O
yǤ�:wӲ�a��5�.������	y���cɷ�:Qt����k 0e-~i�D��.~}�>wˣ2v˂� 9+pu��zD�4�lA�6z�Gl����/L"�A��r]̞"��T!2��3Ȅ&E�K�g���N\��w���h�[�7�U�����1+�ᥒv��O�'�ߩ���I��+E�r ,s1��HR��B5���ZĿ󺒧��r�$z/>0�}��?�{8	԰��=�ڴ����Qꛕo��������N;~چ��j����R>��H)ʏ�Sav��gk]y�bRp	��X���{�M"n�ݔE����TAп�  K���۳TIX��i/��m��&(�?��Ģ�\�%��!֧	N��B`Lh٬�2;��Th���HU�>��L��`��M�j��ٌ���C����%�c�Ǳy���E�1,� Պ}9Y36��3���>C"
=k������/	�L)�㎭]8 y5{�O�oz	�:�2'��[ɵ߸�:mN���k`��_?ی���'D䯭��@~/5��GU���\QৼL`���z�ӊx��}����������t��u�D/؏(j-ʹ�23N���A_��ri��1d0��liITO P翤<N_��j��<N��7Ȃ�A��JX5id�@Q[U�����xL�#x�K��EO��>m�:3�O�3h��NW4���Ax�SvZ ��c�}ryMje��^ʐ��A���(>�@N!#r�o���3}3�?�Z�(������YH-�HK��8\�vLRJ6�-Ő��L:;W��?G&2w����4{���N�|��i�
��`��������d�j��U��Dz�Iݨ򱗍qC���!eO�wm��Llx��	X�����9<	��x�w0��~Q��L#���a �ả�� Z w������[�qYS�a�x������&��L��GB[9��=."P4�=�hsl��iI`V�ks�C$�C��᳜C7֩�,e���-�cw���`�'������4��:�xI�(���`d�Rk9�� ���l%�Z���m3d�׺q���< �?��Zlf�!�W��s���/�z��Gϴ;>\�+���|��Z[h!^u轀�yI�'�xs;G�m��@j'�O�������y�w(-�X��vIҭ1�.'�%��.�ҡp|����6]:J�����S�[��iJ8Y�;���4�ե�ٝ�lD�pK� 3��	_��!i��:(�ޘ�O�ttSNg�%ˉ���N�AΗ$x����1��ב����ċ��hr ��t7�bd\*4Q�ď��%���:)� '�k�^�ٓ�	q�G�7�};�u��� �4��#�+��}"5��\տk�t���c_�c)���Kh���r�}����u]}��g�����O�%_��g��A�ڈ���w�;��u�\��*.��3x��J�*r|R��Ue��CB��Ck�����D�u4�V�
�{)�?��T�<$^���z�	A��$���T�������+m7��G�%&�8dVd�@�Pm���V�7I��K�`����:L�n�Wk�;A���5��|-}Y�%<���i�Wt�%Cq8�I=%�
mOqB+2�A�A	Y��t��;!J|����a�<��vsF���$�� ��|�č����nL��!�"@V�­*��H���i'���b����j�Ӫ����L��;^N*�N��w��T���	���tK;:��s0�\{@��䱉_�o��s=7��_�z���Ƴ�!��*�*���|�4wZ��,ֵax��āԬv��k��0����}&^�/��� �~2�-T�os^n���R-�{�,�;v7]���� ;~�>4n)�ۮ��]+8���iJ�l���,Q�q�uĮ*��Z��<
L�jD���|���Nq�/�i��$�i����rQG$sla��d��bj�M�&$g��	�6�������ĳ�{�Q��}�L�V� z��Y��qv>)W�P��¡G��r<�j:���Z=�2[�F��b#V��y\�����ٸ�W��$�(#���Q8���Տ$�a��˔�(�p�u8������IT��of�H!�Ճ������G���.��
Bj��>,D���?� Rz�`c��ʦ6�Q0� �!�*aj|G`M����[����64Q6&`k�9Ț�L� �]���8�z�7�D+¿ ���8���7�V=�����<��Ȱg�n����/,X߰� �ַ &Y��#��m>��'M����C���o�
�/'�@#��~0�v߶u7�u!;���,�)��
4:Me8������Ij�+&ȃ�7��Jt����E|	 |;��#b�nMԲ}w*ӱ��F�����?����W�'�>RE����O�jTrt�@�	��WQ��UE�1��$�0,��T�x���7�\���I�����,�t��JP��~�l�C�<�77�w���.�(b������xra�{��P�EX!�?����m�.��&�ЗU�F���	r���Z��F���Á]]Ҟ�8،�mL�U��<ÂN�ƻ�?��+��?����7�,y�W�ܲ���#^�d��)؋;7pϛ+_���-��G�X%�.�����A��{6i�cρ�,=�o���O���,(Τwyz.�׹����UW��E4���K g=�����dC岷*�_�ωKߓ�U���ٽd9��|^�6��=X�2Y�IŇq�-�8Ĉ���J-e��&�43ƃ-0���p\+t�Zy���k���Ԑ�$�pI˫=��:P��*��V��S��)6�u�b�Dg�Q���ê;�o't�T��+�d���I����>UZyGCg���j��<�m��}:��]�";fDӟy�MN�!�9�ǫ�<L�{��j�|�uzUVz���d{i��8�J�}��j�'�a�c�	�i���m���"�~R�9�Og���bi�QF)c���%2W�DYA�	�#���ܴ�DFm�̟�4�O��D;� *�r�Oa8���d����w�6ե�Ɨ#6(#�tRhܒ��W^��d��I�zw%B�����V,5.3@O%X��x�B�gE�z��� �x�t8���G���}h���b�!-�V�<��
�2��l��N���$�ٗ`�|)0�~���b�6��j;�� �j�u�bN:�+�T���&��p��k[ӏ$�Iv[Y ]cb��&X�ÝJߤ4��+�ʵ��y:��U7���F��x!��;����.��NJM��L�멼/;E��
��~�9�o�e�-�&xX0q:�ˈ�GM
���/�,/=E*i�
��kR��裘���P�;�jO;��Kޘ2���{&�ʗ�+}+��4à�b���gi�;.��U�g ����iڤ.���$Ԉ~K6�êeV���1ں�����P��x=�^��0W3��k��qQM1٬zd��#7�.I�!�����s�]�ҍzD�|�}M��
%�����"
��A��0�ڌ�Hp�R�̵�H�	�V��ݲ��`�[7<��u���gF��x`����)�>"�j�Wu�Y��S	}8eӬx�/�F8��뙖��m�� 3�J�b��xN��]�`����U�e��>�RY�)��1�R��W����"VG��WϔC1�;�*_FH���H�9@U�x!ӕ�^���M�t3�s��=P`b����\a����(�M#����ێ�r��-�tx
�vį���Ρe��S{zGT|�9�5��f��l#�]K��(mp]���XـK ڳ`l�f���$7}k�QQ��_aLTIZi��>�(�਺�^�ۓ�2SP�}1��a�g�~Wsy4���q6G�)��]�s�wHXp��GbJk������D�*�G-d��po�+5+VvI� 47O�8'�?.��J �Ĺ&��A��[+�.���jE��;�3�8���,����9�'Z�s4�ᘡ�EY�Y�4�Q����E�t��>E����z�������{��K�(k��]�L {��0�Ks��e\ﲌ��Nmx0Y�p�����Hl��9bO���6�$�)�V��췼>)��)��̜�"����|:`� x`"�c(���`^G�o��&~su�>�%� F�e ��>��2�Ű�<��۟2���2`�4T���9�\�޷�4��V��v=��2�S7�a��4�r�5L�$��-��-���y09�w�:
e`�g�&�-��$�hk�>o�I�a�O�&�&e� |�+�����G�rM�7�(dh�A��e� �_TgЂ[z���1]!��k�UR�11??k�؟�I�ell��Ⱦ�Gw:Ø���/�N��[�[��^�\��)2sz���Z$oȳA|F^��^E������)T�8���? 0�Q�!{*tL�~; ދ6]%�|�p�&o^�P�Mʵ*K��嶝NZ��u��ڍ���JE_yY�΁�B$b���(����䢲i�7��͊F��A��N�sn+��6
Q��]�r��W�6��!R9��+�QN�lt,��Ǖ��%�'줭�u��T�n/lv��Z����(X�88�%g�����0>�+�hV��M�z�+|� t�� �i`���������B���e����33����ӧ��SQKՁ����4(e�0��u�,�"3�vf����]���<~�<l3˚J�.�mL���dh��x��7���/ˋ pf�h�i���!B�]W_C��&���W��t'�ѿ)��V��5bq2˴*M!ĩ��"��$��sw�{&@�@4�ъ�X.<I$��h�]#h̕��Aې��R�;z�v�&��4��l�$�=d?^w�cvD�n�T�����D�@G��kjܼ���f� K��d�}����sfF�8P�2�����E����nآ�Ɔ�ʴ\�����U��g��?�U
ڨާ�f�,B^�Q���p����T��9U��r��E�����ŕm�Ƿ�$�n� ۿ���g�W�+v��7�=�Pu�h�5ױ�Z��2��I�-���%���qs�V�x7�0j����k[�Qv�b����'�@��Jz�h,�|Lin�@h�0�1��%<. ��P��D��̊�x�2=�D.������L`Rض��H�fF�Þ�[�-���]R��ɳ��M�| �vO`%�_8�xZ����s5_u����H�������E?±�*�a��I����[��g�)������/lN�M/����z�g��՚�wjR���k�<��E7���B�@,�6�̩�A*w�jP`dHV��]$���} �dyW��?E�>֑̄t�[*n���L�ܬ���=iz:9J@�0r �=��_B�O��!�T� �h0�������Q��V�>��C�֎��@��S��#E���&�Bz}��D�쌯�o���:�Dɂ��	Q`*�&��z���jx����d�F ��\���R@�+��J��tlj����\�����m��I5I��H^��R	D^�hOJ=Ho�W�{�����`��H�r�6T8�p�8�'p.��1�
I`�x��Ւ7��@���+\om��4sKr���{���m�#��*���!� Lbk:�5�t��L�y���2
x�D���w�>e?��R�{ne%�E��ޖ`�����������^��r�u�V��1o�:���I`��V!����S�]{�N�k�R:�|�{�j�4�����s�؃t��)��/47�=f4@~��eV3!�W��]1-��.Z�U���1����n�D=� ���g���f��ϕ%��O���C�E߀ŕ���>���O&j(�C���6�2�i[��Q�U<ބ$���Q?r�|����|�ij2C[�V�\ O�\f�'���S&�-�Y�� ����������PCtD�f��ovto$��ڵO����q�Y��q(�/��(7�3^R�j���O��9&Gy_�'�q�����{<���6ZJ 4�ߋ]�Y�	�4^Ca�.����H���9~Q��SCX�8Z�(��=����q���!s;�۶�:R�A##N��<;H��daHE��7���=��H�miB�g�F���Y6�� ��-m�e��I�J?�!_��ul���nR��]�e9Z  K.�g|E���ePm�O6W�d���;z}�hK=��������r���˨܀�Q����e^�K5fti��E.��rO��wS*�Z���:�oEZ�r�G�U-��X�R��˗�.�8^�܍������E��{��'Pz��#Z����	ڔ���y��������ѾSG�B}���.%m���V��hp�j��&��9�_�pǅ��Hl�$@+��OG��	��߉̉K^g�rA��O*�������?:T6�tW���w#z�>4�9��$^ٿ�X���`�r�� t	&G��ԇ`|��j� �R揈1��$,o9�=��n:����l����PU5�D$��x�fum�D�AIg����B���x[�YR�_A��C��`_{����/6���u����.\y�3]9Xfa�	�.桮k��ܛ�B�J��}(뵛|+\���g��,�j�ןJ��p�{�=��p�}�1�����O��D�J��d<+���?LV�e=i߮_ef�����C˧�&�����Y�]4�$d;���|�$��G�qr{���T�v�*Ũ*����Ԩ	O��@�� 3��ၘ��B4[/���Wag�֍c2�[u��mˀ�@��vcF�ǯE��?�go?��m�epʅn'mR�����~��&,���!���B�|c�����pr#���p�l �w@oW��B�@��x�){����a�+�� Q(2%!�k0�m��[�s���s�� �+��R-[c
g�XR�q"��\��,�y27�N$&e)z)�+��{�{�����%��@�7��h��:H����ZP.�A��B!�s��e� <β@ج�|����[M8����8�)�m��<��k���A� '��W�~	�����N��Q>a�Tm�M AH۴�A&ve(�$n���+�L6#�)��ba�3��$Ǳ��v��!�W�p��D�(�S��&��5�n�{���Lޗg��E0�^�[Wݨ��Wrx=o�N�j�p�m�3�f�fl�aU���Cn��C�x}Z�u�u�
q���nҷ �%H��C�W2�h��ncW�eU�0K�q�N1�6��)k!�����4�7���n=5�����u�Ku8�D�x���(�s�"��W�drR�bP����}�?��*�q��h6>N����0y#��b�:#�F����,}�+���{�8�\xe�z�\"�;&`LQtД"�R��4�$�6.<&�.�E���[q�x�t��J��i�y�Z�d��3�Q~��]!��r��֪]�F׵������L�����X�%�aS�J�X��,��Mj�)��m�S �_!W��e��O7�~� B%�o� ^�Kb�݊ɘ2�������x���};��nj�^��DF;������M0��A��n�C���ܛ���O=.0�'�Q��㌓#���G��G��j<���ĉaPG颧���b�E2��UcC��[?|A��׍KNmb>'�H���355N���\�3�`���?[��(��c��t/\g�|'���1x+2���o��<,�I�ˡ1��9խ,���ͻ�B����.�ߕ�07}�����z��s��R�gl�YڤE�z��8�|��yQg�a5;�����5Fu��Wtc:�tݬ+l��g
	����4�;��]��g0�� ��*���qe�"U�\�|}HT��`��s}e��i�1��2"w�DݼnԞ]q7<�؏�bQ�i�Ja�[���J͇*=���Ý��f���k|o�V���̻ZO5!�@�q6#�����q�D���+����A10w)Q��M�3,x�^�N%z�����	�y���IG��l���*ד�:R��C�����I��I�Q���ٿE�]��Y��%�e�`��Z��:J�(:c�hB��V�,���z���4�v̹?\\���<����L��+	+�EӘ�a�E�<Wr�]Ft,�V��V	�h0�ia�b�IU#��I����!�z�	��*k��t�~�2t���ŝ��s�_��{7y5����7{"�����w��Ȉy�;K�a�l�o�cs�S�����#`p\&.���c$��%��w���z��r��M�O�����a�p��С� ������D!B�v!?S����E��<pB�k�"��IAT��l^���Uo<x�v� 0����Y�56?��",�X+c�ԣ>Τx�<'� f��9�o�|^�(��Zq�`f���w;s��&�r�U��[��t����z��M�g1A���JWL��;L��6Otl�Y����5/'x�ߣ!��y�UAÔ���p��Ӥ*����M�/p� �*XBd����'�>���4�R[�`;��3�"���L���e�bcŪ�B݁8�d��$�/�ic�?��6o���F���2�����	�Ù�r�g���
��9E�]����]dC��A^�xM}���C���֧�'ӻ�ö�9�����x�n;'ş����J���ע<����3,�/��OH���=�i	�C��L�R�Oݒ!l�5LV��|/�t���'_H��3�末����]=b|xi�W V����G�4�Kd�n�	"_����";�z�9��ݡ
=LaNՎ��r�*�/C����Z�1�
��W�zWӜ���'���KSE�q��4����^J(^��5����S
L1�G�K���=%��'��2�'MD�퇡�������g�e %��zH�P%u���vg�������(dK
�sj��h�%��
������L��N�QO�����j����nU��?tY˝���*�ə$hF�4J`{M	Պ��cT��ܥ�! ���T�����@jH�,�����������E��O�mΚ�E<�*�I��<#�W�r	�puKɆ|���+qu5�q�}bb��/�3���
��N�z�ĝmB�;�)�3g�X���i��nz����Ku��g�h�wY+&0s�<�4Jx�A��|���+˖�o��b �;#ʑ6��M�:t�+�x�s?y{T���(�|,�{���\����5)Y�4gU,���WK�k��6п,C��is�~Г���7��0a�Ku�t�����h��2�%��_��&5���	^����p����p���l7��ӡZTbq`C�wOU�:�?���j[�,BfA�a�!��E"�ß�
i���%����I�֭S?��:�+�ְ,/�.�ٶ�i�}	�0���eȢ^ֶ̂iz�n�����~L#c&?Ck�\-�0ZS$#�f��+���`*Uvl��P�`�����q�-�pG��L@K��j;�g��J�2�0�x���w3��Q�	���o�����淕�<W㺖����]�P"���}|��o�<�G.[~�����/4;�|0R�[AO�>`��ӥY���ޗ���
�6[6u^�x �6τ�2�c�У����ŞJ�}��P�]���-�ٵ�C�}��:F��?W�e߲�/p��E���	�<}�[�/����oF^ c�,�+���ao�槲�M��^ͶD���'�|`��XO9Ą�v���U��qs��8 �w�Du
���DX���Dm���f -h��~H��m�8M�/��JW�1�}��M����`��>�����giTj��*s��CX����l������ EZ�6J����rF��S?�yz�� n,�	x�h� �<R���ՙ
\n���z�zP�Jt_�h�ܓ��?׫�CJ��D.�&��ZA��gj&��$7K^�(ɽK���k����d��n�R��@�~k������ҿ�FXd�v�s�2�[�NAZ;���:3h;�T��|{bd@���$Kpj�J ��c!ػm����G��#��S5'6�/�Q���N���B�=)���$m�䧾]��&L�Y9�(,���sH��G�:�W�5����9��w�s&E�-��8^�����9#*:�ˠ�r��\��7�-ڷ�w�=��7��~=gBO�S�����z:L'y�e�˃���0�C�E�jY�c7h��Ob�Q��ųJ���{*R��f��Q6u?Kv!/a���aG�G�y���q2�P���^L�y�[H�цVfUM�Ј)d��@H����T�v
~�p�t�3f�f
­C_M}��0u�y�e�Q1�D�]E��|�p4F($N�vn��V3���	г~L���|�A�_	:�г��e���ߥE��6�i�(	*iu� d��\�*������[/���έJp�!_�Q��ֱ����N�S׺�vr�-����x���h�x�/�L��/LYzf2.Ѐ��+�����73��"G����X���}��)����_�	���y!����+��C��9v�����:�t5��d�_�.8��q{.�6=�ژ������'p��&[���M���^��J�}4����K�����l��'yn῎)��<?�m��ΛY�:�&vm�����:?�*К�"�t��L��I���$��N�r�d�u ���5�f��C�0�l d/���:���Mt<��f��GvS� ���K��q�{�4����]������W�%�T����#���H��Bw��L��P\�Iݻ^ 
9l�D2�Bƣ�o�n�Bǻ΅��|����a���xC3ʿN��++b#[r���3�A�d�LK���P`�c,H��A8���Y��v%�'@&�cؾ��c��r4c�������`�D���O�)Ek>��?.3w�Ժ<����k��u�I� �Ài��^���g`Є���3=��0��qq��d �e4�P��U�h��SZ$}�S3�֐@����6�g���.�6�.������?ۣ��]���x?�5*d8�8���Z�X�M	(N��/w��;��#B�ָ�~-�4�"/�H{���5o��*�2��P<��?�I��SX��ݾW�g7*����}��7��4��Xe ��[���â!�y8����v0�Bw,�A>���̐��ͷ�H#Ty��?�+���:�����}����T��ϱ��!S)F�y�eX�N�Gy�4����@��o,�Kܔ�iN�Z¦k��
{Lv�8r�=�I*z���<�vH�W���hHY �MiJ����0f�y/:����7T�󰰶��g>Y�d�5�=�AP ��(>ey,]R'���r�y�X��yEhe���c��i���=@�[�NxfS�y񅛛[�GkӤ7^�z��!@�c���[6^��OP���.��R�}�A�R�^y��j���ٲ�?C��s�Ml��n@B�ۀ:�F�7�t�;|V�kJ��m$"��#�yX��g�F�-�0�Val�{Ll���'-��c�ٵLY�;�wvZ�yr!���K`����^���%�uY�&�U]E�?�<\qm�5
��u���4�DP?iQO�k���ܩU�t�Z�v��]�>���o��vm�X��ߐ(4glaΡ��-�ZQ���:̅�h���rGq��G�j)��A�tѼ�5د\�l	<��C�k�	j姚����0M<�����tZ�׳������G(\��n����A6,t��~�>�t���B���Y�OVm�䝠�H"
֠鍊U���1ol������W���3�Aq,}���u��'��olW�r����_�W)���E�>���^���L1�kn�ǅҡh�:�O֮߹� %��	Z���ϓ( ۚf@�ߨ��+[l{a���tuU��S
�u�_����:�w����]�T�)��g��~�I�Vm��}�Tp隣��A��-L�b�ƃKn�Q�vLaA9�N�g��1ʻ���m��ԑ�|ڿ���3z7���hS}�V��Zd����r�� }nR�w�_A�p$���b|�`R�En����a_Q�#g��[�q�	���)'=�/ý!u:��Ն�y^Fhc��W�0J��4�Z�%�V��[�+s�?�ǒ���j�*ʕ����5=�u*#�4�Hm^V�=N�h\U{�%�/�����Tq}�7{���"
A��f��R����Х���i��g�p��Wwy�d�;��@--.���Q͂DGP�������4�v�9Y�M#�Z�?,�j%⡑VG�]O���6�K��X��"Q����z�?
I��%���w��`��:k��W��5��З�c�M��E�7�z�oc���:Y{.~�O0>��-�rJ�eX��T�tᑕ4�Q���V�8�l^�k�rV��9��o6��V�Fp[Jy�`���B1�&�� x�f� QשRW�{�`�)S��eaa�5^d�Ah,.L��K���[�kl�P聮�����-�h	+B�����.�������h,�q��),��\=u<���Q�a�~d���v1����X�(ef�n��C<3���޷o�~�c��:��'H8�����-{W����ܧ�TD9�ю�H�S�9��b���{p#��#�߾��f����STt[Ռ��}Z�C�׏;�������\a5%��,�:�D�P��b�ѾU$����g ���=x�{��d���r�pl��{�c.���tV��ݲ�
 �(�k�Z^��`.'m��QfCr�z�e�?s$֡���t+�KU�i��P��jy���Q��M#���5ŮL-���~_��W�ɔ5Z�,�7/�J����m�vҘ)�?D�m"�L:��˭Q��ZB�<��L�i���;FE1����ki� ����8bִ����m�2#y9�v�z�+�/�E���ʪ=���?�J,�FЌ��[� &[��ct�Ϲ�2K��'Q²G�49��,�5T^��@�Qۼ. ܶ����Fr���y�D-��?� ����
⠑�3q��	���$a���l�M: �yex��`H�E� l�XB���
�:4u�*��g�c"�C$�[9�^o�J�p�����)X��+
&NK�T?��%��{���&:�ڒ>�v��&��>�8���le��p�R7�Q]��&�;S�>͍aћ:��Ʊ�W.��bs�[]8T�����*�A��H���8� �Oj�u(s����������ߊ�k��� ٠]���ğ�p�r��׳�lfa���%_�l�����h��r��n��z+8�W\B�������\Ϧ������5s��);��Ɣ��Q�W��r�@��Xr�sjE�l���C�ޠ�=��^�g��B��������_}�����	�6.��¬I1�R7�wL��#�ZA{��|*<!2i�g����P����G�YF^SY�po'y��xDq��u���?! ��t����KH��+�D�*��1��nm�Ŕ���㾤G=��#n����ٿ��*��{��$m
OG�o���
&:{�͢L�]7]6��@��2O�H��UF&����Ό�oӥ��:�%	�K�Dۯ���Xb��w>j�ARr��sfr���^>��V;��0QT/]��2Ed���E�s�� �boU�ѷ.19.�A5x���9�iq�u�8�%w���U�}�%�>�m\+����Q-ڐ@�apt�Z()R����$n�����#�t��ĩ�\�p~�e��ƕy6&'ǵ�2���1ĮPh�*��������t��ah�`Vh��S��0�S�ֹ�O�y8�f�V:�\�u���+}���^���B��9�具��G��Y[�}Q����A�D�S�<"�����kd���o�� �|$x���3W~��Zh��Zȇ���Ӎ���U	���-X�K�\e�^{�
�'R�w�]�Yf��a�wg��	j2��{1�2M�Vg�"U���5F&��@RS,5/��)а���O O���4ml|��VA��V'�9~�Y�N,��%�\;W�8��'Z����i׶b���ɱ@zNT@�}2�G�|7�(��Ų����^��*�WB
����#-�+8��/*$�=�ώ�N78P�9���7��j��Y_�.q�4zzTϲSZZ��,�`5�A㕉�jj��-+m0�%�4-��t�1��[޾"*��������a����>�f�>�0z&DA��u�/&��O�BSL���~��`e�o��s��5���ӄ�a�2��w\�<&��P�M��&0�&a}R�WtC��J7�����nm�;i5�۹ZW���Udb�m9�~e[m4I�;)��ϯ��s��+P�L���(w�oћ�k4���B��!.� � '@h�:ᰧ%I@�Am!	�uAK����2g��7Ϗ{��U�� ����]*�n�C6�<KY�U��Es�<N��mT��gcϏj,����(�<4RĪ��U�؇-OlW����-�	AY�(�`���Zz�Wȃ�e�q'�� ���ǿC,���i������	@B�T-�Z^w�t\�~�8�%�6��ҭ��q���e�]|�h֖�k�9�_��qef��yӀ@ hMDpI�3�y_Tbq
������n�q�ӝ���_Fɳs�sO}�%07W�~�ma��\;ޯw�^Jv��bp��YEG����
�q�i@�_���y��a6�|�/��- :"4~�����K/�dP���|"![�i%�j�i����|C�*_El<�ۏ�9(�V9E�u8)�څ�*�Vńz�C��Q��&R�O��X��fT!f�	'B��p�r@���T�Y��Ԛ{߄f�}�62���i�Q{�z�������y�����}��v��P�j+�Qv�Zޞ][W�����"\a�r����y5y���\�4&�K#!�L���������6j�?$9��S|�O�a�]���D�icC�ݞ9��ƣ)���ݲ���sc�&���<>�L��߄�M��SÊ�J�D�A7�M��nj�@���a�ɧ�㨧7��ai��[�o�U*t���\ .��Q�x�����u�V ��U��7�}��<�QHL�I�%?X�d�W���Uω����F3\S"l�x3� i�䜑yh�n��<e�T�f6x�����[(� �z.�xkq�7�,49N���S((.��2����y�{TA�a�R�;T�d��g���)tw�n�a���A�1&w]:�n�s��{����.�I��DS�tk���8w��i>KZn�]X������];��n�L�Yvb�oO��n_����˓��J�Fld���M����4�$��of��kZ�S��!�ݱpL�EA��}�<�C�`�?�Eg�r-(�Q�|�n����ڐ9��"!��ӿ�U&�هēg?mW��ݝ~'�!>�"��LߪW�B��-�&�ert��Z��Y ��Xn�<�@q�?A'�1�Z4��9�����n�h9rg��Ɉ�0������PA��B�wI%D-��V��_vꦊM���Vu�ϫ7�O"�g�K�����ޮ#�p޵���/�|��E�)Yn�Ώƭ��S"Z�Gڣ0=��<�V����:ϯh�e���R��h��F�3�x�lm��5���~�|�)H���a����F���_����w����Q�{E�z�8_��*~!I�zb--��0G����I*��Thx�r<��{���y�z�А�o��M��rM�u���ʚ�z)�p�`�(��w������D���3 l3��?�iA?�){X�R� �#��G+�U���O�����~b�:�A�tf�.PD�E���o~/q˄b�����Q+��O*�b�����zC�!B솖�riIn����!-;�����mg k=��3v	f�k�4��=���iQ��'.t�*�"⬛��:�;��u���pp���9~ж{�<f��ן�����cy�~������!lȐ���9gL��hBk����W��qE@
��J�-$D�\lKp��2zY^�JO���N�k�f�Z@�v�\G�Fs�Ic-�����p�j�9~i�}~��3�i�Ԝ���t[۟ж��KX
�Y��HG~x��ч��tond[�8��%bF��*"�b�ߟ�e��ަ������&%������L(Ru�0�+,�)�� }�P?Y'4��٧po\�: ��>J�s��·��p?��'qƂ�I�nQ�	��9s��p�W��8��[���./Vcmz|}o�r�����i+-��h�6�J��s5]�J\��z�K،����F	���u��	f��wn����ӓW��0�j�0d��!a�W�G��,������_�,W��OG�a�N��̷�z{O�no��#g[d�Z����d=�oBa�0�������y���ÌqB�/�X���F��ڳ�t�>m`�.7�u����6@W�8�v���c�z��L�=��~Ŝt�Ʊ�ҔE���_F�Z�׆��cf!&?��\	Ӂ	� ����N�������.{\f/���3��]�"��X[�Ғ�̓,@��I�̦[�c���e$�x�� �5?�,� O�m�	{S#m.M� �A����������dn��6d�*�6JQfR����`Μ[	���2|d���%؛#�i�ÀN�6���WI�^�<�}3�Rʏ�qr��NA���y������L"�k([���<<�#Uh�Ȍ����n�)�
�bjLxQ8fc��Cx��1:�"��N��ȣ0u���U댑�t)bk��z�^9>N�/|�yD�Y��зܭ��p��'��]ja]��G�R|�o�2��Q;�&ը	{E`}+SK�&B�OX4QR�<��J�o�sx��H9ǿ�vʓ�?#����At�hU��]�L�y4�f'i�]��T 	KS؇�D��$Wy��#�A�3����W���}I��I�k�x�]���=�����'5�Z1t�D��E��Ѐ�uS��!��Q�V����;�d����=S}����U�Q�[%6'���Z��I�j�vӠ��zɕ{���L���'h��&dG1VIp�}��Z,�៊���q�ܘ��-_�A�|��n�Y֎�9���N:��"3�+OV�ΘKz�rpjB�2E�)Ix==�=���Z���1�n���1� Lw�$����ʗvţ!<c����5u��f|��-x��hb���-�hR��5sS��ϟ���~Mt��������;쵀9��:�ļC��F���s3�sϳ���壾�V-L�&�7P\"��������	 ���-U|��,f��x��ʲ ?3�YA�DF_��cCNh�J͠b:��>ku}�!����7��3ϻrJɥY���C���'9n�72�yNk�z���"��M2jO1��17�S���a����\����?�<}��s����\����g�����	
D5;q�d��N��Q�0��E�_�=� �[1��N�c[���!崫>7�VXXj�=�9�-��p�E�dԍ�`#��2?Ü��<�m����P#�.�׹'�.�Q��l�!�FF`���.0��X�
G�dϨ��i��Q��� /��8Hi�Aݯ�<���k>Wpv�A��_�_)��b�M�����\_��_[��}�-�|ě�_�b�U%cjj& ���DJ)��kÐ/:��3�8^��W��t��/|�H9sTr�Ats�x�E��ZJX���"&s�~#Op��]�Úny�Ҥ/��=:�#�!C�a�����B�޽��.r�q�T��x�~8�1�*�Z[�ٯ�.���)�8�0�~��D�B=�9F����
�5��	iė�bt��K��*n�`�6�h��d�(' �cy3�l��[��*�M�{y�k�r��:�� �w�� F�S�Y2��e�O@�.����C>t�8����X����B�d^��{�N�<*��Y ܷ�?��$yp?ɥ+O��������#�o4R��^�_��#0�h0o��Ȕ�)ii�R���L�_��s*�v���y������H�l�xB޵��n;U�l ﰮp�6�#!H�g*�D���(��q ��HL�� ��ѯhq
�T$5�Rd����;Ԋ,"MO@A��N��i	U� עm��@tX$	s�/��
��'~����PW'(�'3��&�OY.SL .\j���uf,dc�u���|!���z?By�>�z�jx�0�ON���y��2;}���ʒI�&Q��i=R��b��ڐ�"��ٴ��+;�ժh��xl��m�^�[<�Q���FF��A��ǄyY��&p���e���-���6n4M�HI�����7�� ��	���9D���\m��Ց��5 �9�+l�
k�w7 x`�Ǽ���1g�h? Q-�ر�[,��r�������ʡ68�C�#�\�񟈄��\צ���?����W,�0�/��XG�48tS,�i�,~��0{��6�sU��^�u�=Ov�,Đ4O����]@M�����=hSs~�����D�A���`2w��G����Y�aNs��|ɛ/�i�"`����Q�0lx�;�\��zD ʩ]�0��8�<0�Uz�é��]�/��;�2���!'<�BʯQᑹ�j�C������\XZ�|Ϟ[��嵲2Y&CӨ3D#��^��F=�R�s:)���ʲ:��CȜ�m��	��Fq�Y������ ��$|6)7���SL��`x� �
>�e�:{���A�L*��9���}�=L;s<�ؒFŭw%ˏ/� �C����/=���J�O�ވ]��'IEsF��H.��{qe,���ba��br�v��zb�+S�R��c�9`_���6؇�H7�q�	�v��h\���w1`P���,�oxaT�����pn��w�=�.JטoR-�\�?�1���*����K�9b �dP'A��t�ĀE/���|e��z���Ǧ�i�:��i���e�G:��1��>���=��vL��4�URz��q0�4�%Za.�����=��kVƓQ4�z�*�L����q�����8�(��Jj�,���v��B��K�^i��7%�%˦�+{�<xv��|��#��qg�D�)�h���K+�:E5�^F�Mu$�A�W%�%j��u[����^#�w��T�D�'�Z�O����@����5Wu��U5��U� ^���L5����G�	evݜ�cm}Uu���TW毈?ᅐ���B�>�n��*�A���/�a3+��J6�<: �Ɇַ��@.G���-� �(��J��b��o/�����+c����Л5	>�������a������x�`<���P�qC��l��/��7�����"Qx 1�*�3
I�r�����F��Y6����x}"Tc����w��u��P�ɶ�Q�'�.z���BB>�Zgg�"W��9I�I������Q*A.��RnՏ�_�ba�PN�
�^�:8��(��� �U�J�����s(n�L�p��

����m98�뛶/�p>Mjm��3�h�>�6Z/���nZFcb�L�Ɓ�&����$b�m�,��fF�<���X��~2���V���׻Mj�pj!�9կ�DC�-4��Wd���KX�� � ��	���G{MO�����2����}���d+�t��E5;�kv��2��RT�+��+�&`������A�!�s�,�N�#�o��� N�f�ڤ��Ɉs��buH�5�o�����a{;]P�����>Zܝċ���.k�m�Ōt)Gs�|>qG-�F�Ք6?�
��y���+�T�|��M}������T�:q=�r!�fM�sf���f�E���2�vU��!����k
d\y��L2��M�,��`�N��Ԗo��y^�f̋1�?4Ĺ�9�|�:}�q(�|�����A@�������%��h[Ĝ�z|�\Z}<o;Ǔ7V�Wi�g~2p8�)P�$C�����ɛ̠��{A���~��c��E5EIu��*zX�rÊa�4���E��[�;�m�ׇ��ݕ�;X���* �hy���as���	�[�c�G�W�`�jo�7/I�������S8�h?��k���qwqI��Tv�ڌ7��CYD�͖�Ww[D� �3��e<�l P���
�t��z��`�i�f�[3S�UnJm�[��/?��̚�C�O�6���+�<��+��X�aU�N�!�1"�7vm�cp�U(�77�_]<$��[���diQ���!I�:���a�j��-,�4 ի�D^TZ��&k��n���<�tem{�Q�FgB"q������|�����p#xf�5��5{�CTJ7�e_��F���|W��$GL.<*���E���:^ �P���dOJ
�:�h玅�������Y�0(��vB{���M�k@�r���]�Y�E;��x��X~�x>l�GC�����ڇ�vڭ����Q�E_��coVa�fy6���1=�f�ۍg���CE�W1��1��L�.J���W�?���h��:@E�%�d�(��m �1l���7���{INl�L���g>-���|���kw��K�]�Qb�i)X�Q�f�:��)���й��|�a���,*<S�IvP��vQ33�6����pn����vhj�3`	�b��|ׁ,ks5�?6�Ӄ䌇p� gh���-!�A�QT��e���<ꌨεO���R���h� �����ڟR}�np�آ6�<���͎�g�����d��S�qwG��N�,¼�AQP�{=[�>+�,f��v�x�<��]�!��u��IIIs1��%�1l.�%����
"W�>R����Q���㸙vQ٩�����)�KP�Wѿ��'	��C4C�a��9���D\%/oV��|��:[3ē�lv�nbkn=SMʴ�&Sm����:�τ-ǂn�$u0�Ħl("Ϗ a���9��)��
V�R�.U�3>w.��{"	��!"P5G��dAiR��|U=M�Xh6rQ�gy� 0�\��B�~��LGeCpW��lY�	']��>�^E��W�)7`:H��	wʂ��Dl4�ۜ'�mهd�Uo�"��/fr(�N��G�ؚ4����b������<A�^@�(�}���'*|�a�ݭ��69�k� ����+��aP�Z֥ꈜ��יw`���|SD�h}e��6 ��z�ѵUz#�Q94!�����? ���և@����fz�����F���w��Q�|�(��S��u�d��_���3�1�(c]�v�L��Td&P*�:RI����<ʸ>��ol�����G�t�I��)Fn�ǔ���� =zQN6RY�M��^��:	 �Zp..�}]���5*�X1�	���6�ǲ��Nc��q�QkRW��Ȯ�3y���8m�����"����
��\&����bEԺ��
�9I1�y�'b􅭰��SF�l@������Q�Ev�җ�v&��e��@�����؟�ab$L�o�jS��x8����H���������W���8�	_q���tz�ϖoY��
j-��A�w5H�R
M�Ҷ������+X|G����~��߀��[J�J�
1{<��|�Y�`Y*�����`��X
�-�:���"���l�~�cA�p"�]3x�M��:��V~ZqhS�T����� �f���J;�K���B��=���4�'+�^�gr�]���v����jUiB?���[/l�3װ�]v�^�66.�n�:=��OJsV���YM��
���N0���E�F
Y��~�Zf�����4W4M�����ؽ ��C��&!'It�����դ�Y:�����>��udR
H�Q[���{fe��"��z�cqD�N� �(�W8��U_Ԍ"�b^7�">gq/�QG�><Ծ���>y��L���ֱ�3 ��R�D�e5���=��d��u�b���|A{z�uGR�4��� �_�}��*ls9�31ˌSX�~>zSi���)�&���g';����#L69�ϸ�A�B؝B8��%�a�4��Q;{<]�o�Ȗ��6�<�Ȩ���sF�j�2b��?��L�+��ww~SyC��I,�#Sj�ѭq��/�wS�DG2�V��#�%��x�e�������'�N��~^<����:��	i=.[5,&�w��xnz��{j���R�L��Ԇ�k��L�ip���Vv\|��!s����M�为�H酨`��s��NdT�&hx�YY:��0�pg.��v��h��]O7��^��~���ܰ�Vwê�k)��`�D{����8P��!0��N��'����h���e��"z�)�D�0����0�h��穯 ��m5[��%���ƅaH^G� }����茳�PI(��8$�v��g��������ݾ��&�LQ�*�����*�՛P�����.�F�L�Z=,�d��k���s|�r��x�K�4"���PA�f�9����tǬ"����.}A��S��Q�=v^�>ԞԠ��YS�x�A��øb���Y���%UU�忮�=Ү1O��� �����:����~�|=g�&̽јh��WK����^���Ƕ��E;��.$����^�I�d�$?���J#σ-¹��;\�]3�����+��K��$�z��*-��uJ2��ayo�~�]j�Dnl)�Wh#f|���H9JS �g���8�:9���*Z�%�7��8���!8�c��å�pߩ�W���+��~WK�#d����C~a��x��nq/drk�P0��vw(f�3� fY!D�2DB�
��n���]�2�jQ��N�F�`���i�! ��P��s�952�6��9�)U�@�n�j�%˭�cϯ�"��V�q������R4X�$pឪ���{��Ղ�>��@� �]oW���U�q T�L�i0gb��0��C��=��@>�EhjBGl��R�>EzrN)}��7�*I	\���͎��X�qI��v@)�r�Pׁ�ٓ�y����$��J����W"����2��g�J��SI�6йČ�6X�$���l���'�����$k�In��\顮{kF�,ҧ<�hzۯDpL8_��T�Zw(4L�{CL+�\�S5���6aK�t/���l���׳q��J�ϧe��5���0�澴A��# ����g��a���@^xV���赡���P��-�5<��pq�I�Ͷ�,�Uz���9<C��{��]@��9���'���hg���n��8Fn{m44,��:��P�Z����l"��>��4�?����ŷ�O�}Z���T�B*��<$���kf�#��t�g8^21�9��MD�Ҭ]>�ɼ�^T��Z�q*�"��!�?$I����[�����$�j#���1�J��a���8�=���,P_�K����c��ȟbL�º-5�"���I�Π�v�����C��C�Bh����k1�t�t`ol�]�ʎ�t
��X�-w�@廝���`߸-�{������ U�ނ"�o$y��C��kd��*�4l�Z�Lv�m���e�̜Z��R�#8Є,B��g���*P��E �e��A��?M�i�Ą>�-U�U̅S�N�V�
q7�m�2���=��&���K�#�v	V?Wc�b�Y��b��̯�b����"L�cڡ2K5^ȩ��y֣�q!
�C�Z�h�-r�K��x��P�5;�%$�g�<� S67��_�����cq�N�}E�J�?G瀒��A���C�^�
��޷�4��{�O�C̭i�=�^VZ*k�(J|Z��� ��&LA���	՘j>���S7���o�p��G�ѕS���l�a�` Sq�g�$Gn�m5��B ��hYQ��ٜ������I1/�̖E�0�FLӡ���G��a��?]����t��*�L���Vf3�e!b�»�����y}*�X�O'k�.�+w����n��Ya>s���v��R�7S)�-��N!`),��H�š��P���������v����82s�@2�Hpg�6�ԛ��`0�2�g2A��ժ�#w�zk�+��+��ׅ��gA��ۄ��-ll������4'�9NK5�P-�Di��&�3���]��5w�W���
P��?j��Z
��E�rcu��<k=Bf����B��Y4�V꿍3/���N3���O�T���u�5o]���T�b3.��y��k�l�c���d���q
��C(�$�p�]N9S��@���f�C%�U���薦c�8�z픯ڇ��:���F������9�ZG]�r��3e�{���iq�tý�U%�	�c�0����b+#(0�5M����-�z���FU�?V��>s��eh�=A��o�vH�&u�,��k�4�k� !F�A� &a��߇�蜷,J1B�=*���B�IԘPP�����@H�5]Ky)k�8v%�bQ��޿%�sbX�I0It0��K������mo����������\��:�C���{��H��h�1��{9����>�;���Jp	��d̵g;��{�?�����@)V�_��)�����z�ȡpTǠ�*a!S�#�FC���Ħq��{z��Ք	$Ў��'��A��?���}f�b�7�\�
�CD�d���*6A�8��@����jX=g�mGS_���3"C�\����EOt��G6�p���/��a�SG��>W��eϘ�c)�R�K_�KZ�T�|`y��٘���	 玾>N׃S����5IMk!lv���k~�|�p��x(/�h�՜%�x��z�J���~q{���-�QF�@^uv�u�>^�x0r�k`�8	O=��;S�~Oּ��kp��dAoj�b�����:��D�
Nr6Tr|k��s��r"![��R��>�VDE��P��pX)�7W<<C��"�Ԥ����� �xR��Y�jl]��N@{������->���6|�9F��xq^v��~�������3v�����}�)��R��?��������Η��G����ҋ��ch ��b�zV�M��Z�F����4�W��!l�[V�7O����b5S��98��}�������c�c�яX������E�㤈��/�{�GݫF|����^f�FrE�� t-�p��A�|�@4��X��[h)r�� ���kR8�#ڼ׌���k=RNi�I�Y)�R9���i�0��z.4x���Gg	�p��)�-�ػ�?k�=4ea�{����NQ>K*�J�����"f�6(zQ�2˸t)��8?V�ܚm�!1%��3m(�]Tt���ܚ]T,�/5��0"�a�;l�
���́�.G�Q5�"	��=�8�y1P�����Wڭ�#@���=��X1�hA��#�k�i#�� �)�N\��a>��Bt���[���Yrq,hFh�W�Uupu��r��JVh��{�����v�\Gס'��'2kp�=���.=y�Bh�5MV�>2�o��,0\�oXF�{�n4>��Nn`�]iq���`�sh-]8Ph��v{`Xؽ?���t������!�$h�����\�sǖF���R�������k�K&+/�B>*h�.�T(=l{���$$���c����8�`��V�(<�x�tx��/���my�r���4���]�_�9x2��n��Y���,+��N`u�e� ��X�f��uHN�e�b�عD����I+L~ ��hy8�(=46ɸiy�\�������m}:5����R�A��������N}��N1Az4��MO���`;n����}ѭ-�+��N�4�gw�91�w���7�+�J��lb�S�Z-��H���y����.!*:��8�����M�}�Ҋ��hj��O���X����(=���ĔG}���M���8D��Y@�ϧcQ�<�>h!�:�Ή�;��dʵԍ�߅ ��Dְ�O�t�X]~S����h���t��b��z!̤�Z��0�Q�bP�n�'���0q����)w�
�h��E̐8W_ަ6�������o��P���(�c�WC�7A���g��x����ᓆ�h���O)6T���|�*e���� h:�Zj�ac$6,L�Z��$�0ݻF�9rK"�WN$��Sj�4�K*����-���h����5�̯Bn��KR���3��o����L=M;��������!H�!i�l��u������B�Y����F�~���4:r��᭞����I���f����TRL�z��J�B��] �:�����룦@�BNm��M@-��I]�h�b���d�	ܹ~9.U(��m�,�i���+�2rcdhW��%+G@x!Z��(�h=�Ƹ$浸G�T�}�@#��U��4����q��D�����r��_�9U��HXbJ|���.+�����No��#K�}��x!T����.+_��ea��S�5�z����莀�"�` p���z���~�;�q(Z3��1���:�hO���r&�h7�27P�E�Π\��q[F4�%��Qf�<����w��d��|��u�G���T`{�2;&�[����l�a���@Z��w��B���IT�օ�yd����J�)���?�����Iz�v	�#:��Yg�Ck�d�8OX�r9tXr>d汔�{t�>z�&fq]]��)�~������W=���pjB�����8�7G���{��XC*��TT,âsk�I���Nr_G
��@���^)L����)�;��]�B���_ڒg`��h���X�P���?m���iݸ�����L�pʾ��a����I#�D����Xt!�n,�|r�ep�|��*���di��_�P� �����~]���ǡa#[q�� �)5�ŀ0@U'}��*;�=�A�{��=	#*o�@IJ�O`k2D#���gus6����jB*��U�����*�2����;��ms̗�=r��C5�����3�N�����r���&�ܙ����.�:_
�s�z�ؠLOﰐ;��aY	�(���zn�1U��fJtB@��]�`Я	8���v�[�~͘���H��ҹ���w���5� `�����|���I䪔D>%���1�3���%�ꞬM�;�3��}��	%��E�Cl���<ĳ;F0��<'����@=�e�z�\���z��
r|bEvk��춀2��/9��%�&��
��m�:�Noc�/.��
����5�"n�?e �(|J-$o���k�]�V ��;(���:�FV�f>�)��Z>E�G(~�cp��%��*{���^|�� (Ҩ���θ@�������peGچ�{�;_�՚�r��?n�� W]n�w��q361{yY�&#�$h���64���ɎtMujR��o#Vg럑��JZ	7���[L��� ���Ӓ�T�'�؆m}���R]�s-1�i�pb�v�Ӹ�6��9
���Y^�C��{�,zl.�C����HT�\9t�ޔW>O5��b�;-�+lnO��ߦaS��-6�xW�oa~9��3V,٭���7艻�$�"�R�G��G��5��#���X�}�T�u:�.�ʉ�Šx���,}E�}M6qM̼����Q�=o�1Y�l�sy� ��HW+�]�������~ �����6��d@�2�BK��rBs�:~.RL�+vX���,go�Y̫�{�F�X�%:Jz�_�*u0�kX���)����C�`������V��<.��������^�8�dE56�/��g�P�qv>42p�7�tzy��Nq�0�P0"�J��*�#��0�`A�Z{�ȱÈ�s�ɛ������� � �z�
y���exR�*U;��2����@s��>F���k�㈳l�gB�����6SJR%Nj�8�,=I�6o_-�U�� ��^A����� ��1}o�68&LH��lE�,<-��>��7|�E��$Os�W�87�����n���i�a��8:ŀ]$�Oq�]�fvCEb� gA۽uj��Wg2Q�Z�ˋ�P%ş%-t�e Vw�����E�T�Y�4H����p
M�R�����	C_��/0�슡o0�5�p7����%i����l�aCa�Ò[�28��B�ST5}����j������� ��pw^9c���d��M���W����:��e�Ã��\"�M�Ƒ$n(�m�*z�d4�t��$�����v��/���6��ԙ�!�%�:�3d�_�z���x��f�uo}�,�}q��}��@����W�x��[��$��c�vCp�3��6ul�Xq���|�e|���i��M�?@g@�^�%���e4�ES��]E;z�{����n7'�%�`Dp~�+�������{��I��OIT��E\_<SrE����*�>��x���@u�თƝd϶�[�����w�}�u��"6S_�tm���Z��=P�w�7  ]p?�k]���3�!!%>@|�����T�M�ł��$ TP�ӍY$M[�՚\�m'cwP�,�����s������5�	�
F:+�.x~��u3��Ɗ+�(���� Ʒ�d��s�k���Yzr��m�	Q)w5jǏ�p�ELK�E��K�ER�*]`O��"�0�L��0��D5��V]� �I!\�!4!��v:�D�K�7M����׽`��qd��������Ʈ� kQ�w�tt�L��w3�Y�T�s^��v?� q�(�`m,���sf�{�7�]	�liey������B"��ّ� -�k�<��(�- �Nq�0�,~�@�_Ķ�JϦ3�)?�,���IP�*NP7��p�F�NY�g���1ȜE��Э?jP�� ����|��Q���j�5�mk�,ܓw��?��D�wOe�9�)ك;Z�s��ܖe�����4��Ĥ��-ؐ�D��'�����������L��Q��uv�=�n��0�W������R���|x>�/$警����|�����D�YO��dzs��.$mn�\��<�Ҭ��F�F+î�t2�O~A3����ɱ�� ��|*����]\�x^����&�)�^��̎C�Ȧ8
�f�����%�e�۽�]\u��Nk(�iqe��e���gLb�T	�����l'#�h0U3��P�Lwq�b)=���s�6fy�pږK���!ו�Cz�4�vP��3�b��T��x��eb�𽕦����s���6���2�U`��}%	Ujn�'���U���sh�.m�x���SҐ�k�>��?k��/,<f���za�rB�Ro�-��˂���/�����my������N��L
ۡ�qo�<
�Zkz��{����n �X��ʢ�������5Or�.������L�;m�P� T{2K�{2�C~�,�OvMyȱ��4�7B$�R�0`,-&�h�[�V�� �s���	�t���e�ʻT^��qn:�Fq�U.�F�g��"@t��(�%7��b���f�b���J��')�}B�]�p���L�������A�z�_��� �Rab줱�0�B*9���;��C�nF��Vc�����M)#���Y/*�
3\������>���9ߍ�Fb�z�%�n�ȕ��d��!�8`Cc
Jg5�1˅c�R.�|��S����X�:�+8t�̹/�[��b��,�g�џ=		[�m;��/��<?1P1�S��P��N����l�X�?�f��m��I�	��@�}���/���焘إ*��v��O+p(-,çy9������/"�-�OR��`I�9+� bo"}����S�<��V�
5Y	(���,�+����r�������~���Q���&J�+lx���_J�-ufc��N�v���@��[�c`����t�t4;�[�<�gP�~���zq�Cn���}O6��͛2�8⢎%4�X�L�]�F���NYU�����9��kr]u�_>{4��<l��� �3��s(�JV��R�d_���W�Fn=�yy C7�y��	�a_�Q��>\����s1�����TޫΥ����;�Z��T%b�d����`�m�!0pײ��lٺVK�jYf#�G�"��`��tc7�((ֽE��f���d��=GE��S{��)�C��N�ʇ���(��'΋C&{ѻx>DC��mf��5�����͛������(�̣}M��F��o�KKL~�Y��q&�h��	� o�:u��x?���ww�54�M�	L�1��L��ȕ(�����}�s���%a&��X4:q�R�S����;��	�X��cO:	 Œ���E�Ý
%�J�لB�&�ƆYT�Y[�p�*� �.2��d�vEI0�dp_��(�9NB���W�CvOU}���e[E����A�� ?ůw+J�D��$e����[s��!�⠹��6�iKa&�~��/e��Q[:��eb�2���;�'�@~���N��U�%��H�x�K/]�WC��sp
�+>Hd�':F��|*|�50ϱ\ '��]������O�	2Tc��u��6=c��nZ#7�%V�Z��Շotyk�x�.�Yń��-�(Ќ�����1�^��KĚ�q�2��+�|i����$j`�@�$%��=�y'�辊�9�����{c�m�6~Q�'\�IG+nx� �j�+�s�"�Fl?0v�S~W�f3�v%�ӊ��I����/�J4��Q���t��qD[+�����?q�;�mo���ʜ$� �{�#�Ҷ�$�|�`�ϡ�H�}��1�KT��dn��O�-�:����l�0P������1��M�!q�M�>�ے�b"�Rⲧ���e�/�ח�
7i�C>w�
�:�ڊ�(�\�~���p!K,����%�-˹i�ʒ���7��%�)���Igu���������Q�٩K1z�����|�U�H�ݮ�ˬ��ͨo%z��\5}�Ұ?��?��b�d%{���9��&�6̹��uI��]a]�]{��f�QH����հ�1k�JS�Y����7�:�]�����'c.{�Lֶ�^FGt����L���ղ�Gς�=��6��x�֍wD�����%���qr��"�ҽ�G��뎛�ђ	�'�SR������O�����0�T�h��'%�C�z �U�%����sW�iTT.Uk�*�}�uS~���ߣK�y�KzX������$�N��F���C�o���2�-�0L�6y1�I���\��~�¨O��fٚ��A���]���f�I�e� F���kn
3�]A#��L�d�-�z	8&�R�w#i�Q+��p�{�Hu��nu!<[?mT�����6M��_|�w-��L���Y�ʦLp�`�i^�;&�JΓ�05�}U��4��搵u��Jp�lCұ�Pse�u{��6P�<��0Ad)�ޝo�s�ǁ�=�ڱ�޸g���сd��^8��pbk�;�as�ű�xQE��T�k%@+�|nIҸ���[����U��Z��ˋ���~rh�5�'C�_R���K��)xZ�ּ�Y�%�ؽ�M�N�� ���l��I��6q���������1������ �u�E����x`g��bt�g&�B-�w�J�g��:L��:o�?�[d╹˨j`+Eݥ����~���}�8t���� ��Nu!%�(����j�J��2S
t��s\XQ��$O^|��=)1�A�8Ʃ"i�bMԧ��9y��Tq����g#��4c�$���з�,�Q�!.���wc�z�y57��X����߭���N�v��"�fo��l���. ��>�,Y�(���5�h��a���b%�~F�\��X�X�ܥ��4���#���1tCl��}�"^�^��8��_S�tѯB�×�=f�};�{�\=�&N�B� �rT��;���򻥱P���[�Ƽ0:��m���鑀�|��ᙴm-��,mV�o>�;���?�u�-7���$�134"���|\9zk�n;B�g����Ӏ��"C!�7��i��*[�+��F�G�IGG��>�ͪ���wK<��]&���ߩ3�cwb���`�$�ǆS��Y3�d�Q˟rF$ �YǓ�4s�Z����ia���+��3�2	�4�/�]ź~���i36�\��J����t~�ퟳ�R�ܖՆd'�<��y|�#�9v�Ѳ�}f��_Lmp���P��4�m��:w�f�E�wxt��XOw��*����9;&�M{����C>�ҁ���HEdV`��"1��aDG %ð/���NQ?U�t���xC+�h�4o�y�1u�3�i�a�W���q�)������[qu����P� 3�m�Ӻ���ٮ���	�@˃��w�5}��G1X��8��L��|�+]�6��O��P7sא�K�����@Y�tx�Y/8�8l��?�'%(�z7��%��sZ|�S�0�a@����S���"�j�`��t���^���a�:tCdc�>����Q����M*Zih4==�c��5Un���P�e2�ʹC|`�u�$���:(z�˄����'y��v��рd�#�V��:)���	7s-p"Y����"t;P�=��W�9rF��!�%NlX�c�Ɛ"�'k�1O�//���^��Jy�ߨ`~�I���*�	�?��2��ԟi�LP���Ɗ�X\@.C��r�����m�E$戁���ycx	W�����I@ ux_n�/#��^�Aðv[$�)Jm<S�`���b��UJ [�(�	"@)��Wq��I��#�Q�Q�dv�,�]'5�����`w2l�_�N�ìQ�p9�D̦P`�즫���YU6�Ca+$�i��щ�1|Fz�=��]�?���r��8�}��ٺ󋁮A��~�Uef���I�2o�k�4="�01�_`!H\p�I>u�vZG3�x�Ez�g��P*v[�=ow��ѩ�"�X�F����A�� �_�E	���F�1��L��O� ��@c��6i�C�a�h8*��h�Kc9ρ�JGˏ���{p[��7	��&u(�� ���Ҧ)���H~�J<��Ӧ�8<L����H��=�yMF�]�P&N��[BF$o�ٺ�^�z��F
��0{���cfp�r"2v��t��$�!>����d��M;8�3�g�7���W�f
U`ELw�ld�6�
S�h�>q�>m%�$K{��JD}F��g���o\SnG�/�	�^+l�� rb^pz�b5&��w�Q)D���=.��8٠��c�l�ԛLT��51,H4&�oz�֊��*0.Ջ+�䃄��#���N�����A�w_���&�����ր�~*����h�"��0?Êhj�kc�SttK4��-`'�O�@_���C}�%ODu��g�-I�\�D�N�ގ7A��Y�CE�����y�ݼZ^����S���G��������t�-�;#^���|�n���^p�2�z���j��>�[���p�����0�Vq�L���ݬ'�k���"Yxf PF�?�aB�#���{giy�݊F�58�Bf�;�hP�>��Bd�U��x3�Y����mƙ�ٱ�-s��C���P����b.{�̤��fK��o#3�Δo`³��[h1����q�4�q�袊�b���/tI.�\�r#ٴNl�( ��]}��le@>TGQ��xJ � �z���|�ƙ/d)P��7��CJ�6-��.�ξC%�<�OIB��YBX2�]{�#PT\>=cZ����e��狼�:��E`����*����*s�d��9ۜԅ��(�S�N3�֎��f��.p����k4��<��u�}0ovc�T�/e�
��OB=F�vhzj�B>��Y�=�v�?S9����S��5A*�4�d4@�+e���O������b.T�21���O[�B����á"�;�+?�@�^n5=��/���jV߳�17^��	&U1����v����	�~=���\ 8���;;[^Q�\��ܦz��BM5��Z�\ɾ��Yt��2%vWgr޸W�O����(�t,�(���&��/�AV�-��c�;��/-�9|���%��9Ȗ��K �˛�2����5�B����z��ʂQm�����pn�����|��I�3C�7A���aRL�ş���������%j]��+<`F�o<�f�V��"H����4>@?����3�<�z�����(3�ҁp�1~�պ�𺿯-.����d;�b�3�T92!|�PE	�خ�C�0��d͖�ZNe����4��y�M<�}w�Y�)a�*ӛr�/��S�وg�Ϻ����2cҝ�Y���*��
'㼕��3���*STq�����ՙ/��|,Ve�W�ޗ�{����G<���@HbB�C厌W(�ؽ�9���C(M���J�Dde��b�JV�����a�M@�.|�^"~��A_Ŏ	�ĕP����%Qʃ�z|���'Jۄ ��Up6j!7�5\����?����%��Bv������1�]qd���#�^��?�Y��<���p�Q#.e�l�|Y��F��]��4-��2���מ�h�S����kg�&�aBN������,��\s]u�wJ��P�_l!����/K�,���#R�X���pL���R{��߶���^AkFh��<1w������BWQ����P�\����KL��[P��P��ȕ\Y؊0HW�+�K�<]:ԆMQ�+i��irf�|Դ��ɣ6����В��EcH�7sdA��_��ͣp��cE�ϐ������&#0l�-X���ꍌpY�Ox�u_VtĞ�:tU�n�q+/b@�=�%���%cצf1��'G��4���P��*�t�������1aH��ϑ>C�V�bS�e��&�� Q߲/��v���A[?E2~�4o�01�Sp:F9���y�����k�����Kv�	cu�Z�~+_��Sԕ]���ےY�C�]���C@8��䭈�B�� ����H,1�j�j<����,]e@�?���Hk
�n�X�*#w�kl���(HdT�A�ґ���=鮴���ykKV�e$��0�KЍ����}�����B�DJ�o�+Q��O0�z�ԍ�Ś}������)��U�A��ù���la�>��ݺ��B����J��|kHp(ĥ���n�ܨ��W�I����2 vD{[�pd�r��t��6��V����������)vW�Vj��'���@d��\$�30T3Ro�
O�ҳ��G�7--pZ�e`oa�~��$ .>����qt�����p0D�-p c�EH	���<IgNd ��j�8��Xlz���e��(m�8{@d�]q��o��Iy9h:;x����(�[=�Q�Ѧ ���T$p4>����/
�"#����:� k� ��c4�Q}�%f�q|��P����g�	_z�?��\[�_	2) T��9I��!\˻�&�CS����������($D�.ő�uZ���x�>w{��BϫƸV��QY�����oH� k����Ȥ6�GT3������Q*y�^s��'<�pVJ+ۄ�B�{��D�Rޢ�(��1��x&��wN���/~D%��.`��wgѾ�䟜�9P�-.��s�_LGm�d���#��e�'g9vh5��0��<�#�m;(\�4X��:(qvm�x��w�E6؈���b�D��s����F��&��h5��GR1a&��G��� ��wJ�Y`�4��\�a&{H�	M!���c��`o޻�	��a^j���e���xɢ�躱6=oѺS=_���3��X��tڸ��t�q~�B�,�E�����(O�*JQ?J �^���#����B(LW��!�E�?�F?9ǀi0�����E0�J|�f��� ϓ���qc�FVlIe�~��ۉY5J��,��{�l1�GMuPB��8b(=��Jj� %@����\�Wqq�[�gX���t���� ��B���X�7=�kM�^���s��rf�(������,`�1U&u�?�	��x�!�y�^�A�5��R>6_0����Mf����Ozm^
Q��Qn��T0e�4)!t�u�&�vMT�.oM��{Ŧ���U�.Q�=��Ġ5��c�)���vg�gdI�ow`�Y�B���jy%x<BM8E��KR=V�`-���Z���t�� 6�K����59����׸���,��8��4�1�g�
l?o��_�w��z$o+6��=;T':c�2C�H����p�_��f ��~��v���w,�w��2@��U���j�U���V��e�6�n�� �W��%�W���1��l�?3�\o��9D`������F��� k�ix"�6F�ʟRzp��*�(z�1bj��0)��
����4�4p�@��թ�Qb�LK�y/Q	��N�{�FؽQ�$�<�٠]m3i�+z/�
h|� ���n���;�cE�d_['p9D͈���� ��y�P��b��Ǐ�~������!C˚
b���w��o�E��Vv�a~�+C�Bi'1�~?�v������Z�j�7�0)O�c�rp��0̅rڶ������`BO��_�˥�KR�b��h�ſ�M�s>���ɞ�.M�� J$���P���ָ�p�[J%m䒽C\7;�o5➥�*�p�*G���Q�͑�dw��q�Y��s�`�O�B�SwƔJ�k�0�M(�xx��R��s?hBw'E���~r��²����� Ƿ���,>�H�B��!�
˜g�����*v��	7�'�T��l���A�Z�m����k`�z�dp,m�~����˄�x�����2��6M��bB�]z}k�{Z������P����썂D���b��[���Q���wy�zH�/�X�LϹ��_��	����3�1荻�"�z��#�$�G�C��)��X���A4p]p��nLM@�Wp�X���Hi{L"��UK�3�Q�(��?.� )�Ԟ��'���l��as��qD,h4�<f=��Q��w�pR|�+����ݹ�0yhsB^U~�^?���H$&N���5��Kr��h�Vʭ�D��f�$'uAEU�Csv��<K��+��VQ�a=Eށ����A�ѣD�*�AB�6-	�2��cq�}��Է/�3ǂ?k�mky�"��H&�G�?���4��5��ʲ�t�(�-��I��x���Ao����0Sh�VGC�挏��;X'C�n8�:�#�큿b�=��(�ˁK���>E	��1m=ח�B�Ԗ;�)rv(��K��:p�:�:-|"�ǀ��Y(���7�i{����۱ny$������z�5NU��.�\��=![���b�&< 4��Cĉ��_EvJ�s�*�����Wy�8R�\?�2+h[\Ў��?�J���Z ��.h9���l?pm:=�B��/W��/ѡU�����g0!�Ax~o�ȣd6��Lh�[T��D�-D
��?�o�{����۱F
�M�,_.}َo_�[�J��:ރV���*b�Hzm�;�Y$�U���H%h�)���\���S%FC�'�Ÿ�4����72��Y���2[�.@�嫧_�ڪ���������@a�Ś�`51��(����.5��*ݯ�?���X��GW�М^[J��@:>0̺�tNg(�	�r�ғ�Le�sجw]:��Y�9�&�f�։_�ω��~j�X�>��O�U>���$n}y��=�G ϊ��ci+��J��(Xҁ���',�}5mg^�B5�d=���P4nZbAK�D�@�)	r��<�Ѝ}�� ���,iZFG\"����1�L�K�b�)]o���v슳p�L������y��?��4�Q��U	T����_&!�&��WI��諯�?J m ����j�AT�Z-W@<�\�^�Q�I_6��g�;�i�tz����C��_5A]�+���%\vc�n�w��`��j��ޙ�ͤt��74
�%$�g��&t��P�?��ǿ�qy����1���#�MD�
���4=�KS������V�m;\r�W#QUj� ��+|�d"��g�t �G�&��>�+P?���y~ر&'F�%2�n �FW~��>�k̃+����"F]��](p��~å��Li�'�m��W0n����F:ʍ_ޑ����-쪫��,��೬������{nLLHIߴ�pH���IbD�h�����nC�b��`7��������J�����*�v��S���m;)�+~���F3�z�b�O]T\�h��s,0 a�>S�M-y2jt�L�O�p�}Ǔ�NCz�s)h������q�h�����/9�2�=��km�P�PA��e��Lp�����C��8�e�8�5�Zi��Ռ�y�C��P��׿f�����=\�%K͜�%:��d�$��N�tY��tu��c�����zL4����=��b){�gW|}���6�v����P���m&��HC`�a)��*�Y�+A"�i�٣E�'e�B�l�W&u|��3ռ�( �^z� n��'��Z��}-ҁ��=���K!�b�1r�q�B���u^�دdl���ҡ�N��z�� ?{S��`�g�G��Z4��$Ot���!�l�nO���=�2ζ�uHS����s��Փ?�=��p���6gi2@�s�V��3�E�%S�*^�?����;s�Z�f.�� `�Z������8��_���m��u�ʿ2\�6N���;��O&m�~L��z���o���kN~�1v0��3Lb��v����.S-�ߙ �� Dq����iE��P|�w�����N�J�L�0�%v��U'|�]EwZ�Ǟ,}�H)%`4����u��}��E��p�a	�W��h̩;G�ՙ�H�����󭞑Hl�0��Nr��%���c5;�3\R�y�T�1=v�|`�,�]aI- 3xQ�'({-7���f�%of�j<'�|W��V���&�:�%�Ĵ���v���{$�����i^�q.�w��xg��"l[��[9h�H,�G�C��AZ�:������X⋼����iV+<����Hvo���)����q�3�>��.�շ+�W��Q#�klH�m��1IS�A(��ai.1"	��Ֆ�yKՂ��_8S�T<�O��f0t��j�rL�_ ��uay��k�=�h����d��jpe>��ٽk00��-m��ʓ�i�0���̌]>�Ws�sd$O�Lգ����ֳ�!�R��=k.KM�3��sRz�D�%���e����t~8=�� З0�ug5u�r{G�μrd.�~^���:*(� ��߆!��������k�6�&N����7��<��K"�M�[�����������73��!��W��RϠ�&<81� ���lryͱ���^�@��	��Vv���ڹR��c5��m��DT����Q�6�h��"�Q�ߍ��h�
h�)�v�~/-*�N��x�ȧD��V'����w0��q5Պ6�z�,{��)���b�x���jIG���b�ٔ0��뻨#5o�k���#h�c���Yہ̑`g3?�7�=�St�s)q��(|\�򱚝I�%P^4C��GD��D��w�^��$�}�՚���nh}���P��ϧta��+l�����,-U�x�Nl(�M�lM�����&��0��. ��۝�6�/H�I���EG3ܿ�/Tg~1��J�GX�3��gI�b������r���V;���*
i9�g�s��7����3�/:�_Kbc/wcC�b�0�^_����xr�}vR��6�=d����Q\�c��`�W..�gR#MGQI7^`�%$��;�O_t�MI�8#�.:sC��6j�I��ه4�,}��8�90���aLG��Es���N��;���?��V`���8�piL������^c�1R�^<��B"|=r��i5����n����u�N�	��+�`�b���*I�3UE�ةO�oR�"��i������lċ��/�j��ro2�i0�K!�$f�� -�{��i#�wLx��QHa%���e�d��j�x���XX%�7ľ�ɸhU!c>�X"���i�~4�,v����BTYP��v�_أH��x�n�o�T���F岏fx�@+j��[?�m�<6��1�ɋPj�G�x�+�B�1xF���`�ZOEW��ܫ�#f�)j �K�r���1u�ZK�<�:K;��*��~�o�H������#oA����=����g�~7�𥩳NN�z���O��G����HB�_!��%c��ӗ�-lA�T���s% �̌g[dN��E8���B��/���!ĆIkbq� ����b��z�|t\ˎ�#_�d�?M�y���&��q�]�؂a}`�[��l����m�&pnp+��Jg�!����g�zT4�����1��w��ɵ���<�.�џ�h����C )҉��I[�7������A�UɲU�[g=>_�C�(?#(WQ�?��S�/�P?=�v?�ޙ�\�pOZ��O��Z�dl���e�{Mm�GiG�_��r唴QǍ&�!ȆR�4�eW��S���M����y��ZRGh�vV� �aG�f�s���Eg2�#W���d�E�I���&���%�6��6i�yx\�x�F���5D�#�qw���CM(�?�f�iU�ܒΎ�(.� �HAGa8G|R5k�p��[�+�JF����+n��`�����鴚U)y�w�jp�H��Ƶ�\�q�-D�������MvL7���z� �}�����#�j��Uo1_�n���i(��\��+���ū�o�80���d�E�75\��׼*HO�U+��U���P+�ՙjJ5�5g���vaoy�gO4 �CC1�w�o1�G;�@�i��o���J���+V�S��8)i��}d�t�&˕��!�^n��>�� x�<#&�����^I��*��%�oo�G�Zf[�(�Hn"��Y@���p�;��E3���AQME�t�A]�I��)	I�8�ģ�j��93c�w��r[���c3�$��L/=�u+ȉ��yr���D%]"�?� 7QS�C���g/=�>'DCV{��U�oL��e���ۉ���k�S��{@B��N�Tz.����*̙I�~��!��˽��	+vD~M����#`��=����$>2�~�e� �Q@����9O�KD���O��5�����.�`���{9#�X�[����#w��d��/{��*�������#�m�XU�W�=�x`�d����wP5��W�ݱ���۰_�u��KJ�on���؃�a�rǩa%3O�-.Ey��E#�<vy2]��U�M}�l�� ����A�뚖��V��A��������&�ZL��HY��j�w��A󢋲�g�9�آ9�W!
�D+��mx�����4��-I�c�>TĂiZ��$W5IL�d�}
�+���=Z���J*�w&��H���ZJ�*v?:*'ʓv80������]��*0�9Ԭ�6�9ˍ�E���5Eŝ��"�z�1`������͉{¬���pa"؀q�Z��;ɵ֚�VxA��{՘p�I���6F��Tzj�W��kΩ望�	!��CxQ��񬆎k0(��`��qk<l;���Z�>j�OJ��A���(rF��mc���&��x�6fBV�T�_�W���.�zt˚�gK(�)>�ւ1%�@}tt��!"[�h�"}Mȫ�V�ۂ�f��:
�x-��LR�6��Z��F���;�י
�\��1���ڦd���2�s�$g��}���)e��.w��L_uQIJB��y�8~<�HH�QD��z�ɸmM>�8�!N��`�s�a������e���#y2�X:��w�ؓ���Q2�#R�����5�<�N=C=��?7��4)%�������i]:�3�?�%�Il�B�:^NuR�����=�[���h�.l� ϟ�$V���?�{�.U]�l,3��E����?���� {�O��3ţ-�D����(�5|�V��V���ba���^���:�,�� o����[t.d������]5�4#�7��C�):g��E]}��ۋ�Hu�-���W䈗����E�o���"J[0��@nwA���f[��lVm��"�/��G>R8|Vu`$��*ƃ�-�;#	h��V���!T��i�Ԍ�u�?�o"�'p�c�)dPR	 ����E�D�����ead��T+�y`3�!�%7�;�������#���bi���)�IgZz�iܘ�U`}u�E"�%�Js���h��"�&ǷC5��$����M���Y��Q+mֽ�$��x�����Ōg�X���3�_,	aƳ[l�"�{FD�q�g�ӊ��3?�G�̋UP%{�`����FM�c�GxA���s���	臭&K�l�a")]5l^H�2$��ᶴ��ݐȤj	���x��^?N+~q���6����	{!�$k�Yp��#�B�r$��ߌ�m�5�}�x�����w"@7]s�2rpʗ�7?�Kհ�u�|�fy��2ɺ�80va]�o<J�J��Ѩ j\AM��<Lltw����:�5}w��q�ڥ�჻;s�\��U���FI�y����0H�Vj���������И�+�����[mŖ ���t`��A����>�n �j5�jRA� ^5"��2�����\;�W�O"9n�~���~PU�)���:�F�J�T,�,r���s�d1�@���U^6��#}*��pMC�]�/�ko�[�[#�.�H��W_�7O<��K)���>)�@I# %-�SB�Zb}���c|�:T����	�D�l%Oa6�!
����L��/�/V}[0��8+�A��q6_��1W8~�Ƃ� f=ź� :�݈GA`
9ފpÄ1D��U���v��#��=F���-�ȃ ��>�l�6����,�4���_�7�E�W�{B7ՔÁ��ʐt !�ms:3�/��Z����,�4W	>��lh���i��xlF�Xg���ŵ3Q�K�E�{u��+�A�*��/�)[몙,��ִ��V[�%�$����I�c�_�h�Μ����#�>�rT��e�6HM�����W)Mǩ��F���'';_�1���~�4���E��xY�bN���M��HsHl�4���jH)6���_fS6�|V�9�E��YZNX5��:⭈+���gF��Z%����
���ƈY iI'W�{��C��	�3#�W���vUP��>���0=F���(��Zr'�C<�~�]w���S%Nm�����~L<̱bTΉL�
*R+� �Ց��Hh�K���j�� Ϳ���ęa�0}-i>
�QZ�����{'��� ���A�� |懡�n�գ�:d<t���i�X�D�M������;��y�"�g��P����<��Դ��|mɀ]n�{�E�ju
v |}0�R�p7���*BxZ:�RT�@�w~x����˾tR��|�=0`����!�*���[k"c&4,o{}�CO�p?2z�+m*�ku�f|OE؆3���Rv�t�̕��4���Q6��k?Ȱ�P/sqvq�������zcG��<�U��lͱa ��C55ױ����@���RA�Q�V�1�q}�}-���>��W�/�a�>�kET=�{=!a�OѺ�P�,.XAt"���D�
'T?_��,�7 ��Z�Ė�^ �&��B����i��X��(R�� ��wb]`�gK����#�ht�Q�K��g�s,m�a�u�r���~���B�lז��3ɔ|���5� *����0�G��L�T^�� �鋺�80Y3��g��������s��+���qy�њ��~Ȝ�z�;��mF��V ��A��\���0��U|q!N��}P��&�l��T��=G�ə�^�:�v~��D]�A�v'ʦ���,Ra�	d�,I��$hN �v��Z���@y�*���4ڄ�,C�wK���tkG��6 ����X`�~<`�׿ޠ|�I��xu�����,�X�r��6\�{~'��Īj�����u�<�=���{�:Y_�^��/]`�qB^�P���!����@�*�O7���kl���q%�~Ʀ��C�z8�MIP�p�i7_X����B�9�w{��Au�/������(���r��N�no;�xKRЧ�u�u����bJ����?�5��H�G�1���\�:�r���}_u�����7EHE�.�����}T-4�i:��/t�+����"H�9��1�/8{�XK��צ�~2y�Ń>�;Ut�[��{E�����SR9ȣ �!^��n�]_b��T� ���[k�`�iR�0��ah�������z ��e����h��0�xp�S^�Ӎ�nD�~S|������50@��(���ʩ�a�g�ՋX��b6�iώ����hOONU���0�\�!˱E�b��?P���f�,�4n��P��Ub����V���E���sfL�w壍��'���6�6}C��yq�W��4��e�
f=X{�CmJ�l�%?D����O!8�=���*K{�fb/J7�Wz|�	g�|;J���[��s0�{�[ⱒA�����Ճ }}�Uܺ����ACf���k�e��q�D�+���?nR%n|��)���_�@+#�E�r�O������$!�?�3��Sl�.����R=�.j!��O���c��_44٪8�
�_���,���%�nHG-2e�f���.x7.Eg�[k@�����=��F�+Z��Zݝ�#��tG�JO�'�
u�6��Qϸk�i}�TpB�aG���
����5�W��/�G�*`�@����<H�~��z��w��Ω��F>�/'�����~�MU�j�/�O<�8��*ᕧq
��&�8(] 2_��ٔ�����XL�����cWg��l1��S�D�M����P=��Pq�1�&Y��n��.s��5l@��i�΃�^���ϖ�*��w!�����di������Kxp�
���~�Y#��5@�;����+��:����f�˒��MZ�r�O����'F��
�?�p
�9FB��[(K+���{�?��.~��fx%�溇�B�%���^SeVMh�<�Bb|6gGU|�Gb&���k�������i��>���)-YzI�ec��"��
�[�y'Q��~V����I�Í��ycI}�9�ƯA��������=N�]�pU�Ņ/:	L�O �S!���Y�7�V���S㣳�n�<�T�O�U��˅�m�O�j�[�Z
�<n�E��6D7�ҏ���v� k3v��l@��4��s$�-��n�yJ ��!���h_N�AK��s���){G��>�W�����61�q ;�*W$xh=�Ox���%s������5l�*��ł�pnU*Os>�^�i���#6����7���t��;?��A$TY�`'��r�>����K��7���]H (�$��u�/�Ž��P�ѵ�㥅kX�Wȵh����C��D��u�&��H�{sJ�Jd�l�j�ҹ��*����vh_���b��֖�	Ue,�1#�ُ�����Oc��B�T�����)×�濽}�P�ӝg(�'�a���A	�L�`�sa���c6;&�m����6������6s�g�������p��-�m0�%�f�d(�&�ڿ*�g��abKVk�;���)2t@7r�i �)+Ŭ�iw}~��a�sʷ)K��E&��(�E����CkI. ��ԫ�f�-	�s�����I�n��֤���I8 � �4����/)�⓴2x82���^��e<���.�L����	�s�UORsz�ą�_�
I
Aˏ�����zm1�\�h<��bR�]D������<��;��=!T�Xk�j\
w�a׎*�#l����_bg�K�mĝ�M�
�a���9|˪"�Z��.�`j�����)D�^�9�m-���M7zF�H��`��b�d���#A�`��ّ5������41�;���sA�_0���)��$,U���15x�8��m/��ZiN��Z�o����6nƔ��a�nN�@��ba~�k�F$i<�8w��ү,����sj瑭ț�tc|@�ƚ�w+�DӢ�ћۀ$�E8i�1D��Y�~m�c�v����0�hr��up�f�/�������!�s�g7Ow��)�B�����������2LJ��k���2��h��.h����?0a7IKNU�W�ͱ��]lMk��Q5��x*<�go5���d�@ss�s!
��;��O֢���Gc_����9�2h�\��,��e�����v��w��/�
~�MQ���#��q/�b����Q������S�/"���D�$�,����}iF�����i�p&_�$ˈboDq�b��%q@�a�>7T�� �lh��ze� �i1ؽ�6	��7|��E(Q1'��M�%d�Lv:3sH2 �ԫ�V�EGޓu���\����-,_���Sl��\m��/x�y�h|#���D�TJ@Mk��`2� �F��y������o�O��^v����;S�&*��LT:%C���y�o���킩K�|y����X%l"3�i*bʂ�S;@{z|��E�C�w�����%̤�5\8�1V��ҍ�/J���l�@3p@��
K�����j���J����k4�[��4bĺE쳏X�YBv���s��� XB����A�3���U��|��5Q/�B�M�+Х�`�� t���"|�;5�]C"܏�f�i~ͼ8��7V��d%��b5�G���"`�6�r���B*"X/?g@��ǃW/�7�Z��=:|��>wx����8$��ʘ��9!�ui�����\sd��H�2�&��U�} hB�e��3~�Q~��DAEG�/I!s�ӑA&`0�=Hخ3^LU���Z��\��r�dz+�;���=�av�P6BL��-�%�H�?9�a��a��n�~E��<.����ݤFa�8h5Rg�IΕ>}b��D��)F���Ç3��*�)'������;��
 ΪCX�ɯj����,kZY���εי֛3��3�i�F���	/�	�0�?
�[��6^6�J��?��O(gB���N��= #�B~�1n2���s�DeE�`��NE�]!��&���5K�(��ΟE��
�4�+�C�V��J ��;'_�(�ԙ�v@���S�d�ﲃ_h��gF�,�c�A����c�}��h mTA�$&P��Ϯ�*,a�(�Ø�� �9t�Rvf��ԇ���n`}���"��$����^1?5W�(n#�%�z��hi�H�Ҥ����j�O-��� $��[�h�j��F>�t2�ἴ ��Œ\�^�i������zi��C�h��kYX*�����$�ߛ��K��D��A��}__�2uW�:6I�����~���?E�_���L��V~��ny`*�`�����X4$�<�C��U��¾���0��D�K$+W�%��Q�C�'�Յ����>�dg�||�L���C�a=yx�^ߙ'�.rgy�p��ƅ/za��f&+B!��hb}T!�c0sF_��]��k�O ����c�ݬ0
&���/��;�5D�����s\k�P�5�;���?�<�nouk����H�Tw&E&JE}�������:��^�LGi�>)���a	��r��ګ�>�il|,� �p-����*�#ڵP	��  ]�w2Ź�Dfx�8.IA/��wwܧwn.wQ ��-���V �':�?����(j:��z�Za:��8�������zŮv�]�T�z�&���B���� +uLe�T�w8�)hJo�|L��G7^�U����+��)+�ߵ�۟�m�Q�o���ݕ]i�f��9�)<����c=4�IY��^�PT��.>�<6�^�F�1��{��Nt�X�C�6�l+���{�mV/�Ѷ�<���S�dn��BePk�2��q�LI����}G�>L�,��|�تTa��`���������b]Ŋ�'�e�v�<�
����,�0�����|���qX��_XJ�8S�B7�r�% ��=aH�4Ԃ�;	U�¢8 �d:��yT0�~^��ط9�)o{�' ]V�F�:r�����B���g@�]��
2e�A'�����GA�ţGS����*9����� op�"yҾ���m��T�5����(�Pp��F��G��qk�e���E�	2QƧA�S]���ƛ��~� ߔwL�9����z��+��Y�}��|AA�U��ISmV�wF�wQ89h��[�RV���nb�	RZưsJ�R��f��B����Q�UaψI��D�ރ�}a�=�6��#��bBfDQu��x�,��`(����:���,���F:�2���9���(�:nU�z�
=�@��-)ح�)"Ī������E(����������%o�iW\�\� �S%�W�㓫h}/�E<�c���`�G-d�>.����Na�����A�L�h�L���@��c;ş�s����8c����g��nkүj8D��H����	���M��r�Ӵa�)kO��P�o��և�	��]����P�'�}'���=i���R�/s��+y7�a���
�݁X��]gl��������Mx+דR)R���\����a"��[2ťN)3ol�z�|��ۊ��Fg{� W�^�.U�B�1�FlB�<�7j�|��mK��B=d�ՙqŤ�:R)В�ݠ2q]����1���y�v�>ԅT9�F���w�Y�qB��j���B��a��j�`�Wn V� .�@���2�_��xR?"eũi�$����PyyV�x�~A�`��^�&_�ͯqyh����_�2{2y�
:����2Y^"���q�rT
�L�BKC�&'�2�u����'��m�ۅny�A�0\/�{�����Xo&F�1M��!�tƸYRݹeI 8c%nv��! <���6v(��h|.�aڱ `2nF7" Š�m	� wX����2D�iъw��I�+��K~�vM2��vR�#ƾA<S��܍��o'�1 �#��q�MBxAI�R)�Ik�b�m�*\�1�LYi�Xw\O��$T���ī/��ː��!ȿsFa�wC^rM'	#E�&_�0���N���Z�ld��c�������0?��b��
�����>ã=K���
	H/�Bv}4qPSLeRF�G6wZFY7ִ�<�6A�m����a~j+�h��L�+���]�
E#�5ؖB�hrz;�&�u� ���2�c��d6���|^��(�� �iH�L�2�ڨ��>1<��W\U����*�F�܎�`����j-ح���}x���#�$e��g���'nC��Q��h6 h�K=e,*������	���0����~��rU:4���%�R����vb�K���FZ�3E"�^� ��hmI����8�����e-�B�����c�+>��4�Cxi,TWK���-�&��~��-�o�55k�)�y�|�%�g�-�ق��+9N���XʚԜ��"�&ҋ�
���l��k��M��Q���yJ�Z'On@���V�m=��w~-̀g�-���˰��a�� zy��>�C�Y������Ł�h%%�I�����`2�uq#���.3��{K�����S�زW�#�MF��-7�N$���p"`uXf(@w�*-� �ǣ��ţ��)�6֨�-TS��~=�]�=?Q�M�3���jJ��e����e�=puaJe.= �RT� �T��*\t��`���8���w�x�q�uc<$�H����*�����e 1�U��� Klٍ���:K�,p������ ku��SZF�Ӱ�љƔ����OWC��(5#tk�v�~XR䃫���:����[�|N!�dU��g�K��D���������P:'u���$(c��Q��A�~6�iΡ1�1籫���Z�N-�np�+I�[�ݖ]%6�r�K��;�#����j�M'���eK9�dM��3Rs�UY^J��4w
C%��z5n�)S���Jz�M���yYxI�Ҡ$]�c��Y���b�Ϩ�Ǉ??���"U�Qn��	L�W���
�-��'�����D��RK�2���5�o�}�� ��N���It��
��,l�~B����U͏��Z�e8��$��A#�le*�S���5��Y#0֤���
�沏�����a�.�����<\�[����q`�����t�P��a��e"Mf�#�b
��RČ67�ҁ�䝙k�{��7Q�G�֜Qb�#�E�愭1�f����0͢릚�������n��K�1�4�x&�����ph�h̼.��1�u�X�Y�ڲ5naz�<ū5x�u��p��#|H�$���mMP��߉���ʷm�j��l��Y����$�8��GU�I��������0���<Z��6_RX�j/���x'�m�e���0I�2�uݖD��U 8���_��{�Z�U��'Q��g H["�G^�{���!`��ҫo�Z�&�K��-�gUyo�2������`y�C����Qw��\���e�왝��'oË�c �h��U!��,2R����w�=�*}K3�~ĭ@={�Z�juz3Yzn-c9�:M�>�1v�+��q�3	�ԙo�>�����Mx�pQ��O�^���7n�O���E��5��nh���%֒_DJA�K
�n����jk���e��c�����|L�'�p�s*,5WN1�e�X��r{<b��W\ɏs�d�K����	$GW�� �#���$�Ӧ�m��8��b������3�^}x��8]W_���:��A �ϱ�M%�,����jy(>�o���g!�[:lV=Q�"��K�֬�M��+�� �E�:[�i�xIgW�~}1Q�*���f��}�Q��1Ѯ��Ը`^f�!��3
����+5� NU=꟎ٛ�������@�'� I��Z�I�xB	|+��9�~�B��Jh�Rk��H�w��M5��2BS5�ۑ��X�J!G<�T�
l�}����~���d��0X1�( ��B�N!`�7t1�F.����esegVOHoq�[����8���@x�ϗ'�%�Ԕ}���9K��+:^&$D�_�.tA�ݖ��ݢ(�V�6��Qī��/<O~)3w|�G ����{�$(�?�賴�Zmj�<�F�E��/|�72�^�1E+LB����.�K
p����t�|5]
i�7�_�Y���Y�KN�KU`�'�N���o[�YP0����[<��YԲJ�o�����ٖ���N�"�=
	�0	��nbl����E}��r֝Y߹zX��l�{����=#�i��k1���3��P�
���f[�j�a0���z:C.��m��&B�$R�H�{E%�&���:@qPr�p+�!�6I�	�f������eڙ�6�)�&�=W��"[� ��룔l�P����N����o��G����P��yT�/I��+�P?���qX���A��;�AW�RXSV�`G烏ˢl�ح��M�aĢ�����)��X_r�*_�I��ް��&�(�bKw7�r}��=A�
N�V0��Y|a]S3u�UB��I���*�#��/�8�_���	�u���o.[Tx>y��o���l�qs�����~-���ݭT$������*=�~����yr�S���&��lc��'�(x�����)?�c�חѡW��xE� i�.²�=H��=��_�xi^O��۫�0O4v��F��p'�~�ʒ�D��Ga̵Ѩ����ɡ#�5�9n��RUr/3�fi>�uY��ӥc��t�2���b�E�
{k�W�]��p��JGb���N ���Y��jhF�w��.?ݖ��{CH`�:�A/�>rA(Յ/�2�,���=Lq\���%��C��zI�F��֧����b����S�_OOiN ��]o�նr<�-���p��#�����cI�nW*6� ~B�u���R�'��`��
 w�!5�>� <:���[;�EP[�������uڪTh�vJȭ �^H���8�D��������	hBE,`\�H:�Q|NŚ+,
��O�����$�@����yP�x:5�#��Z��=��~M���K���֌@
�PK��M�|]&�t�d�Ku�+dRҝ_������6Ɠ�:uL��0Q��������i�~�-UT T��~�X���-y�ˈ3�%K!q�M��qy�
DR��+P�+�#|*�
�!X2�oA������tȝ�K_�F��I���B�b�R���s���u�5߰�������7���)�:FZ6a�5��ă�`ⳋ�H�V  >���:��Hb�iյu��)��*H�v��z�s�'��b���}�5�����v`��4ž�3[��h�N@��q�
�&��2��\d�Z��j���h1揼M��L˪�cׇ����;4FGĜ�g/�\��!��t�I�+�I��Wq
�l(~�k_��1�$ث����U5��u�mǧ��s8/���r�h˞wt��6NP!c�f�<���i����Wal�t�v$=��
.[��"B�yfBŜ��=s] ����#@c>9��V@k���	_�Ė�L�-*M�;��*h�,�rC��A���JP�.f]�ފ,EOCW3��|��xd��������p�P�ڲ���=�k�R�9�(��3�r�7T��\m�&��|�!qj#⟞ؿS�w���& U�)e����\!�(l��P�u��oc��k�@GU��]���k�AƘ��`)������h,��}�$�3�$%e��sy���S�{��A���еY]�&ϰ�A�\��󣔚�_�f��?�c�4��<A����Wf}0���Qy�}��bshm?ӽk7��萡�/��K֒c�BbCݐ�`]�V��6.]����h�G`��0b)�Z�)]|X�zV����zp���`�Vɞ�b�f;�K�� ��	�V�8����ُ�_oɬ^�0y�O}S;��`�A�����e~u���{�ћ���2��D]�P;
�H�5��Gz�!vX���I��9������TGԽ��X���h0%�d)t�?���Dg�q��f��
v0LG�'�d�������=�s��s�-��0a��i-��C��;�e��8�?k83���L3*U�'܄��$?g�de[��B������9�XQ��Jqz��Dz{O��X��=����cQY��4�7�թ��P���^�eK����I�|D�F/j��$�
��6?��Kش�!)���t֊j	i�Q�&{^r��I���b�DX)�x���Yơz��^>���s����M�����u =-"$n}�߉|9��.
�0��]0��5eTsZ\)��T�k���
�'��΢�Q
�A�wu~�"Y�y�'�G���D�����u��_g�k���OJX�2|X��tsGy���Q���;����B����|�/[/���X��sjmj2:���ķW�y&���ɽ�7b<��L#�xP��]}�*�����WuF���r?l��6����Q��C��o���� h��+���4�Zߠ���k�|5����G���&Ym*�Ϻ%(�ѐ	 �~�u!a�%?&׮�k��o�� �S6Z��	|$�M13}l��y�C��i�d����^�br���grA2AG�-�3+V�>?�5���13�V��Dk�<�b���|��w�R�&�Kx~�����?��盞nq-Tږ9@@/�Y�!O L�i�ϱ6�Kȏ����?["�R,�:'�����y�$.�9���p0�ꢨ9�Ǔ�6�NTlo�KT�q|	�g`QNʇ"��� �r:E��j!vY=u���W��z���GL����l^�<� �¦nz���(����ۿ�~WB��9�{i����:"��X�vzD_��O_�8�X�֫�_3�4(ۀ���Tc]�9N��\��QfS��1$� ����8�w���� ����5�Cpl���#a�Ή{$0�j�bz&_E��]w��� �����%��N��+��Q�������4N:;�054�}X�!3K�F}��B �O��b����<
��˒����r �r�X�&wO�i��!��dD�Xǋ��L�G��5fjO\�P�o��y2��մ����C�Z	�DY+P3��b��"�u���k���w5S��� a�)V����i�黡`��3��Q�<q��(V�y U}����V��_B��;�|��'����>����;~��s��"��e�Q���ޚ�K��oc긘���L�t0<J.D:)����ci��*�ˋ2�3�SúT�ܬ�%f�!m�"��2G�ڧ�hИC���m�w"����9�n>hAt�_���e�F�N��*_���i�{�H'1ފ7�*7�fJ�p��C��Z�$g�P�8Wn��^/���5��e��+Q-���(����4��XQ�9�"�G���j���-����c�P?�!��v�K&28H.��E�nY?X��Ȼ膔(op��F�Go��v�$�Mjgn����������d�i73�Śn���IL�Qw�i]�%�GKR�F�/�_�� C���vU��a\�g��4+͜=�N'Y"��&ڡo'��S"�bb����Ad7�|�y���T^䄰Z:_.���BrW�3���aI���b��(��� P���K�~��s����skJ}��i���uQ�N[&����|�	|�����B���F�AB`Id�ꑍ���E�2*�m�ʚ�⒯�((�̴;��A���^:(^ECoꥆ����PZJ�
��X��^�}m�z�0w@�O��-in�������.�ʓ�P��/(
E�˓O��rR33�%�--�"�)M{�;�"we�O��Y����ᑀ$���Ԡ�����-��fa�Z�Yd�nr�F������"��$�ǰ/����}G��Q�Z�V�$|�w�-F޹oL ��+Aqڞ���q���6搼�s�\��w���o�5�R�r����M2��(�ɴ� ��t�XKL�DP�K�z���lnIP�te�D�h.9cz���"F0��c�'Vf�Yj�����q��j| Qj�Jn�'쬨1ɮ��y�*4�`%Y4�X�DZ#~��7d
�X���l�7��P���<���vI���M�|iv����@�(���������q��6$ Ðb�
��cX³$��(�=�Yg�z�%�c!��z�L���DiK-=�\Q ��8gdG^���� 3�^� s����^آ���8�p���%�6�v�.��ޥ߲��U�m|�3�A�ڋ�dƕ�^>�{u���Xc���fz���}	i� �NU�<Z�@C��z��=!���p���dC娄k�8߫C��wI�����Br�oJ�g9�D%f �yb4��"�wzV&R�A��Z�8�N���`��43��W
��=�7�8Y#n��eP��jI��ڭ��.wߗQ�Z8x��R�[Z)vY�!��|S|	�ۗB���N�>��嫶N��|މ��`f�c>���9��<�0�_&�c�����+�~����B"�5�h<K,����dB=ȩ��66`�]Y&�"G�E�� �yI��e�P$N��ٰ�g�녱���M~I+7-��#�Wc��j��U�������d�U
9-qG���S�κ�?�Go��@�]�i��ƪ��1D��I{ H��ޯI��W��dJ��mUJ4�i�}������� ̆���lfg_�u��qqݻ�m^��2�r˫^��Y��8S;�개(fq��_��c3��Or��ٶqv!+��uf�r]�}o6�f�<��n.�W��n^����zW�C�j�J��z�Pm��a���ZnT1�Z]���(��U��2���1�CzI�hYh:���i���Fu/@��60'S�؆Z	٪���WM�ʵ*-�iF	�G�f�5�� FhG�,W���eT[lõH��ՖU����r`��*K}�Y_�Q2�!�J-�!$fW�k��q}�s��5�  �zYEڭb��5�(��	@3�z�}1����#��~�LE�L�]�9�_6)��/�Ӗ��Q5u^*A	�Gƕ���
b-����P�~V�.ҳ]ܪ9uUb���8���|�).���L��,�3VN�?cMB����Y���@�u���>�\�?����ȊC�##HI�s�{*�E0jy�:�F ���g�b*�V�=%5����0�l2sDn��Y�U:*�|;�9��`�+�5�� �m�~i'{��sUO~��� 3�B%?:�wޮ�	��x�ר�p$�i/�����=n��/���a�#ŧ� k&���>'��1vX���=��������㰪�1��͜���4��N~�����CxR��x	���F�T"k�4��z�|�'��j�o�x|���`�v	-��=T@�e�S� 2VI��q�_���ǉ-U{�t������{��@��J�=~�1��8��r
�0���
�y��P�'4�t>�F��O���ў�r���A��KY��`յ���XXX���S��1��h�#oU/���$Cю�9�$���%�x�q����D¨����l���P-��4�ϭ�c]�X~��Ƽu��=��5}�qa�;�2�/��=�-�K�#���qlY��E9��G����hRa5D��r�܎ת����cF	�����4�g�^��>��H~JvX*��=X<Z���Y+�G�:>l�����v%M��S�zgg�%R���y�޳q�Fo��=T�����#>Q`9-'D�>��`d$B�G}��Z�g��4��<2�����������4�ݎB�y��b=9$ZI�� ڑ���0�`�N��p�M��`J���pp�"Va�����1S����Bu�p�����!�o(�%T�>�PDό�%�N<�S�	��T���u�h���;��}A5��bc$������(�{��}�Q�G���/[:���� �8����?�`�#5 ��ꡚ��5���-��������e�ND�%m%3�[�O�G�C�-jh�l��,�{o
?%&[���~"��Q��a��@�*�A� ���$2�A�`-�#�}w�E�g�D�GRb��g��}nmӉ�,`�)�>$UN�V[�LJͱ��n�ٳ�`��v��]-�`{C�ƺ?�Q����MPF�&Q�g��^�vǹ��?�I���V��W�P�'*�v��FD��֓+;x�9�
�ȝ��v�[u�h�s6!{tAv4рճY;�j��Υ���ﯫ����wT#/�2G�A�A.���S�e��Z`���!.8㜂/���dB�����ES��8�0/�T���WD�0T%ͬ�-�7i�I#��j�ꋏ/ʉ��g`W�/�9�"W[0�'�P�^�S���{���1���+~b�_��+Z��q	���Z*�9#h���L���F�3?8;G�h������%�{�7�?��x���A�F)�_�ܧ�/�8��}��E=��,!�}�!#��GC��ۉ�$�m��g�~�6�w�"HG~/2D�k��:���G ��>�2��r��Ee%���#g;93ɯ��Nsmd�u1����Y���$����f$��"{\�6c2��!��LV������<��W��9�����/���0\R���C`���5�`�a�l��q0׆��ӗ�i�f5)><&�cHP�b��;�|'I]�	v v|L�띲���[�B��t�F�*�Z,��ٚ1$���(�Z(�iQR��䰏�s�]u���X�ӗ,���Ɗk�eJ�վ{�k�a��2P�v&�����+Ӝ��t�oix��o_���ys,��2B��U�/�Sџή�m��~�F�&+����2A�u%�<P��N�����@�,�6��$�J%zA3�N��E��"x]��AOUDF�1�cb�����;Y���7�l	��{5!� ӥJ5����Kr �����>�Ф�B��JFϽѰ�,�7�aFXN*�T*I�n�.?ږ�h���o��qN� �|u��+)��Pz#����,�k�r<�*(��4�I�D��(a|���Wχ.������@s��-���AJ ���[�/ʊ�`&��z�&*������gԽ�������@��DJO%�M���E5���џ�o�v��DR���-�ˆ8h��^���O !��� ��}/,�ɝD��D�\u�ǘL����_Zr4u��/5HxB��3@ځ�0��bv���lV�M��� �.#��8-)�����XLW�P◚榛�0<��k��9����ޤ�,�(򙀌��|�����~9�N�KO�+B���rVB�n��0�ye������q'i��oHeU�{"TKp�'IǶ�4�����Ʉ[٣�(��D��>Noz�`�P��0�f���{<������j�Z���v�24/kFr��h����T����]��T�����6�nsv�*2�����]�EԠ�|[d}��FMD��z�L�Yc �?fns�1��`�j��#������_����I�<�k1�0v���W�8�#��k`��~�+��'݄#���l�5���zVy���A|:=�&E�yJ/�����t��L�I�,W����e��~�"*�s\��<P���8]G%wz%6D|�*�� `�1�7�%:}��f�zQ�)�� �WIIH;��Ұ��iN�Q�e���K��tOb�Ig�Si�[j�뒎u
-Gu��+ԃ�:����4��/l���4���c��|�C��]/ [M���I��[hI���c[����h�t�����B-ZR��<�i�� ���O�I�6E&K*����V�*�-
����6�B�'����p�=t��%v7w�A
E[�����2j���E�M�'&oW�b�.];l��u�i�F@6�׸��p�|3Ҁ7��#���M>��z�bg��	+;�X��� #�nJ�PYJ0�g^t��6s1�o¥!"����uP_(<H��n�S����X	g��y�#��0�p���KQv�?�T{�qt�����P� �YB��eA��3��zI,����+H@�hu>Qä�(`˖�F�ڃl������6���E	��TS��@*�(R� Rj�#W>B�ir+���B)�I�5^�n�)��d�$�{f���|*��u�2�ؤ?^�z%������b����]�%a�z��`��C�B\���"e�h 읺�|*�A�!A7	�6���}�b>6C׌�4��m�*y7�nU��?��~7h�zu����I��G��
��S�����xly3�[g��`��Mt�)��d��rF��Hp���1
ek#��j
&�1�f��(e���X��Xd	|�
6G��w�Ƽ��c�+��}�����ߟ���� ;(P�Ԡ<Ll������X������q;.���*?�a��Y��cB�5�u�겍�)L��Z�t�BARB$F	��p
���*g�|V��4��/)������J�;1��l@�->]N �a�����:�qb�: E�Y ��2�J  |l]��C��a8�����"LDRRjƽ �\�R��n�Π�!��K>p���#��f��D��.�m�~�y |��LQ�{�:�3��o%H�n�����S��:*����se&�X�>�C������O
��1�,�-���
[��j0~_7����A�2��Ӵ-���p��p��~���zC�b���?d�M �F/�u��V��aC��j��X�LT凟K���#��b({�{�t��t*lG0�����d��}t�h����-FLfE��k�y5����N��2�#27#���F�Y����^�Z\PG���P<�S@���g�Ʃ�%p�=�B�@�Ý瞽��T�y/g(�`41���PR�[:b��}�vJ��G���f�h�����A�TJ<���\K�z��5{;��6QQ/�u��� �(G��pb_��d��M�p.A�#�^Z�N��f&�v�V�mu� �y8{��T:Y�B�VSyP=�x�Ԍ*�������Ehc�%13�.:No��&��_��F%�J5�,w��]%�ZNJ��⁔R�do5�%7���f�D��*}Q�o=8�ﱉ|c�S�3Oݽ���C�9U�3<q�A�E�n���ڂzj7�LK]sba5mCn�:|�����2a�:�-﹟G��*Ue����,Y�u��#�*���oa�8}���@\Vl��͊�B�#�m|��{��.�{q��4����c��KvP���6���`�RVW�\b�v�����K$������QA�>��XB��'������WM��H	u�0�0��Cc��ƛ�(v�&R=���n߳�S�3�'�o�*GQ����4��>;�W���&j�M�v�Y�X�����t��0�
��{�ӏ~�pF�(#Еm����M�� du��K��YJ#�`�H��^|=�F���[Ѷ��T�q�MK��rh�1�y�P"����eb�����C�6Fn�	j������e��o��"h��ww�-�('LB;Κ��;����:iv�z"f=ezT%E��~�hX0�k-k��ش:s�khc�&n]i��q�G�b��1	��ƥ����F�~3b}�{���	��XnH��{�҈�7`��a�'x���)��������Q�ݹ+ԍ��U���d3�Ψ���6&��5Dv��]~�e��8�G�q	�#�L�S�AV�����&����,�oF�p]�C˜�h������,F%�Ӳ�R�Ţ�?���Q��P'p�Sm?�׈4�|4�0�j�9f�^�KK����2�	��q��&�/�f�x�"�ŏ@�w�q�EL��WC�)*�=�r�A%ݷ!�Be���7 ��K�\ND4M��X[����asg˛���(��9�tֲ_"!ZtJ-�	9�5�'v���|�x��t��}7����Jצ�u5������c��Y��0��\ʹO��XYJ���<U��X�H�"r�
�������΅���3����sYDU��H�lX1�ʖ��A~�=�*΂*\9���8�ߩR����|���2�a���|��Y�m�t��L�a�)�Ѣɶ�������(M�хLx��z~м]>u�s\���m+!$��{�G�йV�����͂��T1���S��垚��L@�5�	���jXVN�Y*쉦�0�_����_��������%�a3��^P�Rd�J����m����Z'����U���DԒPfp5��!2�/J|$ o��i�h]ψh��q��^���/�5Ԏ��7`�ϫ�*&��sO�h�U�M��,�̣��*`�.�2�/1=w�]���(��&�|G�YJ]�xMA ���kzHp�R�$��� r�p�Tg��R�b�(޶i=ܹ�:���$���&�=�$������e��~~
C���=b�f� �?�c>)���i �J�?g�3���Df��=�
��<g����a������-O����@�(��N�6Uܝ��O"�Kf�����*W�MƭK�V����W,���ڼ�`��5�!���P��/�
.|������C��S�� ��:��p���E/��~�߀�ԣ`���2��9�/ܛd���R0?J�I���2��+���=s�H���썖�^u�z&�C>%łN�i9���]n�����h��6J���%4AП�Ee!���3f4{�n��;�)�D�gPx̌�ve�b�u�J�
i�U�zx-7~5UX��u�9���1�x�?�*�;�T����ȥH��X����Dt=�O�&��'��7�G�D�7�ν�[�����o��Sv;�N:g��v���=�#�ㅊa�&���7��^��>\�Ѵ�ۈŚ�OA�,pj��X��ݶm9Ա�`h=�\'`l��Б�d�q� �c#�h���M˄���=��г�u��g|��P4gcǝ�5C��EFrM�vÅ�`3��HAZ�����v]g9}��|�<� /�8�{��.��[������DVBO	��-JO��sh���K�V5~ (ӻ@�&$ L�q@�%��0����s5_$���_0�:}yF��S�r��)�Ǧ���C�&�|+r���W��;���w�N������W��`�ݽ۾ΟL�5gD=�ɵn�J�^�B�"T�$��,+���Mr�Yj� �d�C���v�������s!T�u�Ǿt��C�j`��<�k�w��Z�j}YzI����G�+�'���uw�ټS�Zt��'�p�X&-?�4�T"Aͱ�7�E!?��#Ԝܚ7H����w[97�F 0�N�^NÄM��)�,�����S�7r�K��Fؼ��R�$t򕂃�k_�Tkq_��@�`�7�d���JD�֑>�4:ݻA�d�r��ŗRj[A�5H��"bqcQ�y�g���-�R�8r4h�!�[�Ph)N��ϡB]ݙ��~
���$vn�d$��Lb�E�i
��b%�c�m���י��d|
$�Vs�|kfǛ.��t�[/�����(��ZD��25F�$⾋���:�J�,q��	f���ZM�������mfl�P�`�9&/U-0�)���g
���ŝ��ώ�>�Gܩ����f�u��@�^�o�����%ocPlV�	p!@�p�j��|"،����q�i뷉m�?Iv����Gx�����Q���^��t����̓9q��F .�[�Z�v���|�������~ ;E$�;��N�	��f�R����m��3U���T&뺋�T
�ɮ�˩8P�'�B�"C�]�r�"B�q5` >�؎I�f��剐�n��B� ~q'\�l%j������'���</Sy�ղ-��(Rz����,�Q뺇��~�䊚��E�{h�̽,1�����N�8+�}��Vt�L|u��LN�!�:{���9F?�CF�iW莃���0+���ʟ�k�!G�Y��K�K{�s�j<Դ�| ��J�o~�����.]NW%�d.�"�B�:�ҍ�P��[���0-���e��"Sf���9ࢌ���]��AR��"�j%��c��@<˧�Lݐg: #D�3�.�{���mh2�q���{5ww��dyx��xV�Blb�)�d�eH��͙��)lR'�fe{�Y��3��mM_�� S=�
�N�qb�|{���%��������#A��컀P4h'1tA��+$�n��Gj�k"�6$-h��v����H��W6�� Yd��̓2��bս���/��Ju��<��`g��<)�6>o�[��S:0�,u�8J������Cjݡ�d6d�,�k��+A1ʥת�ᑨm������p7�����ĜT��Ԯ�޾�EK� S�.��Q���@���TO�<hn�AF���P�+���)#�5���s�#/
�~$.L=�N��}k��BH�JU�=ZB�* ��
m�Ź��잔8�?p�'o�!�W�N�%H����=���(ؖ� @_ �D8��[ꆚs�ê0���y��V��M�\�̽�r�/�s��_*۫@�|肑�ie�4�������B:[EW*<oh��˭�_�[�c� 2��S�j#ug��gf���ixe)	�9zd��Զ���O�$�y7��f{<2�JϡX���_����%�i���ђ���iչ:��:/sێG��N�0ӌ�*UQg�Y���0:C�ˍ�(�Ez��u&It�;OKN�<�3�����m���(��iý|���/#x��ViE�?yҜʞ�Ö�V�M��-'=��W1����lZ_lo�VhE�o�b?�v��ϋ-L�l���, ��|��q<�4	�[���]��R/<L9J��Β��l"Ո�҃����ϬZ�x։x8K��!Y��W����ՏP�w��:�|���˭�^j�*S�Gh�h��
�G1���|_HI�4����1�?�&ӎ0=X8�`dX�#��h>���"n��_�8�B_�`A�E�z���Y���=��<x�4Wx�,��a:{Arw�ץu!2,��̀��o���҉BQ��1M�Ǳ���-}PM��s���j��~-��x��Q"
��[A�/�Z5w!��db2LsG8�#~���Ǽs_q��|p��|e�]JZ���Nc������q���b�G����ǀ�-�6��֕�y�Nx��+E(�D��*:�_+lj Up��,xw/ڳ�2)R�ɉX���Պy4��-�_�G'�ll�w�`��X 2$|.� g��X�>�ِ��x�<��?��B��,���O��3�-+���d��6'�w������	�����֔�(L]�0����{�C�ԡ�"�4������|аS��'X}:C=���@���m��7;����#���.�\O�[ L��XFêUj�0$~?�}ȘkX�EqU��bѰ�-����y�M ��t	q�z%�-}Z9���{�C`h�\�w�״�0������m�*������4���)�y��/�.�L����q�:!EgzC�R�+��	!�t�h�� �
��jt���{[W��h�/k��+T�
�_$t(�Nw��@MS��)��e��>I؈���t{9j�;&���b׊�b�n��lyt��D�B1�#�/��Փm�Z�9�Ȗ�ʌ�-�7�*��`��OcȵP5k	��&�|��'ڸՅ ���)�w ���n�WP�u�N.���q�\w�F�D�Jڎ��^��j(�i�����(��`�E����"²���	(�X�uaI�w{��b�Y�gfuR���J���Z~,j������=��y*@����ڙ���g,�l�&�䈻��:W.}���
hiE|9d6N�@��N�p
��OU˿�T��N@���*�x0DL�����H�5L������r��]$�	����RK)"���r+"�L�жK'Z��HXK��g��OI��Ula� �_�^#����h����* m��S�z4�3\�����1k��K���y�G���O��V%}P��Z��NR�5i���@`�ߥ62}���5��rpii�X�p(��$�+h���%��3���
5wq�0U�w�֑ekGs=��O`�(�В�ͽ� �Z��@�[^K{=<������4p}GWxL������IТ�1R�� �؃���p��*K�z�y��j��٥����S�ߚ�3��$^ �RV������~�˛��+#���5�e��h�j�V�����S$�&�\�:��F��{9�,�Ƞ�Ը\x\����RNb���j��	�\���S����0�W����R����w����~t�z�F<j��L#���S���s�a�pV���a(*��Gl���f ^b�C�l��j��a_V/�pER�!�_��wz]0�ׯ���te��Q@�"i��ä��WZ��T�eO�}�u��|��E@�]��͠!a9�Ar�?��nf'�6W+o����Ȼ�2�Ytj���i�Bך'�I�/��t���7`���p���Q����i]����{m׶����Z�?�����d��5
Ol\N	ч7�x,r��hD���C|�?h;��:+賜��߂�������i�ǶW�>R�%�׊�ֵ�̱:��c�1��RM�́���Fuڅ����?��.���m��R��~�w����B�2�S�Q<�9�>��
"bn�8K�z�b�x����HtH6��+�S�{�Qu���a��+eξ?�m��LJIg��7�Ω�.�C��h��M�E9��:�
FϷ��!jz���E=�,�~��9���-�J�y��p�o ���������_������H7����P���x!�.G����W���Nl�(��cG�����ɇD�Fyچ����$��^R��S��w秠3d�F���q;G������DPs{�� �Zt>e��)����[t�施��b�נ��n�;8g��8y��Ө�~���[���S)};��h���g-:	x`����P�M\5
�U�{��V�xV��"�nG��&���9@g�2��ʎ䍝!��H���_��8	��KE˩�&5��T���Q�o%ᴕ���Q���[3u1S��w�8 ��]�f���#�������h]	9b*�2�%�і�a<�kؗ�[M�Il$�H}��s�v�;�k���+�p-rS�9���Hd�8�s�,�u�̔>خ�#T�`��.ѻ9�/P��,d�з�Ơ��9�ԒJ�A�+m<z�w��0�k-�/�6�2W�������/�C<�+NP#Xrc�̀�S��L��?��<�ji�7�T��2�O�+/��η����A��q�����s�ț����H�~B��d�嶎s��c���#s��yV���ц��*V��DѱR}�RWa ge�ّ�l@[���c���QCq"���A'���W����x�8��>E�L�z�L��B��q�4� v�5��~�v���X�Ւ5u=�K?�,�;��:-@�a�QI_k�T��3�+{�����1/Z{h` �xl�	�t�����q:z�Z��4(�U�xC0j0
F}���=-�����QKm[�W���T�W��������pi��;�Ѹ�@KC��#��iѶ�_��(��d�@�o�x�n�yѵ�]\_�'�Y��bK��$y�&��{'�<}\�C��l�gQ�z_ܦ�*�t3��³ae����non��dn��%�+X�I�q=�"�U�Y:(�R�W_��:e��|'��E�9;4]�.����L�"�L8uYz����*%�.c%��l<��*�9-i6�:|ț[v�0�L�'���-�G�����5�M��j����4�V���dK��DL�Z����H�]���W���ˏK��6����I�փ;�����e���YB8C�y3��D��ӑ�o!����g�x2]�K�2P�<Z�u�μP2oV6���jN��|Y��=+�4�^ۭe|~Tg]+�ыdn0����,��2#�L/�9�mB�X^K	_�����Df�u���������(�𫽱T�/�����vg;�夲Z��B!eA�"r�-��".��3gЃk4W���;�q�X�'��n}�Ń2pR�q����p[K��7����,O	a�%��9D�YX,�����}a���Z[�v�4�,m�vw���Zh�9?gD8�l��^TG~�~����T�b�_ְOF�`k��x�k�P}}��&x.�!JY=�%aU'��t�U˸;JU[�Aӧ_���E<�VVigOR��6��Nu�����4�[��gFcy�D�����6�8/ņ03>F�S7T���KmR	^ڂ�=�%e�Y6!� �)�O�l8ƴ���3�h��a�~=.���b%f��vgǙ�XQi�g��?���1�A�<Q+��N��U�;4�F�	6N��PW�gR��֖$&�"�����E1�E��������Y����7��6ޔ�]4����6c�!�ý���_\�V!�V��� %�������������S���\��mXvB��������@���Y�s��1;������gf0s��(��>Ţ��ʻ�qM�F;�V��/�$�i	G
��;GW�*C[��`�v��$
|����~��8|�gk��帇3�D�yf@����p��vm�!�h�NCOBX4v�pSePA� !g�;�P�A#�'/��L�f1t��>�ͭ����q= �X��������y���:3�"�@DAo�Ie͊��X�9��&J`|��/��;<Ser+� F6�V~�2�����ٌ2M*��j`B}5sK�NzO-<����B�x�����z���x<�C���,�>Tߑ��&�G� p��z!_��fo9j�F��%Os��V�AP	�eއ)A��w-���t�*��}�r}���"�qj�{����1��8������^�jH���A�L�B���S���)��((����czӢl@Cj��b���2(�]"���ٗ���en�+g$��O���f���N��T����ḟ�9w�rJ��9��~�������m�DGk��B�xN(Ur�,�P<Q�^�[lfp�D9=����N�d�(�P@t�����R �k��^�2`��*�.΂$N���M�p�P^��<
��̤U���76|$B�=�
Tf=��t�5+��ơ�\w��"�27ME�-:9J{9�����~Nؼ�G�l;�C7*�rU|r�
È��Í�Y��W7���L�'�x} ���(L��f�������� �r�8fBD�㼋b[�
��m+EIM��e�PG]<���դ��Vun��3!�P����\׎y��^fy
w+� '��� ���%GE>ڝ��jW����i8bK�=����I0F#�k3����x�x*���<�:D��|����^�*%f;�\�G���1���yp�'���� �v��0��4Y>�@I�}h:o��,ᒧ�
(�ȜD1)o�w��~c�$���C��_(ʴ2���l���: �K��O�pkL�(��~:�݌/q������Ȃ��qei���--H���E(�����yCH��Ђ�.��'"b ����6)pZ�A����J��9-
��`>�����l��_MK�w��Tr
R/x�nO����KƂ�_v`�h|�-�P�Z���g�=���.�0%���d����0�ʱ�%SlR�_O�d5��YVÌ������A��vN�;?8)����b��+;K.�^���l��I��<W��I�**�jӎM�jO&W�g��t%V�t�)ф��y�>p��O�]�M�<HG���/���О!�a���㧹�˨Q�����Hv�M�&��1!SSAy��!jl����q��p��(G��AK�|�Z5�Aj'������:�{(j_�t)�"�]� ��&.f~¹�ä�nndcMrݐP�I��@�(��G�c8���0-�_ة�{5!?\a����0��������A!Y�=7��[�fh\*gen�X�k/�'�n?�C�'>f��������1Q�,�tn�.�į 0��;1̽�"aq�"F�2ދ�B�+Yj!�Q��#�D�f���A[����	0i����<��׍\o�����S�voi����N~��^�?�>�E�e��%Y+�˅�
�r�q����bR��:7�X�Z����/�:;j��V� ǅ��s��W8S`	L���rp?�*�� �j�F2h	�l��a�P�����r�֢��$� ��n92�H�]��̨J/�.{A��X�AW�n?��%���n9a{�;��,�%ȇ�UCB�%k�`P��U��yWB��Z�A��BՔR#�p������R����z�Yv8NJ��;NJ����F�F�tM�T���cĤ�^�d������hz֤�jg�#e�LQ�����E������E��Xn���c������δ[�8aY����N�m�����6K�"�л-��ȴ���_�F�~�%����J��vtm ��gQZ���?��k��]6HE���L1H��<��ë9y�n����[1��%�OPE{���k�.�����UCw�/܅x��N�k;�`�I�/���#�Rm����i��|gM*�RlBg���ţ:��1�pJ���EZR1-!|8�#���K�C��ْE{:'�[�gU����&�|��������VJ��H8rP�^������'�u��Z�7�g]�Q��Z��'z�x2J�ݯU٬���A�31m�͒-ˁ�(�D�^"��\R��U<yu�x?lgR�I45 ��o�ZN�+-�駗dؖ�?��kY8R�q����<7dc��g	[у��y�.��<%�w�����٬~	�u"�UF]6Ko¼Jb�H�E�G�v� 9IX�x���d�\(C���V������� �w�ЮA<8�JPH0�؋{�yX �a�>x������~�(�]+�%MA���JR��Y�;$�9�d�R�~g����GgM����(��#u��>���,�BcV�������^.i
��^'2� ���ϼiZZS�<�"1O�k�Ml"e�/�P.5��I�҆�a	Ml�=	�m?�:bK��$v�Jl�-�)��G02��ד�.m0�p�����r� ��_=f�Xfq�f�UU���t�d�x<��2*�^���F7���RiR�]P^�}L#`��}!|���N�+�۶_C葭��"��e};���ͅ�g_���1�sA����3�(��Oy�O�N���o ��68�X���k�T<��I��d-��
 ��L0�a�8��1?fn.�ǈ�͇�c�SD7����4�g���UyF_"�7�������&��z�*j�q��e ��gڄ���N�DB�����yIUv@J�w�3�`|4,~s;u�Ј����] 0N��2z������u%$(���L4]y��{��QE�
��W<Ё�9��chۢ2ٻ>W�6���j�m�*/�Ey�ڵ��U!穚sKq���f��*�e�	�6-�����,�U��Յ����6�1��j�+R���/AH��K!���o�n�������6*�Os�� �>��1��c�:jq���X������p%�Q~��y��L���o߁Up����Bc7�ˌ��! �G_���593}���������˝aVȂ��7U����O�kVwkW��������~	�`6�
�w����t��l�u ���ݛ�q">hA���k��du.(7e:Z(��%	N�T��S�O��u��dd\�+�i|��Ъ� F3/�U���z��W��.PMJ��de�cjX8%�
;�>3��r�T�˅�Y��\B�m�-A39jM%wm���]+H����T�
���\qc郭������|�I�P��m.I�g��F�G�@<�)��č����g"�Z/;x.���J��Uf���� �x]�i��OM �?|#Y��M�<Rc
h|�y��=�p|C��V�������@����P�XsV�'	��|����}���d4�����cʠ�c��bܙ_y�n%��/[(��E.��*�۫��> 7�t?-�5.��I8�C���c�I�����xM�2)���֣i%ב�Ų�d��e(��5+���2i�D�o�8s�!�o�k���(��n�8���R�}�Ƕ1�e�5$���8���Y��I�b����QhZ�=+d�+�^,����bctn�p��r�����`���͂''��P�{Y����q�����&6%������U0=�å�j����D�(�s-ڭ�W����l�89c�D�h�r���/�Q�<��nq�KD�ԛauM��&R�.���l�y�z,�"�UJ���K��O�W5��\�{����6�>�!4��8�N�`FՂ=�)�d��Z�MR�[Z�2t��No#�VWy$��%3v׍c�l��ه�@.���ql�����e���SD�� 0N�3��'�����9E]�Z4w䵞D�*'K�6F�!�f���^�XJV�>02(�ŀ�^r&�?�)֐�����h!b�Ϡ�+=�P���wXF�
�5V�!�u�Z�����P�H,�8S�0�E��L�Y��*�a���G|��QW�D��^�_� i%��א��-�eN��w�G	���2TB3�V�~���k��s��8���k�<��s��0������`+JQj��'ʪ�鉲�c���{�����G�<c�漅'6��4��H7��瞮ϣaZe���q��G�]�m˜4.d&�[F.o\�+X�i:��	%|!r�����j:�*a"S�H�wF;/ui;�|��u6�K�aN�/'��ى�HU>�R~�r��=�ZZ�Ӂ�g�~z�����I��<�Z��W�H:��XQ� ����P@�^}#Q���� _�9���G0��@
��0�4�������Β�%�}.o}��!���L��W�(��a�2����N�Mf!T�%D>]D`Jd�?D̩�)� ���A&Kz�"P"~���3M}!q¼
W��~�P��6j>����o�zT��"~_UCt���˦�6x:����J	�UdU��1k���z��AHz3E�9u��Yj�F���,�r[�]~���D� u��q�e�Nƞ��j�%8T� s<�.�2��'��cL;(�%���@����M�&ZQ1O�@E.��:J*�t�p��H�'F��� ���V�L���`&Fg�4`�';4�f
�/��{�ܠ4��DJRZ�.&S�Gހ��D2^xl	�v�i�8ۚ	)��8W����Z}�cLq�D��*:�Y�[���I:�qz��h������'xOkd���ߢ�T�ƚ�a�����og<��e9�P�sO������k���Z��.��Q��L�ps!������cԫ���^�-�<���b�D��8XRl#�eMkK��TJ�B�]�l[s�w�M3+��?iz�k~�,�Tj��̥��+"z3�P+����Ȏ�k�>/�������;�aȬ�RA��V��m�`W�$���)�]�*SE�̽�����ҩ$q���H+����\爹w�(*�3�$�HF�Zո&9�����%�tEޟ�p�U:fYv�Z��<��ნ3�M+�k0@#�.Y�����[g���M;�!�H�\9r6�������P�G/}���}]�&=�B=e����G� &I�F�sB4v� �ĕ7N�_f�����u+�����6>����"���]�ݸ���j}�^���������M1��`�8��X�����ϙm�
7�&¾Nh�vi�$ň1�������:	�u<��`�%ej��S_j�W��8{�g>&^�"��%���Lqr+;��#�P��E˜Z�?Oa����̥Q'��7��R�÷�*��4:�$�AH�I�{�0�����R�?ڎ��8��Z�lx��n��|�A]��P���`*��Ni}:Tkka�ï�F�B�j�i|w�u��%3�{���mt��17�v�Y�_, Lp��I�H���d|:��[�X�/�+y|N�sz�d�r�r��'=�᭛lfl�_��c�&6��4���eC���	¢N�PP'��į�_��&��O���	�-�$re��P�L��"_��Ey�|ʞ22��';���߸�u[���{�$]B�_H�+&������{Ԧ$�X���+�%�s�rUM~�6@��*�[���_�kh0�1}���������|)Ou��:sS����%�͠L1�@��c��r@&t�4\$�K�
]�e"���'��I�	�_�y��͌oY�`�1A�)�5��7]��E���O?m� ;��v��_:@4�����<���e4�s]	Ə���N'��rs�po]Hb4����,�^7Y��[����_D�ukZU�� ���k����TЋR��ԭ�����v�خ�)�*?�G�a�LԌ�湀Fz~�vE�{α�#B�Q)� ����$Ӗ��M��`�tH�S��F���S�W��2�<��9V/�)��癩CC^���X�=b�6�%L��;k	�a�6�D��d	T�c���~8��|?l�V.���?�9���~: ��R?~S%:�Y�Ī����h���
��/����%�L���U1h#�+��-�锜)U�;{H&��iG�K���̝a>n����O��ۘ���Lg�NO�A_�C��S�{�^#�V0��)�b�aȲXD�6p�����F�s��m�jΖ#��/��9�q��b_�\.@
wQ���S�kOV�o�$TN/�q�֠dD��?�+S�R�2%;`�m�53H����d	c��g��1�AG�̞f`����B���BW6:���9+��L'YĜ%��[o���.�U|=C=�7�_�ʡ�JX��UL�ht`T����4t�p��9�QL�
Y�u�TjtPm�'v8�%"�O�:vs�4����
���%U]"ۄ3�6��mF|��Wiq�/��i����G]�Z�3�ҩx|�:�8�u��w����L�$J�)�e'�pq�����(2WY��D���r����[pU-��K� >Ģ���s��]�]XJ죺���ܩh6�+�����k'+<Nעe�UZJD3�k��cY�Y����[��b�g���_�B�G��.�r���MEB޳��y�k�-�Up��n��E�X��5v���u��y'Uh�:]�\� ˞�A���.��%�l�`���#�͐ ���1	J�n�}�~H��	Y�G^�~xu�Q�uj]N��-"or�5�8�`�5�{������h箧V��>�u�{ǵΒ�I�z�z��L"�Hgc�G�Ք�}!�x�Z���
"-�W~�V�x,�j6Ňڑ{�5#&�������1I*�T�����@�a�?ư�0�ͳ֚�������l9��
�9�#���S:����w���9�Y�G�Hik��o���,��
(YC�I����R�3�*}"�F�q����B�f�&=I��*KG��Z� 5h5���-ڧ�n+�N]'�ŗW;�U��\��t�v�1;y=i_M�>6i�b��ps�Lpٶ�Ͱ=P��:�H���m�gNCԽܯWP���^�85�wا����d�^�,i++�RW�]Vf-�@p���z�"Y����6�����,4ΑY[x3O{�j!	��L���Xπ�s�D�a�>7�`�B���Udww Av�������kRY8Jb��t|��K˖�/�VG8IYJ}�0�?�h[��Fľ�X����@�j�
Ko�5 )o�-�M�o~�1�T�u�f��� �����_.��WK���v�ņ7�*�&�j}�8�����cm�?�x����/���B`g�� ��"B*M�3�>