��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:��������uA��@��y���<����xDET>��W�����C%�=U����3v���hj��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O��^x%���c_��$i��b�q-����O�-~\�MRTHx��Z�\0M?)���w�`+���AXS'��28c�
A���j!�ng1�-⦜������Y*�5��F���c�ۚ㏏��� <6`� �\�N~ɄC��+���>S}}�1���>Ac�@]en��}a�˨�ګu\��ʌ(jx��sR������/8Ew�t��s���<.oi����Ѿ��jZ��E�<��B�^ ���%8HY蝈�%���gK<�����_�	_)q!��w.ml*�DT&^~~EvT`�3|Im�+�z����'������G:���S��ye�K�X�M��hr֤�Ƚ�F�^ xC=^g�|�6@
8FH�~���o���p�\�u�o�euuM���Y��3w�=x,Y���q�Ia�7=��UBQ}�dܭ��r��Y���"�W�m9�z�<�ۯQF�9�4�*Klܫ���A�:��ѹ,���vD�G����U�楇���<4ݎVP��rs٢z{�����|D�ا�|Ƀ<�Z &R�Wqh������6�3Jh�5��F�{ �^�n[��bA+�V(-9��'ڞ� Jj[����Γ��o�S?���(v�LZg�)t�� ,8r:L���6�W�ܣDm��	�v3r����w7ɍZ歊�'@=�K�LZ��0��4b$�������.�7���Ā�2��CV���snJ�-75���Y�^c{$��'��?j��:�N	˵y+�a��At���$�rgc*I3����>�AxTᵏ������\�Q�G��T� ��H&�� N���*�,2��8YW~4��hH�Ja���N��ZԦ;	��Y��S�{�4�A��O�� ²�x}�bX5Z?��e�������2��
��)�
A#S-����A)�u��ά#�?.S�,�%�(r�&s��q����	V�P��YWp�a��:ꎱ)����(�?�-z�AMz5� ʘA3X m����������*�z�sN�Zi�%��i橆"���n���O8�G/60$���t���tS�9s�	���nM���M%G��R�_g8���-B���'0�_%Ģgh�UDa-a2fƀ��U��F`k�򦨉���w�u��Y��5����o���q�"�e�I�f�	��L��O",
_�7�) �iu~�a���e�N�B����}}�qZY�}�1Ub���5��y�^��J 3���Мؠ��� m~%6��B���!B���̱U�}l>�FI�X��J�:/C��E��
�3�L��-�7i��8��P�j�:]4���wK��e,︱���]*|0ah�_��!u&nz�s<%ӏ�R��[�[�AW¯leY���'�,�l�hz��Y4f�`6��cx!�pY]%��^���k7P�1�bP��6\m�͆X� �-��J�h�Z�b�,�M�8�Õ�L;��j�\Ͱ5e��<%˂ �8m��㞵P�
���z:�'`g^Rv�QDE�fD��=g��{��q��ҟJ4X���T#��n�t���7"�nTr.��"Dho�'~'����T�H��ECbUy�ބ�"��/ӌq ��e�k����B�u�\�X?Ѫ�����K�k��Nb�#�T���B�oO~�\(�VH�v��&y��/�����q	��s���a)&0���[{��=�F�"�JlT<˥����7��)��@���4w=��qb`t����<���u/��Gf{�H��HR�[��B8:s�"#��/�{5�e{`	�(_k�����īU6������2��+Z��e�f�e^�k�F����Wl)Y�gfy�'�
i.w��b���bV�S��36닙}JF�!�i��$��]���f
�-�+��<���Dせ%9<˞^�*,I0�f�9@"��A&���Ww'}w��w2e��ĳ{�/����ф�O����ko�7�����A{8�`f�9H� �ի�j`���4��V<�q���}��zcǏtw�#��I��6]�=]���L�M�S�M���?���.��ft5tv��%<?���n����ʱ)R0
+�ˠ����]&�73��e�M�5�G3�WzT��7�kH��XE"�K{���4Y�ٚ(g�?n�cN'Ի1��=r������ے��oQ�|��P����YO�HΎgқ/� �){��g��u)�
��:p����L�k��Fr=ƻO�>�]��e
u�We�/4O�V�K����}�O��|W�M�T�s]���d��U3����9�ɍ��,[�M�*��)T�%�rg3ޒ*�^���_�t��أAotv���*۲⏹o��3=gԅ�p?���Ш��w1����3�ŶG�����Y��Ȑ�q�ɹp�c
�~(|��=(��X뵢��Y&�n&��Y\z9"\W��^����.�K�u�	�"�y{{�Ó$�����M�TJM�=�p5YΉ��G�fm���?��P��S���Ԥ�%�,�q�+6�N�x�4���!���P�|��)�v��9\'Lp�C�1G�9�dnF43fdr�x��>2�&s6��o�z��/�V�hu	��,��m��2!�¬�ɶF�8�3�$LM�c& ֲ�:K���N����p� ��,"�Q0EŕՆ*Ա��Oa��	�5X�.�#���A�6;Q�U�$�n��n,t0��S[0�H	���.eRFg�y���ͪ`�E�	JgE�8&<��(V�f�h+Ў|�yVr x�A`F�ե-���H~�h
bڔ!Ӧ�cy뇇�h�h��Ipr�4����{x�.��O�#�F>uݵ���
�.^b��Ȃ!X��81j�uq�g��ql[N*�3.7T�(���;�ز�5��F�Hd5��x�Mē*��X"e5-X���%�F'+.�{P��D��]؛������[����~����؇�"�1�C��f7����\!����0���ӽf9pIL�� r��i�cm�����榥�^F%FH�����d�6QM�1�~��/�L ��Hn��s�Xe,^����Bg�ď�^r��wGߏ����?/���}����K������GFE{�&�ЎX�K��_#NZ���M|�lrx�GU��gy'C�pNZ��E��������	u���o|��Is�p|@��lꩽ/�P�T^��fø�UOWBt;O�&<����	���.':�'��f$�f�F�_�t�d(b��yXh��t�������1��mr�:%���s��eo����Q����Y9����l�,@֫|�4�8��J-%�r���ƹ���ǐSʛ3|5V�5���'o���]����,��(r2�F�Y��*ʊ�&������I�������1n��lB�0]�Iw��渎��ro��3�x����}��z�5����%C.��nb5_>6�@R���g��є:GZ<�P���U.�r��3�J�`�?�W$n�c�`lSt:]k�O�Ky�|��#�"��ʝ�~�Kv�	+ڶ��;?�ɂ�GެH��Th[��K�aٍ�����H�>����3" �����I5(���	�l.��h���;�t��-=T�[�!�X!)<�F\�L�������K.n��k)�
��xL:eT� {�z+z)�ďY}�q�S��+����`}���0�x�n�4�kV���$yl&���zOF��?��ǥ�<̘��m�	��2����0���*�!����G�z�vؖ�z�����RIC�k�8��5����� �z'곆�͹X�)�@�i�,�^.V�,1�tn�<��
(J`)��C�k�b�׳����)��;l�eq>�8��	$���Y�����=�Iĸ��3$�{�B¥��V��"�ۈ�'4��ڿ���W!̼*+�^�����5��͝�'V�8g�@���v�D@B�dFB��8�̌�ׯ��;����ʎ�kP�LNw�F6�&	�q�QE���B�7ٱE�`d;QH|���8��*���w���OrSb��Q��a��E1|����|�<Vz��������{��<�+�HƠ���;P�|1ܿ�:=����
��գynZ��~����Bb=i��?�sc���	iS��8Y�-�"[|��ք�KZKW:~�� �L*�e��}�uJ�ʐ�&�|VE��\�RV��� ��ae�7^�IN�5�B[W~�b�8&'��h��jP��4\�Qg8==�>S���of�E�p���6�ş���}s�wR&�9(�����'c����̭��������'`7�~n�-9`Y�ZA�$X��j�����S�U�sg�<�Nv'P�J�-�����Zk)������#x��S`|���h"C���}��&)�#����QAoWz����ae�(ʂ�ɐ�ɀP[Dp�f�~_���3:U�y+W~(<r$W� S�4�@I)�K��^M� Шz�W��P���^��4,����PcT�f[�>#�&��z�V�a4�yq2�+H`<�B�(�@�����),u
�@���B� ��A���Z���|	S�w�md�{��ӏ�Y8�����0���1/����y(��[u3�����@�6�υ)�X㴸)����d�s�'��I*���OS�Z���#X�qv���F�[���P�Cƫǩ�ծS-�KѲ�x������78ue�>L1�ё�F��@^�����/{�pBP��O�~eL�ܔ,c=:��Ӑ7���oqx�0�{�Cе�{�k{���95�g�e�K$ю��Ւ���f(N�E߷͒y"�1�"-_^�� � �d�1�qΪ����ܕ�5�_�&䋧zJ��N�5�ls,9�:X6��W�{k�]��J1>�����2�zE�Q���,OX5�,"�F.��|��1�~Pe^�:�9~�7Đ�,�#�)��V\U\菻8 M���8�\l�C]=^LRz@��M���L�ņ�>���ou��`U5@[�+B��KoK8d���c�#�	-��Q�o��Dg�ޡ6��jF&Zd��A��f�����V��II�����T7���ԡ�A��RM�b՜!y�ֶgg
H��)�3�#ً��)�g>����&g�Sʆ|�9ݠ_�ߚ.(.n�-*�a��1�ڰ0%��H�P� ­�#]��gА�O���q��t
G�%�!,Ǒ��t��u�9+奡��D��N��R�b��j6�������q���Ԝ����i\V�Y��J�xA7_�9嵌;�Oe�t�Lv_�>j��>Zw�+-n���U'd�'�����4/���	ƻs�ۺgj�Q�c��8�t�V&uTT�z	�mľ���G�~��1�:i�0�g��`7B�ZS�k��g��p��-4u�T���9\b��e�����;�I؀�\�C�ۅ74�L6�U�,lW�'�D+��{؝�gy����ų]z�+S]�O?u=3]��R�I@�M�hB��*���,��mnv$��]FD�-��
���{$ˣ	k��Ơ~��B9<����́�Zp@�%�JM�@m*ЧV�T�����G�\�{P��݋�s�U�Hŧho�\B�׸��M�Y~��=�%Mcb1�x%-�H�e)U���q�&���'�]�ir���!T�QDXcXA2��vF@\^-�k�t�z���c��n"8��0�y\�,�mu>qP�Dy��_�q\��m�.r~�4XL��W����բ�	!��L�{�����2�qJTX?�~��AzjV���jZ�X*ݠ[@,��.���N3�Q�֫��E]V��e5�R��c'�*�	�b�`�"bի�:4f�?����z� �}��FO�2��� �T3܈ċ'�S�8�U:��ؠ#����c�Rw��Os��߿�c���6�'2��h�����|�R@���&�����h�\���x��QZ����E���>���!	��m���郯52�#� hÙ]���%��9�ɒ>�ȶ�^Ŧ�8f�Pj�6����>5SK�7[F#���gV{�E�Ϙݥo�
���%{����: ��N�2�U����XN� ���/P*�!l�u2c;1$�P��QI��(�h�<�A�b��cBW�K1�&��w&�RВ�02ψ#�f��Q@A��$� 3lHf�]TEXu�gX���/�6������u�%u&Ĥ��-i������&���m�#g����ba+��2"�~}1=q��6������B(��,�u�]�Aw�����V��M��>؟>84Z���Q��TmC�O�Α���_��o�q��x�.���/{C��z�-鴏.�	�.|p$��e�T(s mk9I۳ �XkN<4�� �܋��𢜢k*ZT�����U���t�Y�d�h6�sɸ]:�?O��b�SU$qa6K��9^�9TO\e#�p����3��E=�.�+rݭ�U�^���?	q���3'��������f�,:��tP2����*�G�X�o+��x��j�ѿۍ���a3�P3�f
\�[p������ByO�y�)'�
����1���KΟ;����5�ʛ��TNd�\��(�ִ��҅j�5�ߕ���4;7���rS��
i۽�)da�y�����Z$9ɇ��>vT7��i�r5Ç��~e\��mdrHr��(�ʜC4%��t�Z2q僞F�H��7��$��݋��}���
ݿ�?�P��m���C{�-�g�f}��n�&�s�	�����K����"�c+���YX]�V�0��X{G��f뷠��j��Oe'D���T@J}}O
�ǌ��P�_�fA'T���tF�O��tw�I��5�|,4V�m2�^x�}�!�O�K;b�4�Qs����m�v��^�B�T88�"�Ps-������"�"�\�
G���..���/�%w��ّL��Ke�-4��i�[k�i#�.�>�%��n0���5q{�V�"�C��&��^|$������޺Y�~��!ūm7�0t��o�Ma8��g�(t=Z�g�n3��&������W�fx[@���c�zb�lm�h�^H�N�8�bZ��|A��c�#�y<?�?�����͏ϡ,:Lۊ��������2Em��H���r�Z����#ߪ�\b��y����(vtnZ���1����Io1����Ă�Fk�S�F�]��.N� ɷgs��2�W���f�?B�+-���������Gm�ra�<���d���5�*�b��B�Єʒ��1��