��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v����aW����8�]�T�]�6:v�&�CMl�g�x�J����l���WP�C8Q�����
��1wcf�H�Ĺ��.���I���v������> B�G��3�2Çb�ZS<a�M�b���>�tE�f��ԏh�����b7 Ql��~��x��P�"�?�t/�x�0����N4� r�b�
���U�v���+{*���� �����A����_��E�r�.B�q�t��j����`����];����fD�Ie������� �C��)h�ChD�N-���8wV�b$�1)�l̹�c�UR3a?4m��>���-=ϡF"���B�����Y�?�ѵ���-�<�֠�}ʦrP�k�?,	���ܕ�����	����.=vu7����8�/�'c��.��|=��n2��L(4n��\u���Su�s=��l)��-�7)V�A�80��o�*��cr�b�307_A.6<`^�Y�@Z�*�+m[�)��&ɘCpQQ��g))(���"��������}w��3'v=(Cby-%blx��p�T�w}�K/� S�Jp�E�)t�$��K��O4�}ڭQ>F����k��+�R��C��� ��X��J�6*`���L2�$�H
~�O:8�r���:B�;��c�׷p	��^>68Ⱦ�x؂^��ɻ��y������ǭӶ]��}N�_NRiAkt
}�̳Ls�1]�,GP�
s�P|�SaHy�dJ���Q��O6�]# KY huD»K�]ݎ��B'2�[T`���(����5%7�]��Ε�L����/�l_	��H���;�~^�xΜ���h����Z����$}�8#�.*�V��.�F�՛�:O��I�/0ڇIP�Ej��(̀���g�?!Շ2�k�O��������rKѹ�%�iu�$CTN�E��V���[�â5�R�ų�rerHx%D��'��[�]Q#gT��e(��.�U�@2�Xeј/%���{�ܹ�U��(�����&���@��,��!���ڲ$��w���lD��_P!ܹ�[�@S�0�f�tp;￩m즦l��/$�$ݜ��Yq:S�����Q�����NWK���k�L]�Qf,���┻@�lxe,�9 �g��:���x�>B��{`�H�t&h���77�M���30W�N3��,�L�??�����h�E�z��ۢzǵYd�.��Wtn�c��j��zg$�J�|��2JN7��P�-��I06ԁ���S�_"����]���q�)Ϫ�,��T�V�<̻�4t�MM�	$�VI��R-k�p��O?PZT��"Ũ�!�ڈ8��Fc���f�â�i����T�AJ�#�["j���X ��:l��T.fڰ������%6=F$
�[}_މ`F�}����!%!�U������]:��q����D���y��L$�43I����ɞޮ�g�q)C�\yT[qYc8���8�ً�ޔR��B޾��������/ۓ!r��6˖I��݋�^$%�����Ut&/Kc�|g;t�`Q��p�*?���l�8$?{�v��n�C��	��Z���߾� v�-,U��{����C<���0H�&^�H�N���_<�ʃ  ����Ũ�~�l{����+ۄ� o�L��l&��q|��8K�H�a�rEV�2;����A�Im��@�|��y��?+�w�r����L�pǥ��Պ�R�&���{NZ�Z��H&�?1�������}"�;H��2^�f84���t�fC��#e��5+�y��5�e�m��#G��kb3/�n��Q����7�_��ԁ-&7�{�&���j�F:�5��4ig�1��>ч��Ⱦe�֟/�
xH6���U�� ިAT¥�C4�PW���{	�έr)������u�h��洛zLl�e-�?�m�y\�u����q؉�Y^�o?�`��ʇ�^��5wtKʿR̛�̳,�t1�Y���fݛ���HS��b�v�|���3��R�� A8����ֽ"�1�!ϭH׵Bާ��Ude�����;�B�H0�����ǇfP���;(�֦���D�]��4�x#�S���x(�]/�%3�6�3꒪GV\y:������N��%<�o��A{3r��x5���d��=�CG}���M�Ӧ|��6�����a$.�p1U�g˫n����sC�=�w��8�&^;-�W�B�v�@��%�N;I�5�-(i���˱V8WXrKl̮ �W��7ܬ��q�Џ�>Ї�zY	ܾ��㿟��GH�{rB���a����I[�	�]����:'CT�V�|$�Ԧ�Z��B��I=�@�tW	�U��I*�`�K�L:B�<�eIEޤ�.\7_��v<�
���%��}�QɪJQ6&��A��l_P�vnx|Jy����)̮]I��)������G����T5�U�P8bф�GM�gNE��<?�٠�U�ٶe���~��\0�넓��fA�  �㭇�_rH8�pbD�����W�l�˹��zE��M���6���G���N�8�b����nHe�v �	�Ƶ��K�7&�>O�\��Z��+�w3��74�T�>��F�ʨ���AX6��\�n�����gĜ����)K\Ӈ�b(�#v�⾹���
�VZ�򛚘v����HB�B���"Sh�KC� �x�S���I��;��D�� ����%]�<.X��JFD1$ܐ�kR����rR�hʢ�����3t�:j8q�ͪ��<R ��.�I�CW�9M�y�r���<��p"��W��a�EB[G�Z^n�%0���<*Ot�1o�+N�T���|-����D�h�`��C�,��N�P�*=�H����K�P������H&��,[0���^��s\6�M�m���23Z�:����b�k��'?�W�'[�O�[��O�|��N�.꾢o��&!���#1�Z̻���U`����x���[K6�t�l6���j��^%�ˮ����r��:zF�EYAȼS�&���gc	G{׋���ѧ/�#�2m*fŞ��6�Aq�G�ƊAF@�ڴ�a^��P����}��I�>_Ъ�G��(R���cY�#��ABKr=T0�`��&�	�)J��pF�3���a���=Y
��9�>�[��ȇE��#-I��5R��e<���w�#D˫�(w[��{� ��5�x��=?΅��h�����Yz3h R5�FSּdܶ =28h%0�A6�W����'�p?��L���J{m`���cȗ@S3DlΕ�v�$se�Sz��/�@ ������O}u� ЂY"��.u�L�? ��N#��۲ߚ[u�z� �������W�eYJ+9�^��,�X;Sw�٢��xQ��i��@���`|��D�e*�Y����A�����١$���C͊wk;F*�+M� ��s�D������|.60��D+}׽M�SO;��$��p��L�f��YM rA%Uu�8W@Y�֮�f���D��^�-���ԟ������h�o/i�cV}}�Ѭ,��/j�IWr��fٺ�1�6j��4xk�-z�_�6�����u"�t�<]��jup�+