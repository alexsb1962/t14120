��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����߰f���%�w�$[��g��
n��s���!~�b��pв�_�nm�<-M{�"EE��+�N 7[=�5/�N�n <3����Iӝ�껋+���f�c4�
T�n�d�)� ��
��S�5�d5���J�2%����}ϺI�C<B�'��~gx��K�Pr(�`��2�'Խ�T�"���r�C��@�;��yoG�9_������ ��Tt��Sʓ��V\�����`'!-�yh@�zKD]ٱY\���&V�|��'{���� �g��)��{ 28��n_%�*��[4G_12g^�Y#�:�v�
�o�䖏݉a%/��#�n�
)��~U6�~Z��i���  ��Ĕ_Ў���n>��lp6��jQ�9W������j�Ɯw���v5�T�Y��9諸K�;[�ϟ�f���l� �c�_�w걕H9O��M�Ӓ�:�����4�����赵p>nW{fvHt2s��h�kRFj< !�5/��b�v���^A+�ѳ+��UM��y�-���[K�໊��8*��P4C����?hף�� n�>݄?��H�K�bl�Q�9X�}�~^�=VMY8���8)2���S�0&��k���.��xTrd�!�w8_�O&���S�	J\��v'z�?��'�/��3C�aV����MQ/�?R��l�dP��!5��8�5ǭ�|����9����[*��2�>��?M��>:��}m�[(��v���r����b-���r�e�䆘�\b3�~��:+/���I($�<�0��?ܷ�! n�4�hV��.1�mpJ�r�����z��k��L)�/�(����x2�p
{�\>\��)9�F	��*A �Fzs����FM��
@��6i�- }��	�����ƹ���C����8t��`��@d6�g� x�8��cWy�с��m�Hbî]�<n'�"����	��y�:Y�X��H�����o�P�6Ժ��w����j�`"
U��9�LU�@}��������Ny�s����h\C�Cr�M֩��ؙ�^��{�똘0������}�>��>P��u�]��=R5[����F�y��_YB�CZgI#�z���6�Xm2����=g��	�K@�es����~�-��Q�A�]�A�9��7D�k�ޑ~Y�)��E�]��Y���Ue?P��l?�'ah��!�׍�J��)6��1ϖo����U7���8�)�N�<Ʒ��$:�gز7�i��nf-�!n�.@VC��1k׸�������s�����Y��z�����ܨ�e�/�9���5���ے�ʓ]�����ȍqz��c�n�F�'��J����)���W2��K�z�m ��x�ˑRR�e��{3��آ����(��.ي��V�AH{��(Y���z�5�0&3��L!uH�JD��UO�".7��04��1�rK+�+H�o�BqgIΓv0�ˠ��o����O�҇���=��KW�͘^X�"LB�9a�cn �Bg�I-�ɠS���o�<�&����!�b�A�#�nI�(�}h�LBE��`|a2s��	4�٭�gk�P��y_w42h"�l���,�?�9�'�9����J����l�ɚH���x���Ά����pK\=O^���3
rȠ�?���9�c�H�-5�t���Z���@���I@ �>�q�v6?�����Ё봓���p%�/|@�l+,nZ��O��Z+�?��>' 6Tjst[�Ygш�U��:��ڑ���:jR��î��t��%�Q%��ص�y���K ���j���E�H���e@�a�CU=d��3U<8Y�m��9�fr�*��Ujq"t���f�9i')�U�XA�K����:�jݴf����Pd�y����o��o̥6�Yז�V�v��d��o���PZ�ၪ�}�f؞}�E'YfĀP��V`'�����jnK9��dq�xg�(+�֡-�6_�y?������qP�ڲ?h�Ī�V����e����p���Dߋ��a�[cD&1�����qq#�5����P D�WB.�2� ��~x#�d#�y,�8g?��b���] r;9���YP��Wrz"T�Y���"m|���`H���N�˫������\��=!��P���`�"��Î����"h��~����I��t��, h�g�~?�_Ǆ��y'�wJ�q���_��L<!��g��	�SG��O��>�Xa�y£-DSv����ڔ�6�{��^x����4���s�7h��I�^���Q^���u�B{M^�dY���J���ri�ʇ�ȩ��t�E/4M+�Mt3�/CA���-RM���-ډC?PX�d�]
 �Yh���l6�����.pD>q��@YKd���<*������W!#%�$���h�8cME�8�#ت-���/V�ћ/@�D.����awb�`	�gW��+�&��l�o�^}1l���[xr%���Y�K�����<�ܗ���΂������n5VZ�Qo�`�7�X�#�a����6t<g#B1c�~��>�~i�PK����Ah7�W��B*;ǰ�k��)"+C������n-�bU�r�E���_���#馎R�C�/������>fJ��PRn�����Ff�ElE��|cY��q����Y�L�-����~���\4�թPdm)�p�_��o~ĂF�d���.��pӴi�X��O�~q�K���B0�2O�������B)��δ����|"����Da)����.�ڬ�@�9_�e�]��N\��ӛ"͙�����ݠ��	(�F��,|�]~Z�"�#�Qٟ-`��g�5V:Lk'չꕔ��8�b&'����{���$�]�hǍE��P.�fX���9��e|ޏ✢zp�M�3�'$$�t��5���:J�El!{��u}S��xoս�Z����G�FE��ʮ�B�F�����G���y<���ޜ�X0��hB�\�m�a�W�_=N���mlᄲ���'U-�"��uP�s�x��i%�y
[�4���ajQ�BM�aՒ�ئ���2�ZlS���C���)�&�X�%��Z�C��1��d�vF�G��(�o�=DG�D��lH�*Sp�7�_f3b�d�������~E�e��y�7������n��B��ݿ9�v�`_Y�ŋ2;��v��Q���q�et?�wF��܉�e#���-o}z|ŗvP�F|w�;ۤ�����S���*(��M�`4������9��&�Dn�)u��+��lL{)���\�r�$1>_(ݢ��2"�a��i�\�3�ڜ� �u�G���@?Y��Ӳ�(�}y�{����C�Γ��0v��"P�!�\2��*x��`�,�r��1��tˣ#q0�8o�0�EeBIdY���S��=�N!�ϴ93������u'�:�fc3bUN�	z�x�&"7�����[��d��e���,'G9Yn�4ږ ��6_�j�fݟ�d]8D?_<�?�ڿKadK��DG�+�T��|#�R��#�ai;���n�;�w��&<��
�n�}�����A��DR�xWLs�@q1�#R#�!_Z;ܬ�UU�)�D�!'�C�|=��d2�����;O�����MZ*VO��m�5|���_د��US{�f�K;!��Ј����y����4�ߓ%[�͢�&~y��9|��j�L�{��ZdW�R�����;��&�x(V�]�h֌a/�����8{ׇ|�>����bx^ݫa�!���|��6+@�C�vF7o�x�[�2(J<�{G�[��<����P��a~�v�DCif�O�
a�/�U��n����6�k�`���f�����v���7�C�t�
t"z��m��'B rJ�?~5	�����E�a��C)G������V�P�@Qڻ9���6����&��ӳ5f�j1��\����]�V�)��������T��iOY�K��ƹ�0�ki+X�W�ˑ�vq,����6g��$�qA|�\���s_lFB��k��y�5�a(���e-O!Ⱥ�'�ɬgS�����*��,L�c��f�ǻ\}� �!<�Ŧ]��c�>ZW��弥1�9���b����n���t��0�oI Ù?�Vů��A)���cκ���,�����@4b=��d��P�I�w҅�{YQF�I���d�Ἶ3����m.��f-R~��h� ���*�� ��j
|�i��v}a?ů�C���%/ӥS����6��Cmk���@¸ǘlAQ/�=�S���ޅG���N�9ٍ��<t;!��U�j�"��)	t�M�8d�נ=������R:y�2��*]($��q��i2E*�(l���&O#$طY["��Wژnv��^�{,Gs7y>0izy�/B�2���h6��	\��R-�B��������u�� � ��S,� �|z��>�o~|���c<઴�i�5���.ÊuL@C�p�J��1=N=��A���3}Ԅ���>��J�����[yU����do�
��7��ja�:a?pEch	�RS|`E#FG�7t����r��WfS:�F��v��ߺ8ģ�v��ǻ��A���D�9v�>�^<7i�d敧 m|7�*���n~i�qER."�I����9.���fd�Bmk����#å؛@4�?1ւ���OH#jpb�{I��0v���}!?�
B��-4DR�J�guc�¤�̐R��A"��NUܬM*6�QpA (t�Luq��E�(��S�3C{!MB�S��K�iĖ�!�R4^�C�ﱲeb=�[��$>ב�b��>~�&>;
0_��2�i�ਸAn_4���6�(x`�r����_ ƽz���im�.�s1씕w��Ӕ�S4Y�w�XF:�S�5�
8G�tURz�{��@��!4o/<-�kg5]����ҳ�ql@�|�km�
�>����`i��g#saV=���T�~r�{�C������6����,���[���-K��dK�Ĩ�/fl�Z��DQ�;�٣�=>_o���^���a5���^��e�
¥��Ɍ��������N-�H��k�w#�\֭,�Av��R�ɓ佪�z����W�eS
�?D����`~wQ�$�/��fS��Q֣ ��@=LX�dhLհ?�k����[���툐��|0��i�z��X�	kU�^��!��F�B>�]�����pح2��6��=��F��:e�h1�%�Kw�`UHDÔ�Y}GO���	�g݇��y��Oa�ޙM��Z�-%!�V�3#]E*;��y��>T��T����zo<��3ݨ9�Ny��G�O(rx}Pv=	���u���C�5�Y D.o~{�H�.�x��]��?!c��{˿��$iXb�	ΣəE�N�x�k���cE߳%*��c9���s`�8`��#��)���=����.g�`s��U�L�	�d7�l�0�egm���=W���t�(����1oh'����v��SL>�����VH	yQrT$�#�V^��ň�t�F��$��P��W����\8�Hf���~���r����y��ԓ]��9&�ZB��m�O�Y�f-M%N������'PD�G��������ocj\��lǥ�&�d����@��K�3C|'��!d*��D���)f��Hy�1J�Pm$����H�v����c�0M��#�_uvo�Z�ֳX��?��mx}��pLߒ��}7TQ��ЩX&� �R����_�3�a����%ؑj��:��^/�!n�;$�ʵ
O����KB~��tBB%R"۳��i��ɸ��4����ƣ�L_�
�8
"�� ���X[�x�w=�N6����`�z���`����=X(5+9�S ���	��V�f3��6�Z�cV����
A/M���f���;�=vF�!��">+F��}�V�uw"퉗����h���^^Z�������i��XJT�V@�1&,��]���j��y�6̑вr�P��ٲW9lN
�!��y���a\��c߇ �.}Վ��pȈ��pC��7�����<�pę(1g���m�~o��Kd����ȯ#ʕ�3���S������9j2*�~Щ�Z��"=[Zgd��|ƄS�X����B��=?�H���t�=91M0_��&�n����������K���͕o0�ϴ$;[�*U/�����;;����h����s!	*=�I�M��z��=NKu�?�#,o�qd��KYn�.sFx����X��cV�c&;2p���r�3�˄F�������Uyj�F�|�����Ѥ;�ux?ˬ��Ʌ����-<d_���������{f�5:�:@���\����M��we��&�p�_��M3QL(��/V>�'+��g�ȇ��y�C������5�55h��Nmj�ԍ��b���?|����d�յ���*�Ui����ߐ��i��}j�����7��4Z��CT��l�#��0��	8�T�d'%�S�\ՙW���ޮ����.z#��Ǒ�7�'�Y<��) $�]3�m�yG���&A���Hx���\DFFq�wuz6��ǡt�&�+�9	��jff���3��N<RkV�����l�c��ӛ�����j�ܨ���u|z��P�+�1@��Q[KŖ�3(qV�mtCĀ�	Ƨ!9Z�8O�,he���HE�>�1;�c��$x,�z�}ozb�.�Uk�~�<����k]L��p3�I�}f߁��P�����`��G����Ȭ��qL�j.:b�ƈ��O�D�H	h�$4�	���,��)�ei�(�(:C��Wb�1N%�=j0�'<T6��p���`�Խ�&�ӥNR��'�n��|�p���Mp�nU:��T^�$D1��!	���&��)�c]�(���}�"�E7+�'H,E�|�`�,���k:;mBݭ����3�mp��Pe�sÿ��C�τ����B$�B�q���b�f}7[!�/mu��.��2�ͳ�'�(��/č2�n�U꣮-���[ta}� ���Κ��1~�ȿ�3X�}ی�	g��¤�9���������#� ��Y®�Q@nO�=e��+BFL��Tts|�R�N ��B�h���kO4�𜳏�WgC �bf՞��KQ����L���^,眔�����V��_���{�$���#�:��;W$n�	��M�~O���A6~��՟Yv�Dޣ�fR��G"���8L�ӲoM3 ��o�{�l�3��pѷp�YYQ-=p;�2dS��l�2��i[��&�UX�ٞ.��&�G1�Q���fGu ��M]��2��}���=��sȠA���'PI������Pq�.隕G H's+<�癵Uw�OPluV.JP���p�y��X2��)���� ��R�����ʶ�⤓�3�י�5�+��~(�\P�1��t�wm�M������C�|*��OS' ��Ʈf2k}r~�Bi��$���åK�Į����M�yLF�"�d/���^�Y-���d��<����j�%Z��1c�:@ {�����g`O�A`����@��o� �X��?���x�p��9��p|Xh���{��yi"F��OH�H��.>����%;F��f/v�捦�����X�A^������<gq���V͕�e��<���)6)
 ��Ш�>�$��i[��R���PrY.��T�fK䋧9���ɨa��n���u���D-%�O���؞̝n�C[��|¹7�G*GpD"��t�����~<�DP�2�
����)�|/}�-��&���>q~F��th��z
�3RAa�aNlp��8�Hu�^�'�3G �ݍN/��T��z�J�S����Ҭ�~�5`�b­�;�E���C�ǡ��P�[\�+��_�וTo'u���CZ��&�*g�-t`ZY��<o9
�3/#�+m���Qv���OB ���mb�o@�(0f<=C�Ŋ�4�<7^�f���2%�Z:��ww�h�y����8"����{	n���)�����q�'�._�Z�� c��� ���v��a��j�Ǳ�~�m���+k��p�pfި�i{in6�V$�8ma������bb؉�����d:N�f<��
+ �{t?�~�#?J%�t�W��2b�#�+�>��c[]2�Z.YB|[^����^I)K#U��{3z+�N	[B�s�b~�Xb.s	G�;q{o�tۊ�3�%a�������
}bpD@�2�s�*��u�*߮�%b�)�������q[vW�H{�� ; �%@�_����1M0b��3N���XhʩG�S�a�M%e`lV>������A��B�����ɩ=_Ȣ5i�pX���W$h<�l����F�?�i���/r�n��rV/��/�
��j�5�@�O~�H�3�}��t����Zutf���`V�����Ox���}qe��ʚ�ԝρ%:a��@�fC�hj�"f�9h�x�p&-h��K�v�*�
��g�n5?����!rO����EG8�ɿ_B�㧉�k`�a��f���b��\�G�j��a�¤�5!�괯�~*��Ǥ�%r�1�Lͣ��ς�b���j-
���}���%��	����ΚG/u����5�'ˉ��X����1m�m_A0X����L��;5ҿ�+�/E����VK;��a��9e~�'A���
*_���DJ���Z�m����;֏+�jr�|dQ�d����a�4֫H�՗w�~�V"�!�����s�e�(�H $Gċz�uO���O��~;�9</��n$��;��������us�>�T%�hg�ױ��ep;�R:0��4J�F����n�<J��^�΁���'�mFa^��Aɞ�y�Nx9�z/��������sf�g�K�s��w;�J7�V��9B*�F~G�;��0.�4��c��R,{�$��-��M}}����D���,^n�+f��k.�����O����8�z�\c����6TZ#fY��,�R��� )���Y���g�:r�B�I_7|9��g�H_4���Xy�n��Z�v	0S��t6͸G�GHYD[�Z�';k�,=/(R2�x���[-�ޒ���U\�T�fQ>��{pB6lƁ� ��h��);P5�.��u��zIR����T�l��ҭs�w6��!	��y}��������{�QÛ�V���hp˭���J  S%�!��mȘ��� ��7[�~9��R@�_���;"�~u�����J�(��l��I�o��g���gG�W��T)]嬖����R4A�e(��/#u�1�U���A^ �urj|�SRS�U��#��2��1*��He��c��~1ﺙ:��[R|c�q��uOK.�k�R�Wx�d���̮�޿b��k��������L.���q�,��KU[p�L�PWVV�����4]<����)�2	=Q����b���4ZFc�F2�N/�_�r�K��I�7�?�&t��c1��z,'�+@_��/D�ntᅷ����<�ygࣔ�=�{Z_P�D)�m�ld��ٻ��<W�i�f��` ��n��{\:WBz~����� G���"��kދ��{d(��3#�n�1M}Y��9������#�nC����@D��_��놤J�N��� � =�{�Z�������u��R�̍)�����H����A�Vs�^����Q�r����h�c����&_&aNʲ��&#�إ�V�M��zI�{��+Cx
���No��=$b�Tj��S��6����-��f�
b�k�3��3NA��ò��x��I�f�?���%�d�����e����3=��RN�7#�P1�!,~n���(]�RnR$3c��a��3LZeC��ߝ�v����aMMR�d����x���Kc�Bй���z7?��	�T52:�_QhV�.���W.���W���G�4�\t[���'Ե��#`<, ᯴���)8�YVq��Hs��'F�i#��;�����	�W�@��:1��;�/<����Ȃ���q�9=�8��.��N�^ �{�g?m
 � ck?p���7dȾd1H��pW��~���?��|c�+di��3{~̎�^��=w�q��ОD����P���!Ck�0n��Da��l�8�{�V!'S����|4�JB�����E�1�ή�H�A5����tk�*�|ۑcwPk�&C��5�������'���$_���<ԇʬ�w��K���Y>ZO�Q<�_%M2Lp�/�r�%Y��T����u���cC�1|��	���|��-��7A���f=r�
ĉ��(�����Z��>�;w���)�E�@/j�P5JV�&�R��l q��'��	~��� ��P���J���]�QO�ݹ|�3^gs�rx�BR�R�~{g�o%Aҕ�wQ^	�ˍlI����?H�N�����ܘ��q�VP�.�g1���9�:�{9:lö)\��,�Uno�.j�u:N ��k�53�VC3u��`�>�º�'��T&����z�
���2��/�2�i�k�y�~�����41T��K^]X_��a3��u}��s����r����8Ijo�c�3�����Z_�R�������b6(���R��:I�&]uҋ�%+��{��Y_+�����>���FR.ޛ�H�k!�[�_RsT���I�Kj׺�L�hb���GF��j�/��x�<T-�$�ŗ����!��(��D)t\�(lj��M3��ļYX�<R+�?bu�a�gN�\���;���<M<z s�Ê?]N�{ק����7���0�+��c{�u��a:Z�%�o�S���;����8ݿA� 	�3���Yv����Q�ʥ/.���v�c�����R��S������ʓ��p�W������֍��B��8�`�چ�D�"��8���Oܬ6bN��E��T���+���\;~����-� ���qh�:��aԃ�D����𻗳���n /�4^�B��5�X�]g�Ex�{���c��A�>u5YA�i:�v�C����S95u,;��Ő�������|�ke���x~�N�� ��z����&Ibq����(�|����3���$T����A�{�j`���� 3F��ڍ�?JJO�_�Ro���Ŝ�t�U���d�蹍�+�����.8B��;�H���9�������[v�B�y&��ʱ��ެ�ޠ�p�4Қg�˲ڮ����l@��04��l�ը5�|��j	1LDjQZ/d��S��$��K��zVUI�	�!w1��Y�%X2��,�u���'��9Κ:�-�#�LY�)��l�q�|�3g�����- k�����v��b���{���}��{����N��������Cl��P<�"��;a��lV�n�>-(8���}<�a�)o��^���p�>, n���%_��t���j.���c�Uo���/�$�m`]և�i J��Z�U4aD�M��J�M�a@��;����>�	F�2�����j�a7>����E�����_�w��R�������e*1�(��w$*��A'��'YTm�'-��)P�I3�O�*���?]�e*W+{D�QRJ��@xW�i)�ܼ��1[x�g��r����hT���E�bH�P�~�����3��SC���B���Sd��x4�j�%#�,	��O8�z;�;J�W��i�{���ev7z��.���z_�YAh�;يk.����qO=r�V�;�F���J{�*u4��:�z�vP��8�E�;T��B/UAhv-6��h0W-D�6)N���;��gZ����"���3"�)�~�	�O}�$حȐ�A��,I�b�j���Fw�]����ԏI�yU�Ȁ+tU+2l��Y}dAd��	��S����\|K?�Q�:��ۘ�s��a_+�w{���m$�?�<�՟:}�j|�L�8b�ۜ1�;�p��6���� �S`o+�)E�e���ڊ��<aaY���RU�����1�E��,!u߆0�I�%E�꟣�N}��(�s��P�P�@��=	���P�C�4���ci�uőW�Дy�
���&yj��*��qGb�w}��3�q��C�*�R��"b[��ȧ�e.���>��F����+�%��	~ gbɡ�I��'��۹6���d-.�դ�JHmJQcѺ��8]l!\}�g,��	�j�#��?�SyG �/eݞ,���n&�����[Y��'Eѐ�4��?�b�[~gi�4���ƙ�B7�l��wq�ޅ��J���	�2��ǔ��&��u7A����`T�n�k�W24 T��yØ$�qob���n;���z�d!@�S`�j
��}X�_���2k��7-%�c��aR��4�A�\.Y�YTq���O���lu@A�}H�qcF�������~�`�i��7 ���%{��ZS	`���s�Bm�Fk5�VX��'��cuh�-W��<���)pP��<��}@g�:$� �ݐ����ͤn�r��è!w)�)0ke�M;b��X����=h �|r� ��8Cpz�?�]����|�ӥ$�5`�����ǽ:Lx�L��v27�@R �s���������k�FD(��WW(q@�<�G��Ϙ&�w/O��r����`���Q1��dE��37p��0�K�f�$ͼ�����k�X�������
�S�ַ�!%��gӆ��?��:Tը��.�ǧ9$�[��s����+㭕,����W�6��&��	���(l�Xz��-}u��%hb�Y�ȋ�F��P��F$gj֛�7�-�l1p�W����y�������]o�f����o>u�b�V��e�������S1ޏ�զG��o����x齦}mɕ�WG��{�⃺
��6�ޖc�N6����1�~�՝��U�jJ�b�4M�qR��Ɉ���@3=ZƊG|hn�=zYV�� 6�T����[4�O��_R�9�y^f�L"ʸ�C��\����O�`�cүJ���p�n4	
t*�_ux�Ht����QN��a��ؘb!3�l�&��vB�KN��z��a��Z;wv2~����aE��7�����:�p]��8P�f��X��F$�R�t*�����c�Z~�:�|�)���O��*�Ѡ�~�X�d�{�*�*j6F�>]{D@�w��
�UWU<F
Ņ��Y��ƫ)O��z������D:�&�Q�wA�Q;��<\n��W��M���U���(���`sC���o�s�;a���^��
��}��9u�p'8⡮��E��<v�����Ab�����)z=���腢ͳ���s]�Cl���s-�E�xYaܸ��R�}iW@Lev�=keg+��BO�w������'������6��/,��������2ݴ� �JXpZO#=}M~q&L�b�� y�*�rN��]�R�O.�3Op]cg���{�T|�qـ��P7#��P��� u#t�:�u�O��?�೽y���2��_��Z�br��Ɏ�g�%,Z",��ZCB:sb�����VM�p33`���X��/���@���!zSNjA�D�!ߒ���5��S��|Ž!O����~������&o�
V����	�>�P}�І=q�a��yLcq���<�3�Bi_>\��{[O�gf+�����}�F���K�k9s��"ŵ��u�|T�Ra8d9*{
�t�u/x�7d�~;��2�����\�Q����W;��v���ܨ~MQ)�9lw��"��JeV�W��@��X�L rQ�Q��뜣}�tN�0��L?Da|\\��(/(Z}�8<N��>��b����p��d5��s��n�n������aD�0{a="���ր�Q����R�-�d��p��X�E�*��-���ws�$3R�a��HeFً��4`zܺIf�T���z�[mQE[`�мQ
����0bQ|�*��T��}���kw�j5ȇ�[���θu�(�{�� �ʤb��c0�5bz�&g�����2Vc���6{(C���J������o݄Ҋ$h%Mc�� h��P{3��/����*�V��Ô&WbU`�F���i�Y�\��ϕv�A���PO�e\Wᦫ/-NH7� j�0�����8}x�S�n��<��Еl��OQ�Hp��!#�4Ȱ������7�:���OXVoO��k�-O��\A�K�S �WR�dͱJ[~=�x��E�J�f����<[E8���F(.d���,�� �L�~���xq�n�E��Jn�>W��h����wgP]�z^�B��D����7�*�z�Ԙ��oż(lF�a �Ӆ�,�-k,ѽ��67���m�}�sՉ�)�$���-unu�D.�����+p�#|�6?�����`:�G ?Un�e�D[�E�Cu9�������rDTBH������y��;ͽӪ0�'(}����� ���L[�9�����aݛ����מM_Og�У�ܘ�;��	nϔ���L���]c�"�I[�y�of=��?/^�5�=i6����%?'��� ����=Z�A���qt���~\Q�KV[�ڠt�k���T�EL�N ���<���FċQ�j&�^��%���L*J�]S`*����N�!��g_��oB�X���������0:!מ	��������?ld�wRi�A���$���c�$�-������������ �����G�5���z6����s�@����7[;\G� D��/S;8�]�\Q��.�@=���������z���D�.�&�ɘ(����"�q� ���i�]���7���;�9�a=���n�6����_aT ���,`�5ν�c��`,g�g-��1�B��_;Le��T�$�5��M!_�/.@I��hs�r��8��XL����۬���k|ƀ��������R�̤i��Mt�dom�I]Vi	bN���}���o��P0C=�غ'��V�(����S �mt�r���'��ۻ�p���	�I5�^�to�b9&�!	����B��%u�/�[Y ��	f,ۊ�f'S�C׊�����Gp�Q���](��;O*biIx��Z��@��h&�~� �P�g����e�ڑ�.��ҟ�f���aʺ��5�VƂ����8S��P
*S���d��P�~�r.���z��K���9S�K'~�Ƌ��n��5�i��ҏ;$oP�����4ݫy:�=Vb����v� ���1��	'�dn���y�~�w����M�ǘ������5��"�b��5�iM�JW>1���o��b�8���赡z9�F�̳V1�v��ʱ�Lq����$"�{*�;lPd��l2�Ő��?���C��V-ߋc"K��_��5�x��i�>A�F��V��1Jp����������  E95�=�#WU�(p�-��V�ӘQbu&Pt��p�,�ڸ��d}k�0T��%"��&Y@Cϻ�s��3k";����Y՘� �|t.Ӕ�2Ȏ��i��CY+���<�%e��'�_ �Ky�Z�q��̚���ͨjao�f2nk?A����/i�����[��o��G���J�?s>/N\n�q!�x�L���u��;Iǐݙ���L��y�#���%��%z�}��#I�g��vLN3��F1�a��D���oȴp����+�"�D|��^�G�c� �TUrb���ϴu�Y6������|��u�.�&F��q�H�<��N�
��C�k�y��EW�8����Ct���k�Ms�2�Zk�1dd�IWM|��`��q�7[q܂�ߞ����G��ȽU�Y
E]���Ziې�Ѿ-
m}}�:���q�,���L��,��p�'�'��G���h�����
&���+�Q�gH�Y��=����/���~3!�kV���%p|LE�O?�^5��&�7�!7�d>㷌Y�]���iu��5xm��l�V��U�r�Qg�y ��AlF� 跾])cܫ�O#�&�����Ot�:����MJ�4-v�\U4[&��R��,���X���}cb�	�H*NbU�R�I��V������h+�Bd�5�d�Z���k{���Fj�q��eRۺ�X�j3�z �EC9�Ǯ�����K��\z������Ɏ�����T,x� �ЩyW��de��͠�%V-|;������` �|ڬk���y�H���6C�*�bQN��}��aHWj��M���K�鰴����?YM���-�������?4G�A��fz���ᝃ���yO�_� �Ѭ�a�`@�Oy���,��B��U�����hqʱΎ�\��O�T���߄����FZwx�@��h��ڰ9��P�7#ÿ@�4T�]^�ڲ<l-֭�@*9��M�O���Y}:qa�`�l�V}fq�vh�z3�"2�!0Gd�"h}+f+��!#@��'���>W�xlx��c-(+z0�Sɴ;�̧Y���{�D���p$�����.b!# ˤR�|f���۫C7�h�e�1�@�[
��2���sz2"�����n��]zW	��R7�r���=�I��2���b��v��Om�,��c+�n����S���z�Zb�W{���\va�J��-s�}=��/��U[1$�ޔ��J{p�����U?��A��:�~� ��5�D��K|��w������Kǎ֟n���+��BI��ۣ�R�6p���N]��ʌ=��C%)�{�I�Wk`���/f��)Ȃ�]}W�����b��<��X5 ��������B@�/4�(���_��ެ��_4���Ʒ����S�(�7()o�������A�d��,�eZ�GLW�ioI��\�m܏]RC��Ϫj�ǱiA���,OVj#Nc%��sv���|b��E|^�d7`���j�^����5���z*� 2>��l�xUP��$]�$7�L�brq�f�D�s�Y��ݑ71
{���jn��F���~9�H��M�ӗmsJO�$�QGtm�8�j���0~*�!H�<�.�;������ K�%{9̛�3����~E�+L�̳�w����SH@��;u��S}"���%۝�*H�=_�|\=�����Sv��H�'f� $hä��W�6�.TД�l����r�1���+�l!�m5�I�Ӻ#�ɴ��"|8�GiE0礆�d��$h��B}���6jQD%׭�Z-J,����7o �o](k��ڱ�Ԯ��T��
t�nO^�8ϙ�Į���b���&�n3�͟�^"�(��X�^���Z&�GϹ�D�mKҔ܂����6��}�g��(Y�����a�Ն��A"AG�!�C���!�\��d�8�d�?b��f��`1�Y�����"	Z~��0�_2|VjY�}R1+�
�i���0w�������ͬJ�=�������[`0-"2����	=N�R���g�(�3���q�tk$,��1/�_	�TR�E���]~��/�x�"¢*�=���c��O�+α�N <tL
�u�l,��H"4@���I��~j��~S�~�����ZE���g2�s�R/��	���萲|���m����B�	�����B����d�=*8�B�q*�H�5�ٯ���er��	�α�?�:oKi���(n�"�A�Ra�r��o�u�_IݞnFv�x�q�s��z�;���4�3V�&��b~tk���lC�b�b��k�>%����	��.`�Z�r3k<1v}��J��L�iqDƭKc�l�)��X	���6�ش_x����d?�Ͱe�|�rO��U��������k�j���c����~�ׄ�ϵ��f�c]
�ѡ?�tS0�2��HN��EvVA=��	D�nW������Gy���7��2`�Pյ����rz��'1c��g�x0��p&�p�H:ޘ�*	�WQHt�a�	�s���ه�����܄$h=M#;��Z����ki���gz�䯍�jX�Э�5����I�����`+mp)�Ov�"�S�9!���Ѣ��3��8<*����5���sT��؊un.	�]'t�$̿	f�5�ve����,.cVV�%�� 샹��~���Z4�g�%��卢���=�%Le�GA�����.���ס�Z��%/z@�J8��������;����C���@%�B��p ���埑������RA�(֒XaF���v����'N�;�W�D�y�"�������#����X����	�
L�y��#г�B��K����q�?��S:.V1C�ύ��@ԟl/ձ��� ���nR���:W�I3BіV�+��Y���k��Iu:�lm��h�=�� ���!�ص+

+z��;�c��#J�P�B�j�ג�\�0�s}4�*p��\�e�
�)jfK�s6!F&�$5��f�n�btR?4V�<����7@���f��bX��c���pU�%��Nƅ�xg?~V'"Q�%&��}��2I�gs�5�X?H(F�}�fQ�]襵0���i.��1�������i�m^ʥ�K����7i�z1�/���p2x��K�좁�uB&7��*U<�)����=���s�*��A���oi���?4��N3�
����}��y��?��
�鯊k�}i�.]��Ay�Q���Q�>q�\�i��][z�w�u���/|Ç-�T�@CErM�u+`�֬��cyB�':d�>������Qc�n���KtZ���ty�S7`�'��#�k�Հʃ�>Uڌ+���bg�g����(�v�'߯�oe�l�x������x��b����7I�ܱ�:�gO���ܮ��~lRs+��:��0J���u�ʕ���0 ��Ϣ��`���;��]Q�:��1����ߩB��_Z��>�w��ꊀ0�bɨ���KM��s���t����z6,p���E�0T6��4�36��!�Sl-��!r�R��~�d{��fx��N�fR�
y�,�	q<�"�[b�o����P�-5ե�mXi�0��_�Ϋa�E�>�M���c�Bv�m�-��\��E�C�!�A��F8�e�ϩ��v2�f�|N��m	ʡ)ؐԑ�8I�$����W�T8ˊD��)>i���/�o���
�q��ԃ���Q������'F��\_�0di!�B+��Ơ�X7����i����X�Ͳ��_�*٪J���*�������%�����V�Һ6���MaRJ<<�2�gߴRXf�L@/aӁN�)&���lj6u(>����r
L�"����,g���}p�M�ڦ����b��~��m���N��o4���
b�Ь<aK�״l�Tp	�K�x?���T��H'����w B\�K]�ԧN��PD_��]�+0W"���+��(
�h�lY�Y�>�wׁ�I3�����B��8��S�S�5,p,EP�Z�uAdI؇P��(�Ehp]��,��0��H'�s�n�w4(�!�Ӵm�����d����9�q};J�+E��-kzA�-�_U�Q��Ё[��$Nf�iU8�T!�4\Z�3j�.U��
��ɽ�<	�ݬ{F��5�gg��~p/��7?��m�ܺ���1�{%��Y��tOh!��_<P�9�����K-I����\);��٩�}���.�Ƞ�����Y,�l5F�բ��~c�;�0	��nE��ߕqo 5d��k�3���Ql�1�GוB��䔑�U�c�ap���{gq���x��[GO��>9]�y�E�[BA���Zi�(��.�[���\�e���@z)�ӧ ��1V�4E����������g��8Y������$n�"6n�QT��S>��8����F������?xԪw�>wG�Bl�30�Q�+kP��M�+z���v�hlQ�D$;W��;���IGja<���va������;X$Do�z�g��y���L?�0RZ�I~�aiBlנ=bF�g�c��Te���&NGh?f�l�Ug�)l�J��R��[�g�En	/;��r�s�/�w���t�U�B���M�$����(���@��2�=��P��DiIU'QW=�F�zt����?6�C�I�{=��[� #�J%,�w"{�jHK0뙉� ����T}��ৎ)f��m�òOP��דX��T��P�R����V��5�H���m�h��~��@W�̔8�ڷ�Y�ؗz��&�0��	�f�q&���'ܻ���2!�Ä�/M��~�*p7ˬ@,�*`�gHnڱ�H!�CGۤv��v֐?�J8���!��&�A���ް��D%]�w���y������gf�o���.(�|�,\!����*�ɭF���us}DA�фro�oG���&��	�Bp�4�r�o*vr��w{����D;���RH�U��A��T�b}���C��yP�VZj���ݦ�������=�N��!A.ft�7�IQ��}��H����%����窖M:ڭ"Oq����I�Oa�z�����ϡ#ۀ��g���ʰ�nWm�U?����LrGߛ��>sa?���mҔ�%$��)�=s���Y�c0lD[?�r�ϻR@��� y�(n���������6�_�_4�U�U��j�����":�hf�6��ͨ��0�:��d�u��q������,�5+h�k��S � �*�v���ڙ�q`�W��2�V
�_�sS<&��jb�\��ā�����"���27�x���u�����K>.���y�<��Ғg�w{x�r�>�kn���'����Z����_��Tf���Ç�G�"gOVB8���r���P�Oxh��,��\�-q����BҐ�A��4R�#�w��N�2� 2Ih�R��)��!)�Sj=�) ���%� uY1� ��W#R'N�_���~��P�(k7�)��[�b+�~��OJPy3f~�zX�% �%������^���F�=�[�'[��"EO^�dk ��ԼN�pP����ѓ�M1u5����D��&o��7��*�߇s���!���3w���G�{F�g����yڈ��-Ly��o�� �YL�
���λ���_����ϫ�3�m	Lsw�Μ�F�,�ū��������>�3)P^Eo��<#�|y��l���>'�W� )}Ú���VH٨���=p���5�J���¸��f��
�Ś�As-�H�l�a33��_�l���b�ɵC�����[; ��_?k�1Ks��j҅��=X��v1���Q�<� ��+��4q���B'LI��	��c�x�:c�]d'��_�a�JV�=a�W@��n
Ma���K�'�$��:Z������IQ��h^{�v%���\t���h�fF��,�L��o
�q����46�?9��/x��=�!�i�)a�H�����O\��nO��8�O|��+_K&����m���)�C��kK�7�π"U��U����cA#9Ď�3`�4�8���s�u7@�̈́�f�|J�弩mbj9�&!L��F^"�W �!����C�^����x�
vl5���3ۢ=�eD<�*�����H�q,3��������U����]�H$���u[�N>��uV��`
�`6���C�>���3��[�����G��D币�t�7�O����_M�=����:ĒO�Ȅ�[9�%[j
D�H�z<O�ޛů8����$>%l��yCOԢ��f�ɓD����!c�b(��~�7|9�^`�����8��;g�%Ʒ.�2�<�F��:��<��;2��ߜ
WL I�8MVPhW�����?Y�O��ND�jh��������@ٚ|��i��k"�X~
\�L�����sX6-��������*]�&��593V��)����
����s�sT�7���[�f��%ͷ��a�a���nJ�g�<��.m(��*A����~�u,<s��x�'I��_���$4�h���*�G��E���.�3H�_���c�+O��A!����Ŏ���m��֙��YF-	U�	��)�9�ȂE[ǧ��\��	�;~�-H���vᘻ��w�a�wKho�Pn��.®=�#�.X�8�E@֏r��K&��y�-�'����N�?f�9�gD�)�HI,eE�I/l6�q�Cb`��7�<������4k̛s�Yl%T��8=�<��ܵf�W:����%���'	�O��?����焄-��T�H�5��x�/7h�J���:´����+��O��'��w����:�y��S"�o�]lj�"y}!]�~[�m��-�I0���:�8WMw�K��9�h�JsG�ͼ����&8����c9`��A�W���К���Y�x76kѧ����I�\�Ȑv8Hbw���yg�A!Ŭ��������e�BU\�i��]ލ
6��_S���*�TY롅�5!���r�8���<���5� I5�_M��YV�a!	�{��4�]��5N/q����#���,���7��oc��?fՠG�́�d.v��v�M���X���r�Y��嶈<�*K�H���s��3�>�~�o_�Y�a��5���#�����b�;=O�0��VSpĻmZ�-���(4�Ba�w�0�>�Qp�\Wٲ;�tv�\ĝ}v8̾�O7�=厃?]���"l�=X8��ٵ�A90`!إY�N�H�Z��q'��,��'Ֆ���kU�̶}����e�I�{?�x�mk )�αTZ��4^���mCmW�4��z��Nbg9ɉg���qES��zB2S0y2T�2۰�D�����x݂�<܂b5-F{�� �og�������7$ȶ�������6�Bޓ��� ���;�-sF[m;���%�`Y��[ϔ<�Z1A�}B��]�0��,i�Z]'��ˌ�t{]4Mm��R�lS� �DZx��%6�&}�Z�2i@`�oᑮ��l3�A4���Z�č+i
�[�]���pã���%o{���e�QwMR����9�C�m�I٩s4����ּ���1Kch0��B#ܶ�L�	EV�]*�.�[��YY��nP;��aw�<�^%�M�z�����ZV�J��8���C&�  �"}w���la:�O>Qt���v�pj�(�6g7����!�#l��o&��շjsU�Q��n/eX���]u����Z�\��4% 7���i2z0��}�T��F���g����C�T*��*�CG�e�����(��9y�[�P��F�kr���CiZ���J��V�xn�g3_b"����c4�1�`�Fh��C��!�>����ù$�U�Ԕ�o�f�T��}�q���>�_��[fcVX�{�)��>|*�a�u8=(H�p�H	���KJ����ߑ  9�bƝy��"���x}~K�-[�sK�<��!����zȫK�9�l��g���S(�?�`0�:m�����&��\��r*�$��$�]˦e�cmZX;����_�SS�0��j�gQG&���R��ǩG�OOrI��$�Z\�[	���x�(�^m}�p�B���Pm1U�	flᩂ����~����׳��-E����_�-w/�0�����g�LY�?�\Gf���B�TL�K���q��U��;��b�c��Rܾ���MS&yEF$�:�5��S1��T���0"���.������[��4��>5g�0 Q�^`{TNY�#
U��N��\�r]-���~�5�xA�74C.S����& ��/R��i�:3���0��
�,�޵+���Z8��l�Y!���PW[��i}E�Ն�l��M��U��~�	�U���ZiBЮ#OTȇx-���^�l(��s��:c(�:�Fcfda��Pu'4d���QL�b��ޅ�Ra�zd��x�	�Y< @.Ҭ���P��P��I
ׇ����uCt�����	�=���!6QYN�/Eֆ�׹�B�LU�뫕q���3ر)�"_����M���rwO�����+N�agU,�@��+��Tsƀ&75-���U���1)�7G����'�#�$:j�S�-�KӅ��a���3N���%�1Ww6qqԩ��ўI�頬5��*�JU� e�Y6
e�T˹���z3y~��nH7�2I\�".z��7��n�X����}��j)�q?j2c\3�s$�~���7+s);�V�p@�@�Td�F�(g�&��U����۳I�o~(��`kcZ`�N��CN4�[���č���D��ߥ�.��9��y�x]���ƪ��d�vSZ�lVIGԤ(�Ϩ��kQAz��F>��ͦL&��>/HCN&�1Z9��	�c�$��i�r�咄�FR�.�؉���v���P��n�;'��O2X�F)	�#�Sލ�ںM_�0���<�ւ��yO������:����1�Tu�l��E�_dPnp	��IT�S�eHARR��d��]����W��'=��*�Lan�u@(��;���;�J#�@C��B�<Z�@���Zud�$fOu74�/����7�t��O�UH�V�m�Z�V!�����-���9D�����y�Y��d��']`�{�B1�,�[�S �ra\�l�r�BI��3)̮E��̈v����@�t�F;9Ym�C��������.�7�B9���{Hw��l�����Sa�1fuJs*�G�\�*_&�ht)�~)f'����|�o��+gt^����ӭ!�c�d۸ED�٘��=��O�(�����OYg̋&��=��-3)���(7�*�L޸��AK�1�8r�	K��}p=��sTsnۥ{Gn-�'�+����l�d��D/i|�Kc����j�[�:f�,ˤP5ŖO��|,s]
!�88���v;,��S7�(�z�������	K��V5�|â�!7�e(9�h?�IwU;�´�/QQ���LWkD��Ƌg�8/�!t�U�T4b�bPAf7�����:~hS6��j`�/���.\��~���D��� 6��w�?���\;����hX �|عr�@�|��+`���VI=[Ƞt�f·�A� .�>�5W�����b����+���r��3J�ȢU�~�ʣH '��p V�~-P�	p�����;l0*���-�� ��^E�����9�9P���
�Y�.���)
)�%¬˜�ND��A��dh.����Sm�a�x��C�&-¸���		�Һ1J#����84W�}9��E]���ɷSу6�]�c�)xv�84J�CL�@^h��i��4��,ޔϰK�m (�|��Ǚx>K�e����L�-0�D���fi�g��C3�f`P),�3�e�-!5�U)#E�_��Bټ�՜�{L:�02<�*T#��W��Kj�	A&�gF_8m�L����9 L��p�0�-6�'cj-��Mmh%)��9�v�Z����S���jB@�-��<5��Zt+9N<pg�4H�=��ݣ�&v�³K�dSI՘�oR��P~�
Ƣ��j��s/X|? �2���IaMj�rт�xϓvD(K��ǟ��^X<m��da
��p�@��t5;/�A�E<�)^�~)�>�������y
����}Wr�[����r�-gIC�{I��o霶�3�7�rW�A}z\���qx�w;��,H �2cUNeM��b���J���d���`�EU>��7�+���i��X�Bu¼�𑢃L��2v���7+�#�vXD���\3��~h���Ҭ]�y�`?�@?!����o��s\,��'	�(��I&$��ɚ�U�(��m�lLƢ�b�~�T���{�E��׾J���u9 >�zx:k��l��ߢV�����p�ZT�͓�;9��n7�]�T��ʯl&����uk�<Q�Z���#eE~p�:F�F��ӡ�Rh.3���� ^�,��bsA;}��A��(���S�6*qf6d���fYCZl?��i�� P4�	]x�H܃�ן^����5�ch�_�-<�+hD¾ql��h������lp[�u��.6�{��V��N�+�Z��g��*�I��ntF>]h�����bw�D�v���`�J�0W]k�FML6�S�|��B^���H��i~�?ř��Ѡ����n�Y��T�[	�p�^Q+�ၼ���9Y@-����/lnvr��?�rR�L8��)��~	v�9�)ލS�9@VT6J�r�r�+�Я��Ԫz��<���8=��a�q����x��}�e~8�e���˞HNVr���6x�u���ZTb�&�_952��5���gV��!���4x{%��=6��ˮ�i�Cų��^7 ��֕��wڀN���Ah0�h7�V�ջ��}y݊�z�jVU̡&���_S�����A+[uJ�Cx�{�c�/�������
4}Кn�E�����<G���'a^�L�V���[�w5q5h[0�@�`�~�}�藥/!W�8���k�ݸb������$����<<<�*�~�<>��ns��B}kq�ȴ�]�v�y����Mo�e��:�%\wO[6lnL��J3�!V����G/Dԁ�*�0�����]��'����<�900��ˤ�l���·�-Ѩ#m�l*D*�kQ|R�C�AŎ��G�1���11D4y�Ѩ;�����.v�_�P��π���J�Xg�����H#�т�i�\���W�>���V:Y��3`i
�ʩ���λ�y?C
�S"�`�7���f_e:�� ��fe�Y������>���Mw�_�H03�����#s�4�|�`�7�
�?�_�%����j@��	�Z����$�j ���_�{^dO�k��`���G�٣r�&H`���+��)�Dj�O�諮���u�=^|=#����N�($���v�҄u��;��tАRl!��z�p����0��p��}ν#�<��8�կ��G�Ӧ�t.ގ:e'f���� �A�'_D:��ϡ,7�p���؈��%<o�)�a�i�M�ػ���s�al�,�z�A[L�,�<w���)���"�og�9?�g\����{��K���^��l��B�{�KE d���Zq�jA�f���������	q�DX��8�u�(�X����9H�tNG�I֦�]0dk�@j�S�<��-l�&�,�B�H�D�����Z��$��5�;��ӶC�!�+n�*�,�/p��C��t�r�v[�鞻�5���km��)��yWI`�L2'^�v���Gmû>.��pG��%s{��倅Ȗ�	j"�3<](�G��?�z�� �ׂx����VH��/n��B�"�l$�7"��N�֩�X�sk�|�p�!��_^n�䏁Q�悱�$��j읗F�D�-�>�����Һ��0�m#q�`�9Ab9�"�7���O�������3t��R�PB@�{�K~u�ʤ�).c��v��˻�E���^��4���U�,}�u��͵m�Xin�a`͆?�*T�1�=�EX�@B�c�Z�q#)�-^�@�r�̔pF�.^'�5V���1:�|��@�Gy:�y.���ɞ&�=#��`��m��n>-pY���8��n�He��ߛ��u�(�M����R�	���YRH�l�d����>�	(���6M�iqM&�3é����/n�0 ��:}2;1��ll猷�(��-ɖ��DJH��	�� �� �,�{��vY��k"���3xR����N��P8�$O� V�|Ҋ�;3T�C
�b��W�D�R7]o�-��:c�v.(�[=
&��*�e(M�R��x>����kV�m�a_��+���~�f���hn���jۓ���D���[���P)�!����������y�V[�sW����RA���%H�0u��1��a��e�^�Bf\���$MH�7��S�����7��$s�xk�G(b-��\���o;����̞Ϧ���oc�SD�%+Q���;���Sm��"���͕)�	%9�S��j���J��kѨ@`t�vt�b�stդ�S�@�6�³_i��6��2��,��DvA/_��E������k�Ջ��diH�EF�s��Mfê3,�l���d��&f�I#_=u��qJ��+�1N�t�CI����gb�$�F�Z���}t�䂤O0��A.��|aT%�]������5`�@Az^I�v}d�c"�<v��8�B/�e-���2V6ۚ欓nTx<��\��Zy�E�(������ؖ��lZv�(��/fu�+�W��t�k�J���m�W�v�3E,��Q��Y`���l$��-E'� �l�X�f���Y��z��	y��v�K[�C�$`�i
�	��]4]U�Opdv��Ĝ1��S� ��I�l~��xt�y��|�Y����;���Dړ�O�ۏ�:�(Vv������ލ��d?"����99�Wf�;�*�qؾܴ��Qfo�9�l���OX!ĭK��J����	���t�������qT	u�̐�g��˔{]�K�4�b�mU����9+�/.�]W.Kf�)g�Mwż��F�%��g�����s�hXH���Eݭਗ��z�='�K��AB-���;���� V�: ��Nh�o;�bd�$�Fo����}5��r��5�?�vۉ�!�5�|���'V§	�8[h�]�@\��6Υ�
3%�l���s+�<
y�����TϷ	��L���sPy����T��v� �gd��?�7�K����ml��|�%'�e7�>q��(-x2J��ʞD�������_lm�a3uScf��.x��Kɡ�'�X�%"�U�S��:�Y�.`�w��-��R���-�F�C:�����n�y�? (wK�y��t�a��+,0OxMaݮ���#r�k��L�t�s��/Ұc��͇E�e��"��?�5�K��/���K��D�H�5��,�hO���C`ZF]�G�C���^N̫
�TN���_Bi�b����u��4ꎬ����#�f��o��P�V�֛�{��T��#�Kr���aP�
���#�Z}#����l�2��}L��5 YC5���b�$�U��g�|�Q�~�n���[�ីm:4�����?K��>��
")z����i���l�NoȺ��C!�������I&�~oY�7�b���� (4B��BU��4��c&����u h�+%X����ä�vbA*TCI�=�pp��`�zhV��w=��<�ݠ塶Dl��вd��e���CI��d�����x�ڠ�w�K�������^��ՙ�����A7U�J�d;~��a�"�i�ԫ3�ͨ��g��q?[�q6����<4���G������i���"�.MR���8y�sy��&����-����i��Q��rY�=�H��0�
��1/:�k���L�&�`�v�B*�N�B�f��"�����g5���+�j'J`��:���c�5��1_��l��:zP8�KYa�Uф���2Pb� �� )�!�T�W�xz&��:�\���(��|����͹���_|!�^*#I銒'��,���]:��2�j-ϋ3'~���\; �X�-����̞L�ڣ����;/]*T]"���xcއ&�kUϳ�X�p.�o�q�hN��n`YF4z/� �E�h#�^�4}зξ=�2B6���N�y��r۶ԥ�vz�kj����!Ѵ9�V�z������m ڍ�I��Ӣ�[[�Ň��'�`������v���p�p@�,��lIoؤb��!�Y3��<��OD��і�4�j�{E��Ի48B6�1	��$#U$Eg)��!>c���i�BT�v��%ݡ�½�O��%�eI"��� ��$쥛�
�
叝�6n@|{�E\�w7��`�1ml���I 1�޻���u!�řTЧ�	p����}��;!qD%E��X��,#��/ Y�c��y5mi��l�f%f��M��c"*� VWǄ�r"c1;��Oh��]dQ���M�+,Z4�#�@�	�?��}Bp��U ��ƍ�?*�n��t�&&y��m�7fT�) ���ͺ���>����O��`����O*y���n["�6��,EDL�}��J	m�E���F�<���_�ۑ�Ș0�ڂ�w�s���shX�|A��E?�HЬ��AZ'�H�8�V]�g5P|��&���
E̋c��I��!aavϠ�I7�.�����xԜM��?D&���z�%ap���7��#=�Ę�C��֠zN(ޚ�w��T����G�Ώ���= �_5{���e�"����Q�r��|d�<�B�!���^�K1�N�[T�BW7��r�����I>h�iH-��<���Tݥ?��!�7.t��8C�dq��bƭ(�!3%����`=����'h���~G�8yJ cWC���g9�xLA�+P<�-,@�1���q#ӑ&$2}1 �IT.��fA���}��4-���` <t��X�t��e���5_��(�#`�$U�:j�66-�1/�[���W�T��m���vU��|&Y��c�;�BYE6�c�w�o͡�k=]�sf�rߞ!�/��\�&7� ��\�d�����}~�;�.X�Yu�U��x��b�����$<O��(e�,�<�"���C�\�'�,̖���F�sNވ7@.i� 539+{-N�E�?Fk���ٝ��GaF��jn�kM�u��}-���HJ~���K�)!k�w�F���r5`�F���Ѭ	 O�X%�I:oLAg�Y�HaԸ�`�U\A� !$ef��|�а���q;��Y@�����CJy�����~�N�bq�	�z���wV��rS۽���Ʈ,7��_�5��A�~���D�������z��J���c����!3��19�H���`�|���
1 mVD�軻tS��!۠�=�"Qیj����U��j�p��>]
[�K�chz�m��kϘ�ɭ��X���ҏk���O��O�b�ҡʹZ�$Sf�^@���L(]�	�fX����F�̯	 �	��<�:�%��0��;y�6��No��|8֮��8A���'�:{�Tr3{�iy#���
Z��[CF����@�bZԭ���G�&�$:Ԕp�f��x���Hh+��[uEq�-*�/�Me���rs�*��7��h��!9��y�61��5��Ʒ�0�qM��q��(_�jnO�Njn4+�ˑ~$�-�jؼ�@�8�{nzZ����c��d6�x��9U�w�A�L B~�%��꼰h�A$�]]$w�sRp�K�y*�*���;�tm3�ġ¶���������`X�P(dJlI�c$� j����/����k��F������͊���K(�����N胐���ʐ
�f�Z���ɸ�Z8��mxW�-��P��hf�	��"�O��坋:�6%�^cbvv\y7�%Fio�J�2�ne��T&���QG�C�Dh�!T7E�m�a���b�{|t�4������G�ck �r���9�)$d�L:����y�i�9���?3�6�t��O]>�r|��qr��ͅW;�K�~O�v ۑ]���C�6t��%R��n���GsC�01�h���AS�^\'���Y��5Y��B뮢g0ٿA':k�n�e:\{��L7��鯎5"͋~Ew�X�W<�Qa{Ht*Nb=�@l�d2����XU�m��gSN9���;L"'���`h,ͬ����5�Sl�R�K�E��v@�����s�7hU���`� ^vA�Lc�ă|�q� (�a��5�3+�,�1m&y�W��f"/�����SvHx���B
�����,����#��Z+LV�ÊF���I�@ZE6�r�y˦�/Q���_����t6��Xܵ�jL7xd�c�/;)]�/Qaz���%K��@&{�E�kn��J�Z��D(�$����5���ֵ�\n�6 ��7)� ���>rq�.�Cqg;�Q�J�+NO�.�r�&4f�7���p�̱B�%���=�ָ=2휞�'Te�꧲̙�I�$��3Կ$�����k�A%� 'm�2�C�1�tU`?}9��I� )�(VEx[n82��FPpk���7���<������Ʊ���x0F���Z4��������Iꔺ��2e�!hX���g0�H�50�%s�d�g06{�~�3Ǌ-Ģ�/�`2tr�Ѝ��ے�B{A�D*;�,P�S��'o�B���G$�(�$�'Km�l~�Nr@��:F�H'G�{T C��q�crl�C�&C�R����*F 4A�y�u�9V��Ӗ$}���>�����U? ���;֌�B(�D+-h�QN5qzV�Ш׬�"��E-�յf��ڿb`kB�b?����2���R��x��<*ىR�)�HS�ؖ���ӵ������҂X$L�޵_J�V?gF�o�!�|�i�U�J�n��J#�*���s+'���J��� ������v`�}��]��ذ|��F�����(%��Ȋ~!��/�״�CXw����!%j=�}Q��Ǳ-���w�nU%k=_�$̱���8�����x�VY]�M`��/: �I�|�lj�
�ͤg��ںʈ�JQ��!8��Ț�@����;d�:�Pq,�\X��y|q���IYi>0�-F��f'�]w���%��\(��M�nb�����\�*K\�#�����ʓ8�%�� �bٞOM8
f�S��#+�)t�yI��h�R��Crȗ�$���h恠��X1���D���l�K�Y�a�L s�{��$��̢3���Rg�tX���>���nˉ�Īu��k}�{�!"�f�E���:@����R� �Pf�/jO��}��f_�������dwsWeeH�-�$���� | ����ރm��tS��H�E1ߨ�Zn��J+A#>V����6�1�1	d��Z��%�������������#.#ޮxo./��&z����)���"FJ�2���6��h��:�T-'�إ�"�?X��,����z� |n�0bO9��[l�n�Z���e�)�ɁsV��W�o+�ы`k"ʫN��9k ��웽o<7��	Q��BRx�O!x����;��R������/]I]�%�m�$\��M=��LP����,�w	)q�Ԝ�g${��t2BRpR��ޗ�4�L�hd�����71�>�m��17o���Ӏ�6f�#�iGq�UVո��>��|�t���jE�0ͧ{w��kQ��k���\�1���~=����ݢ�F�lsۛ���ށż?�;ad;�VUo�S�-���v�ƫd8��g����\���4kc΍�rxQ��?L�q�em� �_�� ��N�� #��+,O����N	J�o�=�.�����ߍE�#ݠ����E���o�a�:{S���o�w���$#���!Cr@<[9���K�\}��f\V�w�O�M��ʔ�)�P����o	Z� I��ВWM������#�!L�/!��Q��X��G8BfuBC�s�K<�;)=R�C�O΂lr����NB�(���\q�z`����?zI��f�z#D��.�{L���J)�������	c@��5D���
��H#�u��Gx���
����*?�5�i�5)�TN�HQ��bI�l�(s��$��V�(�p���1! �vD��f�L���,��P�sʠE��fZ�b���z��tE}	ܦ�s��0�t���m)��C�F4��j9���\yW�;���0ʝ*s��2Э�E���1�o׍�Ф�v-3Al�wb��cga��0َlgN��,�<۔� 3�����2�91]heٰ�!P�M���t�Wo�Y�:�E�x�l�ງ��D!u�N���-��,<ޮ0&��e�ɯ��;EV�y��b�X�SW#�Y��!���;a(P=	��'���:���)�	w�X�������0v^ex� ����5����K>2�_�N� ?7�k	���:p�/J���JN�b�� �N懝�$5�5�{чc�_m".�^dCa 'u�^\�ȇ���¤�6v����SaX)<E2����W����9-ziw��%&?�E֒A����Xsy!��-6�ז�uӮM)�dt=�J�2H5��<�-�v��@�5���n.����F/4�X���C���gh�шQp`�vc����˕�Rju�I"��mŁ�c����\o������� X#P�+Գ����3�/�e��P<��M$��U+�r)^���
b����02���U��<�4��hK��ϾU��������M��;�S�@>WHx���E��qCo��C��p��).T)&r��s| �Q��L�~�,�@u�����٦�Ƀ�2ͦ��৔���i�����~�Mury|ٙ�5��׉L|7��u�d��ט�WFُ��l��p ,�m�������ϙm���A@��]���ʕ���Ͻ��B�Q�no<���=�yJ��O���+$�,�#���qR�%fׅ�FF~�Ӑ�ј�6ͨ༺hT���Z�u�Z��Cz�KH$��*6p���d��O�3 y�!.����S�r�͚��㸑IV���I����#��ra^��u�t�>��eF����� x��5h�}D��1o���}^���8��#�܍P��w�ipf��t��{Z��׻�6`J�I܎@�[e�Sc�C�'����$@�rW����$��+�������(�$��`�e�d��uP�
~��&D���KSW�H��A�]G�^&sA����D�ڂ�FV/@���t[TvȄ1^ �[����Ψɒ���p� ��<�2��mKVڶ�Y�}t�<3h��և�qq}� A�b|��{�����A�A5���dz��9cX���R����(��ٿy�� ���(��!��9*R��=�V��q�����o� �f�?]}B ����;f�f��Ъ�����y���ˬ,g��w��9��*�5�+�v�3�v+�3}�/�1����_Ú��-��ߋT�m���n�\��
o�A��  �84h؊� S�������\*�������_5gc�
�~���3�Z�ʣ5QP��-�H�^k�`ykl�fs=@˂ò�T}!�L�ɱ���5� ��/#�KY�2����u�R�t
�6М������6^����#Ѷ[�/�\`�,%��
�V�����[K����^�ĕ׵]4��&�Sb���0�����^+�A{���n���l�t���e����7ZIP�btnʦ�np��(��m&~�3Y�l����pt�����s�"����U\���q����~IE(���6��Ă�$Q�oS0:[��B�þ%_�r�� ����k� �U��&�{ylg侷��K�M��z�w �`7�K��t�?I�PP����滵�����m���l�wE�� s��L��q�&�|ՄN&9$�L NZY�(St��AS-���w�7�M�f���5&��!�Թ�C��4��r�73�T/�4+�x�
�Pm�����`�s �@a�
�t�NJ��j��W�_�d�����|=�ϑ+~��N^.��#B)�Cd7-����.@�&n�s�|�q&�+H)�aҏ��CC �>~ZZ�����l@����U���P�}�B_$	&II¾��1Յ�� w�h��߆I��]9M t�+-e^4�D�L���*��aa����"R5O�����8D��1��6Rf�׭l'�&�C^��J"��b���n!���%�C�]�j���2�Q�c�qTU�1��a�
�0�#C	�|!Ğ��?I��I�nb��, �
�?�Y,��Ĺ�̓�D	��	j8�{oi*'փ�Lќ(MK�p��,<�G\��|_'o?Z��ތid.��H�8=�o�췡���U��/X�S#�r��A����fdE�2�&m4�8�Y���㷕8�"gG�CZ�u���&��^-�C�����e6�,��w����J5f::)f���@���:�*����=�H���J���������9oF�ϕ�.����-s�i�� ����ˁpMIc����D�+�M���T0Mރ��Ҧu����u�'����G.�#����Zi{h�v8U�]�����bEY�s:�,�7�[����޽*��u#��`�J�ڝ��1Vs�FTivW�x3d����Yc`@@��ூy2�DU3�����m�Ϊ��afî���b������e�/a�]�Y9�"��:Q)���)''����},DG�K!�@����).U���AV6���'�9=ɺ֧�0�4"F͍�����gj?������Vb����e���i�'{�� 5-Y3�S~y�����
R_�/��m�ja���K���HYB%��}�gh�jd����j�+��m�x�;c!�`��[k2an���[����@*n}�'`_�-P�W{s͗��>�xv҆���:����K��}b2g,
�N�Z���Ś��4�_%�-^�E}�oV������@��_�sYϕ6i��&��;6Te�m�� �(���8�܊��"){}��a��E��{�)��03��"&O�4e�j���o�Jm�:����������C�M�$E�/;����[1ݛ�xuΜ�Ws���s�z����/��h�]X$ m^<z��·���'�W��I*�/�e�ʪ� ~� KDZ�q�f!�'�ˀAn��Z�w -USȮ4���C��:k=��C(=��W���t�o*ۏ�p�bOHOֈ�aA)M�Ogtt�ۯ�
lK�
���9O�l�H�UFy��y�����M�w@�0���|�������"�S_˅�J��sԨ��Urv���#�'�ʤ=M=�c��n����	Ӑܚ(�>5g�~1u_�z�	�t{j|��9� ��A¼e
�^]��+�.���o}�3�7)�Gg>��F9;p��ݩC���p`�����ׂK�*���C��z����6�X.��2L���]���7^@�C���Ľ�s"��P������Ţ�,c�O9������*"cHRH���錠��� �L�hHWQ�b�/8��K�����0&q�.��y�K�~d�R-L���\LI�810�F$)yL�a:���I����4$<F�X����	��e�Hn�\���!L:l5��>iKZ���A��|B�����7�d��6`��|����JH�-"O���b�v�#���Y�\H"�f�O��8���͉��9��'�PaѮ�"�P��~�����P�ѓ��%�A�_��7=��;b|6T�Q��n��9��Q�]�(⡋{��U��/>zb�/�*Պ*d��H4ʿ��|���E(�8��4�a�6u���;:-�cԿ���Q�b���ΔN�u��� ��.��A?��A�4[=��=!�B#+����E$d�{�Sa2L�L�e����	�Hv��