��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~�O�qs=�  HjCa���-��M�j43�9HC�:�y��~ܧ����	��f~��Q܏w��*N�"���zX�W�7رW
�<�1�k��ǁ1#,��]��D��@���>MX�Y�[��G_�y�^8�Z�ӗ=;?G��M+ȿ�
�l���Y�If-��¾L��i^�2��ds��(�0��"K�c�kE*�co��q�.�յ�_�ˎ��8Deٴ���+52��R�r�N��&��_����E\���U�?A*>����@Bj��N�+%���+�ȖEs�ғ��!��1�������גo7
P'�	eN�g>k�=}*�!�B?a*�'L���$#v|��7���e�����/(
�����	MRe4���">��c����%� Q�j��h4EJ��|.l �D䒁�<�0�6Ju,�)ؖV�u�I�����?iϠ��oA���(8Ka�������Rn�z[�I�'#c���键�n��n`n��?H\�;G\}U�6����P��.�(��)B�r���0�m١蟨;h���p/9Y�H����wk�R�8n�
�l�
�f���w��A6h�յ�".5�a&��׈z��(����ք������1�k�Þ����^|w��my|��+�+_�;s�G��\^��@�J�6瞃�֬_螯F9��e��oAH�)��5�����*Q�;bL���:�2ä�̔7�������Wt���j^Y6���|y����w�OX|��M��[Pؠt��QfG��r����e��lB��4DX�P�ilMŘ��Φfʘ5#�;�sq a��ʔ?G�9ï�a��Z~��̝\�k�wõG�c*��D����Έt� �J�n���x:�~ �j�J�iy��8��O`e���yL�	XzF�T�!�|����WR�5��l(Z���������;�{xz� ]�y��7.@]��`"E�>��B�#1<]�%��G7�T��"��)�@��5��&Io��>,,s~����{��(t����]�ך[q/�س4�����c�B������Ơ߂��ډ�ŀw��2/���)<�z��dǚ�@�$\�ӈ�?���Vz��ڋ߉����3z';��$���4:3�%b�?�%M�CipM��Q�̬��j�����	:���zx~EwsN���1�g;=�L�Yg#��?��������
:��<�J�﹈4o�XA�Eq��<�\�� Gd�������'ڋG-�Z&��=��l�}��K}]��T���	��0m��X��%;��	ɵ�Ѐ �����,PM�Ok���gfh_NS��S��`7�|���5�g��<o���<M#7��ہ>�$�0�䈕��)N[��Z�t�g��vB4��9_�EÊ��wx묁�Jm�$�29y���� yt:�����|0�K�J�9ԋ��m���	�چ�>F��.�~0�����f=Z��-�yG��5EC�h���$T�/���a�[�jP��ee�	��D��k#��h
g��$2�ҽ����Х�ȈX$�����)`�"h�_��{�}l����:<l*	�4YGM��S�ihmK% E|%�������y��E^`&�[=�Ů&y5�O���s�>TYB����t��1�!�a�d�W1�J��#�4��|d��8�&�4�a6�H_m�y�(�[� OOo�������P~�#��w��ωmJ|i$+���6�wk38��*�s�KQs�I��3������WYK���n,r���d��w�Ÿs�����GQY� ������ͻ}˰=��gIIS��ۅ�v9�N�� $�)|�#*\�e�;F�b�+�Ȍ/:��Ӎ6��9���d�%���ɹ���N�_TR�ݘ����s��y%><��Od����"7蔷Z;z�=d���P����p����B�����C�,�O��PU<�N�rrg�T�8C��~��x#�4q|��� Ǝ&��Js�( A�*��� �@j���Hu��~�R3�xY�r�14��Z��8��d���5�ɮ��%Zտ�U�x?�K����pQ3eS�:~?z�d{�p�*k@���pR,��#}�j�m�U%�I"��>nK��#�e���rn�0�������h�F3)=�k�����%"��
z�n�"��>�ZU��~O%N�j� k���)/��qk���1o��0�x����=�٨gmI�s3���������)���l:�%s�+<�˃�/XY��@�J�T��\�?�F��Y`�96"������ 3��D ���e��Zo��5zH�,O��-ZS�]��W�M���Ƒ/,^ueO�A����i.�	�$��^�^qߖ_��W�巉�88�S�p\���w�?-�1��Q8�|�3#.��ӏ������É�cD��&P����l?hd��|_�ߧ�?�^6h���a�C�758���_������^�	���B��|���+A�L��qe�����d����P�+�g �m��IŒ��y�E��l?B�v>9P:�H:=�ljc���U\�<6�������A?�����`�\���ۄB�]tx�N�0˵���k������)�ꗼJo�������1՞��d�����s��ӊ��?wL�%�&2�1x���M������T��_ϽN`9�o�"p̺΃Q�o��2t��a"ᆝ�Z�@2�!
�a��!w�c'����G�FZ%[.���@��Ƭ�(�/<�SQ�d2U��q�� �h��I(��~EJ�����|QQ���n�
n"��e ��#I�X�z̙4���_1	LkB�p*�^��֨$��8�Ȓ��n���("�'iݷ��Q���ڇ[�|W9s�֮�k`�C�)�z,e`E��m�Yuǎ���?C+:ؾ�=�0&����= �x�F���c�����d����9���P�|��jΆ^i�'r-,� 7g�<���N�U�[�y���P�1,�����J�0Lc��:��Wh�{�$'��a�9�g>�����-��{� H�nw�[5Դ�%���h8�����.�nYa�ࡤW 3��R�񜌗�`e, ��j#Q\[ۻ<NT�v���D�q��I�u+-����ĄN5���������=`Ύ���oà���I�&�%���G�
Ƀ�:�=�0�L���;7������C����df��Y6��x8��ݰ�xFi�7DύX��tZ�>���k5fth;͎mKMM�E�N��^Y+�|V��ʳx'���R+i�5i�@7u��v;��b\:C�i6��KZ��U^�poE)�3�n]]�"1ȼ�OV�����C�9dd�;�ۼ��y�
fÁ�✾��ţmP{�ڢ��Vu�g�aC�xȍ�Yb&���h����-6����B"�.��̼���]�K�K:C%M����If��z�Cę�g\c��{��Y�_<-�\|�V�yl��(uW�WY	f���L��f��s��4��}�+"�S*����֙]��H��gE�h����Lҷv�fS��Ҳ�q+R�}k����O��~�a8�Zc֓A�i�E����ISW�\���\�x��$R�|��뗺�n��7%<w#��k�|M��a���}I�X�r���$}��["V���:�]K��1�BM�I���1��A^���ͫ�2����S��#�iF��z|�(��e����no��A�b���,Q�]-������ꨧ�6����AX���%�YZ���ğ��E4�Ǐ���f�`?D1D������B�yUT_�2L�Z�/�):YV6�3f��n����n�i�2y���(u�(���J�o�+}�U*���$���C�Bڣ�\ᰬ,i�Ś�<Aegْ,#�o�Y����Ka��1�v6	�s��B���d�6dЊ|�]t�g��I��xM�����/AԢ�K~�_��/�N��|%Fg>�E�iqQ��4{¥_�i26��cj�㹻���2*?��W;�܅���&��!�a�v
��V�P�7'�㳀C��2��>���i�:�=����G��hL���T�*�D�b[�^� t����xEi���+�[T�9p�f��p��T4�*���D?�Bo+�sof��֢�Y :����A��\�L�Ekm��\���N�1�y�삵	&��W4 o,��LA�v�l{���En�V �}��k�)��)ȳLkr*��~֡��Wo��'��l�ob��ܼ��c|�CW�;o�m��\����lt������r�/y�KzsO�J!ыV7�,�`�l�%J�/|B���{y�U��7g��)5�3��;eٞ��O��,d֐��v��2d�& 	:<П��=m�&w"���gMy�O�l�@��	Ē�)wtX�od�Oi�Ɨ�X4�<�����Uk{��"�}|f�^��C�܊�p��ѷI�(6�������Ύ}��]��u1IW���	�GR��K�0��يE���"7�q�Ї�2gc��[���߫8��2�w��9Up~�]����
K��t=b����3�D��+N4gm�d,e���1�}��l�I8���*;��F�}��̈�z���}ih���@Ի8�L/��e��Y*+)6��S�o+ؚk��� tAr��^8�����z��'�&�6l���L�2��vpk��/�{~K��
��`���&�-�u*��c��6݄������ysC4q*����Y
8E�A�[���3�/�[���'�R�8ȗRz[�J��7E���I�b|j���������d~��P�T�-T��I�� Q�ؖј�A\w��7 ቍ����F@���.��4�N,�����"�Ϟ����!������}��R�1�Ꝟ�nTI�����X��9q�#h�M�6g�E6Fm}���'4�R��-����^��Wc��B��?� ��-ix�`[7�7D��{9ih	�$&��3t-�Ҩ5Wk��D4��ōf�k�n�-�38�5�s���o��_��l���
�	�룀�[���*
��ű������o^�1!�u~G:,��ʄ��n_avJ��e��=���1���~�A�&�L��"���׭���=�����D�EyϥN̓P���N�4?\H��Ew�n���6s1eg6���1�������� �'j�*�E��{��n����,�ª������]�<o�2]oi~�%G�&�YC�&��hE�PH�[�^s�����9[����sM�g�#Y�8fh�y)"50�t�A`j��\�w�BI뮁!Rv�yAFYگ���k�fl�H�z�*`p�e1tA���+e���k|@i˱4�ˋ�,�ڍ�8�[�'C�)9�-X��Rv_�ͽ��,�¨8�n넽x�?S0��7���]��E�(r�b�/��N�r$��+u��Kb��s�齚:�ӕ�Zn��{�Y�P!#\#���FO��~��0�{�����+-ɚ��+�����K>��"��
[:!���p�E8�vT����3�f�@���ey ����ۘP$��@�y/]����U�� ڝ�$���ܨp�eП�֩��
xj~�װ�!��1��uW��A]u�[I�&�Z����`��i���p��M��éL䔂,���X��Y���<|TX��VTl�?H�\�!g7r�:E�$KV��q*ț?�J0$L��QMĠ�k(Ds��|�;Wd��ٿ�84淕h&�Ъ�yF}��p��W���/t�׹�R�VA>�R��KJ�����2�RO��b��8]h�ÆN�n{V�洶>�bLD{���gm
8L��iy�T��U�&���^���QG����^S�Ơ��_�m����喺6���Ś�{ 56#!P�Tp�;j�C�@}Ox����II�6i��|�U������K{]ʂ���WݤQo@��U�4[�S;w�B����f �k�#�H�(�
�ˏ;���6�g:�����ڶM⛜s��CH.Sm	�$�#S��k7H�Z����C�6��Ô��f*0>��HR�$cJ?�M�)`�]�����k "�A�&o�`Ť�ʤ!������6�U���V?{�>>�Lg�@,�[x^�k�[:�,������J1�b,,ߘr�XHM�!��s��5b�7(s-"Ue��]Px�p	��ϫ�D�V�W�e��HM�b�stoD3 r��8_��j��5�5`�&�8tމ���yp��W�#�v/n��o0^�^�s��[�=^�++����U?,	�z߮ ����i00<&܄F[�E�������r�����^ݧ�]���?�c�-�|��?����+��6�aX���`7����(o�TՌd���+m��bh�T=�3ϭ�S��-i�C�o��M��W'A��n.�/����S�Ԭ/��l\���+nX�0��ksO��Rn�YlP�`+�+P������v?}BW@xD�"��X���cx�I/눐U�D�Q��S����ލ��DF&y\��k�v���?����L����10d@y�B�P�?2���V�6��"��R���<�X�����c`�k���p�%By�4��0�ޚ�Y��Uc���@����T��u-dٟ�A�}ڦ�e].�r��@�����n�3�m��R��������}���9��A���/����Ӑ�6ŕ�����jOtjR����D3�/����b5w-�`����G?�=�÷��e�#�"[�����%]a ޥ�f!	�o��R�H�u�6q�g���S�<C��R�Ҷ�!�*$&��([ ���g��IO�/%��d�E�ᑚ#�s+�`��h:�	��H�ԡ��/���	�eˮ��:�u���: Q�|T�sb{�]^�cPr� ��b!��6��F��wK9��Q��x��Gjat�OGb�L����6C�A#8��X��vǕ��D���m[viWћ4��԰�m�uy���23@VtL۵���Q�e�8J5�(̧��J���W�d0���T*Z��d�"�4[�iu��~�g�I!ʰ�����ೇ�H�k��S��B����.fPzN����Q��J=�]�{�:�6c���6�~Ucr�M�~�����>a!�����2ۊrW�ڎh.qu�#~g�$��7�g:�	��</dD�R�t�� >P�&�	sފ,����%Z��B�y���1��h�I�p��E�؟��̙�f��'j�kd��(�w��'7V�T�Sler4pj���,!s�Pa�k�	G��O�qep|{4����-�}��#�]�]������`�vK�ܞ����~>��XX���\�C�>�@�1�Y4�I�88^�T�GQA`��g��SY��/�Nz^�C�s����=ꥭh&�	V�G�6���u~'3' KI�4n�
�-]ȭ�K'BmSHN������_�g��(m��Vo�7#3벾�
/�E?�im���s����`�`��"PCl<��;�����0�Sjl���S\�a�tL��� W� /B�m���8*1.{d�M�_zP����7B{ˡL��tp���xYz Ǟ�2�m`�s~:��(nL�ڄi� �.��j禤�~���&K���;���\_����2��o�ʷr/d@R�JH�BU̜�#�t|e���t����#҄��>҉��ɣ��;��v<�,�o�&���S��|D֌���E�i��!���p���B�g�;upڵ|��2��bc�~w1B灝�g����1�<�~	NL�����r��g(��?y��4��8�G����=I��K䔬7�ve!:1B+O$V�8�^��d��f�G���p!#t|�������;IWe/4���e����������!|�j�Vb���dvt�� %��l�������Z�w��S��)�
���3j�R~�;�
u�Y��K�pWG|�����v!�C�߁�vϚ�%r+���#��-!ď��:��|�`�Th�Ix��k�� ���N \K���	+M<DJ���qpͤF����0�N���Rh�s_�>Ҵ�%!M8BxX�齝[�ˍXB�22	5GJd���� ���,]0��$E�������>��@z�Xw�6�?@g��(S�b�����߇$��]#�v�qX�����x� B6�<�׊/.�W�#1.b}!���5B�O 1���?�(�%�D��ݻ# ��7w��;Ʀ���U����ަR쫕�0��R��1�m8�=!:�4�IAA���C�q����E�
�
eݣWZ��p�F�c7���I
�2��tP���\ �_�L��q���#T�3G't�H��BYA���B7'b�DzD'x�|�t˨7uڨy�)y���J�{G��yֈ��K��g;J4gx��I҅�7V$���:�o
�Cv;m�#;Ȍ��q�U�`AEAHR�ћ49e���L>Y��7nfiJ�}��1);{� ��֟_χ�����'z[ћV~�g��0�6�4���,7�V��9��^��掜���B/C��.���>�N���|?nh�ÒC��N'X�:G�#��ڻm�d>����ֺ�)A�D�ɵܸÎ��z�G��Sw�����H�w��Nө����_V���M�A�D��M�h�夋=���g��^�����	3\	ךͅ���	��O�\K��Po?��z����O�&�{�J�t�=2w��q���
�,1���Og��d�&�L$}���[�Z3�Oz��Vbh��d����2�=��&�}>=��^͹/�-D��z
>������(�9�X.V	�|Hx�p�����ީ����q�O���'�� �Ejl�
h��g������JJa�Kt�c�ܜ�ɢty?"0!Sh�62��P��T�.:��Mm���������O���zѧN#.�>�S����[S<cA���|oI48(.��}���}�	b}jӰ����"�S����7�4����!t1�7��U�W��`mL'��y-a��]ف��d|5��0�o�O�.�2�����C�\?d2��g���c�*z�6ߚ�'b��� @$<��<Fsú��J������`��'Ku/3N���\1wc�U��'D[v�y��� M�.�<��}�p��~�w�v���.�9�7t�I.m+-��4���֍�&RLS��������i�#��ë�;b���J�{<�Z�M֮kJ))<�b���"�Y�Fh�����������)=f�\o�Xp� �H�Ps.���jEث�����2%y(���x®�_�hk��A, =��^$��K�ɝ����;�p~�kN�xd��?�	w�WA�����[.�[����4�Z�)�%���@mF�����v��[:��7nd&pc��ǒF�� �d틥�����U�V�y�\�2���;��������z¨��>s9ȮB�U���-�
�^
.��a0(Q/p�ppk���}~rp���A 6_fO��Xk"ˎ�?��u�#T����\<)���=
����)Ҏo�s@�zBg���|���2��	l�P�E12�P���`�m�H$x��<�B����{�V��=�ܤ&ľ��n��{xe�Q;���RvQR!l=4h	�4֟z%�����ד��r|����$�y�l�%S��A�p<&���_�W\���>�H9��V&s�����Z �qr��U�}GP�'Sޭv[[I�!����)��=W�@%9z�@;2l�m�wsM�\Q���D��M]�Q��ٳ�k"u��-XB3"H-�IMu���4�gl�
�����������G�o����H��)��3Rc�~b�5�-�J�[<&�J��HN���v���F��
D�N��s�[W�8�N	>^د��b����n��͵
7ه#��tI�Ý��;��E�\��[}d}�_7�3}B���|�^MjJ��b�X<P�Τ�V�u�3V�M!��*�1+�h4���n�$��vs�'0  S�kO�P��Ѯ8��7�m@�P}	�Eo��T!�o�l@�p�B����6�=�~�f�ͅ;���s���ų�D=8�W�gEJއ9���W��� �%���k���%��yO;�f��Ƨi]���A�s:ئd��Q4���N�so{�5�Rc�Z�{��-��Η�3 :�'�s,-��&�zTe���=ߣh����2�ǡ�&�`�ٓ���߯�6�Q��N�;�R�3U�O����a۲EL��<��+5�e�������$�0����q̔Wm�������8U�+�ut?ߛ����K*���τ���{����Q|p�|{�h�����ϳYO �_ta�j��N���,�z�Z֬@����|������q�
�ϊ�¤������j�{ί�9���zZ����6��D
�g�sN���~�����z�I@�g�b�yZ��c��e���s��e(ܹX+��=1�ٓQ}LU>uF)�dF��n�Hv J�b��x�.^OT� g��'��o��X�N>�?pQT}���0B��F�ijډ߱e�����L���UK��wk�(��]�Ѩ�3Y����&Ŧgi�sG�Ң�f�aА�8��_9�t<��ҼM�Ye)v�J��ȢfL>�P�gTU.z-Qa�,��v%��\oŞA�T��SJd�e��6��uvEta*����E�*�6���v�Tp`�>�'14uY
�ž�K�O%�,�� 4�^:A���Ľů��Qw8�fy�Ƚy�53����[�ΟY�H��(hSl0T/��#�I��7��l�-l�u���rm�&:�dD�ζ�]��&��B�O!8S'�K�;ʜ�9n��,�ˇ��瓗y5C��*�zeJ2����ql:�!��jO�6Y�ƫw�W�@X��/�B4�1�K�"�H-�7u����6pҐ�$E������t��E,b_%*N��� a%X��_0��O*�OE�`�4���t��\���a�:
-R�)n��	�Z�����Y>��"�?cW���4ޕ����ka�h_�S�K�=�b�*u_��⚿��J���<B��L��Թd����q�i,��CJ쾕�z�JR&����x=� c���?�����d�J�W�vO'M�XW�o��V�ŋ3�~�(��GQ1;���ne򋚠n��2�>1�&�zx3�Z��_%O��乞�G�Z��[�ji��E����C���f��m�P��S�m)��×���>L�	W0hr�~j	g�uA�߲�-��wSpA����'z-x�">��
�%F�߷<�\Us�*z�<���
�< ���EQВ\�6�V����FE��$�B~H�X_z��M���|g�۩�@�[3gɽ~�I$5�R��	���"�"m-�h����!�fr�|���_	JݢF7^7C{�Q��px�B�B� �����,/���v��f7#	��j�-*��;�� �R{�8)�}Tۮ���ŪE=f�5�P8{�㑫8�A�غ}�N��s�/K��i+�2��\�!�d�E�ɦ]�%+o��X)���&�,�A�m����n׺��再�ؠݱT�t���Q�_0k��O���YK�Q�}��X���M���d�E�T�N������0�׏�%Z��y+X�c1��>�c��\��
_ L|A�e&5���y��u,a�\�B�́��g{ڈ܀M�W�̢��s��J廯��D/P��rz�\HS�q�!�@'+�Gè��;ȀQ�)��!h)s�Y��L�-H	*���5�(-t�	y1����jf��� nw��G��+�ѽ��3r$�&Ƭ�ĚРg�vclF�o*�%��stQ�7-���-v������죽Xc�<��!��(ͳ~�ɹ�!]�4�N6b;���%w-n�q�H/�~���M����X�b�F%(��s�qM�9�O#�X���Wf�B8� ���XC�+�4S`ǍJr{�'�R�ŗ-��.�
]b���ːP��@��i�u�A�_�E�rn�>gV�P�����lcZ_�Y3ˏg�D���y7史��6�<�=4���en�*��2i���R�W!���S��:O`L�N�>�Jo&&�_��Q7Y3��nV�i幭ĢS-�a
�f�������E����T��؈Gn�j3S~�.*���}�A����)H�H{�x�c:�դ��Tk<��w˵�/<s43���'�˗�F�+�}(��W�M����)(d�cH�7�>�����@�f>G/���@T˵)���^���`z^-�x�[fn�qX(̡� �1W����nU�|���oQ� �$��l��;�OC�#�������u}�]�Fi}*�sA;�"����S�����j��T���԰���r�ߋ��Ǯ���4�Kd�|�+#*��
k7��leh���&�8a$'c�T�.�6��/��e�K�j,�sH˔d�_�nc��{^-�ӪJ�V�i���~pTofǮ��y��cj��c���3T=-�%v�Yb�`1D��α-xx�u��⓳Wf��,X>(]	���2��"w��_ �nQ��rl�|֗�l�S��ɭ��i,�:��vl��r�d�/��S�J8��@]Q��q<��I�"��KP*��nP5�,�+�ؗ�
����������F1�[R�aJ�x^���3{��s�b9G��p͑Z�n��ӆ-	�MW�RԪ���;�9����?���i������*�t�Rl�+�Pq��Ġf�y��`�B(�<4̎U"���?�ޯP� ��wh>�Y��k�s��>����mi乯Fn\L�^K�N��u,�����<m�ν�����z��j]�"�xK+��:��aͬF�K��EZgZctw+iO�2=��/����q�c��r�w��X��f�C� :2I��F�����0x�n��
r˿~�΃����b˩j�}��@j>eb�cl�p�e3��6�T��i��!/�"7��umg�ҳ�ӿ��IjƀR�L��]ƈP	��������h��p�J\Nhb@D!�X�v�]�^���K��Rey(��t��=n�l,�4"!f��������ڼ����{6��
<�
�� �RV�l�����F:�&u��բ�.���dU��=@�����&d�P'�#�"�;P�,�h���'���҉�ZWޗq>_�[�Lc��tLv&��]�/��g�p�f������-%��5��*R;���o�1zW;�(����ÝN4%c��dovpw�Mu�E��Ԋlj�^!ȼ�����/���\c�^[c�>�ٶ�q���6+^����"��ƃ���V'�N�+�e�KR8����<��蠙#�v`#Qy���Ƞ� ���՛��7s�Dd'M�B���夈���Ds�0�V4����}����1;�4ܔ�ã�s�8,)�{��pdtNX����$4��t#�7PP�������������[��Y+��w�=1c����۟�_�uc@̛��a���o�}�bB#g�٦{��9�q$A�����:g�	f��T�%���j�RY���8o�O1;�#\2���
]��v�z���p�#j׾)Si�#�~����J��xr?�p�`����`c���ގz�BFG���+��=i���I���u�+X'��7
�h����;cw <��_��B'����\םa�'�������L��ϸ~���GY �@&���AԂ��p�ΐ���loَ��_F1q�5q�%�)��������L�0��GKc�?e#�w��k��y!wyZİ� �➷�4N��(!��X��(���Ᲊ�m��i����zӺ����A��Ϳ�4-�@oҁ$& �����V��ODyepk��y�^E�.V��$�e��e0�Gs�!��յ_Q|���'z�P)P���ܹ�����T��`�l%�v=V���!����T�����;.y��c(�-��f�͕���3Ơe�SN������#�V�R��&��n��~H��k�.%�Q����$砚w�=o%|h�GL	5m���A�K�Ci:Y�}�oxț�+�2w�&�Sn��5s���
�bH�D`�4s�r�2 �R�<7�ύ[�d<��(���,}�����o�����N^y��dz�[^�܃��f���uC�x�͙7�5�s���դ�Ǣ�veoڇ%5��d���
�C��U�����.�{���C���Rf]H��WX��&��͇At�ǋ�y6d��ߺ���2��ᨓ6)ϛvO-;�
v�tQZ�}i,I�3L%P�������I��n|#�Gj��U�!X�!d0`vh�*y��5�E��f��s���5G>����M%�O6��8�$_�SW��������ԬB������N1c���b�KvO
�i�Y�d$4��VH���zG��v܍Ɓ:�+�2�}Y��'S���8i��y�5NeKso��X6���ԛ7JғMBUC�&v�Ӆ���NR�@�o��}ҋ������j�'p��N�����L��{������-��[�E~�WQhM����v#ޤ�����)�={)��04G-d�PxI,}�I�{��e2���G���q���B�����<d���3-�>�AYRG��R*�J_I�X؉L	��Ç�;Q�?��u��r7kss�E���i$���a�I�U2�X��}��Ք�lჄ����R���G�%���3-	X��S�d���X�R�k��Y���A?8qƘS-[2����˃O�(	{��o�/S���E[����e�h��s��σmZ
>
w������A�U5������h��N�����b��w�[{�:���>�=�A���QA7(��,
�DG����OUg��c� ��{LF��_y��b*�l]ѭ%&&���r9��W2�p�hߪx����1\6Q+���.`y�Z�ŋ�p���
��`�e��Y_+Rs�7����8��at�ݚkw0�#�6�5K��8�������w�u݅+�'���O����l����9��nc�#�)� �ł`�KV��*�9���WK`0��Q���D� d�D>�����}T�9�e�m�}f��(�ȓ\�x�S�"7�������J�EY�2 �����_KAh&�L��Ó��n=L�g�s�C��%-�;���=�m(�DK��<1�d�$aI}�*�}����
��s+N�(���G5�~���K�S�	����Ze��9�"%|wl���Ȋ��/>����pѭA«��3S/�v�� �.-ͷP���s�zgV��C�yz�2y�J���ڻK2_� ��;y��<�p�F�z��"0����ط�->Y&iM�z�ꂢ)$�ې�6��3��9�;@�θ��jx�xc�kZo�ل��x�����&-����Gk�8dc�tU�c�ݦ�;˟�߆�|��w{���w�Q|ȴ_�M*�-�v��Q"!_+� �O��%��2ؕ�L�9:��>La�/M�9�E���"�T[�۲��%U��.j�����w��-]�r�
�&�5hj̖vl����8*�-$Nf��nn+M?k��V����Ji^�(���'סz�\��T��8�ɨg���%��@��$KiA�z�rgkQ��	����!܍�ݍ��Y���8*ze۴�	+��l������l��?�Y\�?��0U0!_��	�r-��G�y%l���� Ƞ��2�vJ������*��1���X�x0�\�-��.e�&�^��?5�S��6��f��,� ��H�f�k��;�l�a@Y��ܳoǏ�^�.�2�����$.jN����s������I�+�\�J��wT��u�7JY���k��&N���O����թ�x�7 �3ig��\����O�y��w�X��5��j����N���GW�X�|�u`.6������<E[3�T��x��%�-�BCU;Z��¼|+)?�����\_��`��Zذ�vUJy,�đ����VrC��	,�����]_���1���ï�7���^��eO4�XOae+tPBx
�I�г�^���mP�$�{�d:f�#�}0-Bx�� S�1J��d���U�����q��]�k!T|�s�x=�g�*Z��x#��e��̈́R%MJ�~�D�r )������WZ�>��`��_0I$0�ͻ��?������^�;s���Zጩ�cO�q�	El���4���2�E�P�kX�']�/�5�*G ^·c�4oGԹ��\̕��@)r���6���Oәv�(V�
��=_Hz�P�ZA���ٗ���Pԛ*U�,���
S�aġ���j�޸�2F��ة��*!�q��fv}���jKdA��6��_���4&����m��G����>�-.^�]�,���sߒUmG�⡬
��`y�ā�Ԕ��LU�M;��ʒ1�^h!�40r�̱OCO���/�K���X���t;���0h7T����A��N�B E�9�:����m�\����c�����ݖ�]'�z��1���y�q���2����j����H݅Ch|�3����V����[1UZ��f��of��%K�KL����bʃ�C=���$G�L�;�ܿ���P&��e"���w��Xa���S�p�5IMS��ٵ>���.�x� R�?$ȴ�����
¿���:��|n��Ƃ, �7�LZ��_���gI_g����eF��n�@5.fPN�=�m��q�Ƞ���D��P�>�� l�a�h�Ϯ!���:^���-�XݦM�3�v��;����8��{�wh,^uR������=����O}�>����-:�g�/r�;`�7�����l�����c�1 �l*jr���t�9���<Sy�����?��6۸9^Rp��� �K2�""�z_�o�k{|?��ލ�߹��lq�^9���d[�2>�'��X?�� |* �Ll��z��_N0&�2J^ƙ#� f�_!Y�'���I �2
v��wG�U|�1Avij�ʿ#����[�!�6���b.Ad��W�cНe��~��2�����=�d�{�rJ�X�J�Z4�&=Z���F[�c@[�k�/���}�����W�5�*U@�^����y��3c�ɢh��/��^)3�#�pzÓG�L�������Џ5����P���>�{��Bu��?�!�4P�Қ���N���N���ÒN��Y�6����yτ=�K��#�e�C���.����P�S���(Se�_�۬&A+��V"�J2�<MW+�0u��$�g�t��+�3��]��=5��5��*��c,��`��}^�R_� �Ḳ��vQ�AK��Ͱ��*���඙���u'>�G��RI3�n�z%"t��UahV����
b=O�j�ڞƦ�?u��+����iH���t�%�r���� �R����x�,D�&�0n_,ļ�=��(@�9RQ����w��| �;���7S�b��� 
#��e��Ie�W������{޷��>��� ^=��>��_"��Z.:3�x� 6Bh\,fyr�-C)��j���[{�Yfd�"�<����?a�kW�(����O�&p�F����C,�F�/�7�����M���bNή�=�1�Z��|�3̱F�����˥�oǯ�2��%�B�	E����1��}����x#�g �Y\X
�'A3�uAK�˕ċT��1���r��{Ƿ����(聨������z�RDG"���7 T�ܨ��~\��jS��Q���LLH����;�)MN����ϒ[r#d
'��?fJ�?��~��78C�M�/�����b�on���1f]`�Ё5�k�{j�-q��&�_�̝�Rg����T��#
E4|Շ�H��ʪR�}��/.����^�2�ҋ1G%=�9.a
�+n#hL6X�8I*K5�W-��Hd3�?�1�)\2�r�D���(�jCk�(�
���ˠ��,eD1/�?x�
�Ԏ�b�r�v�/��{Ӏ�3��?��x\?F�P��y�o5&X�rS�"��vX�?���LL�~_OM�ұ$!b���k<����5~h)&gm1Kb��|�>��|ʖ���H�K���V�+�7RKab���x�[�Gl��t4���E~ ��:�)ļ*���:����ġm����o@6�{Os@z���_F cf<ۘ"�ƛ��7M3qY�%���a�YC��-��vuc���4�.�A�^��$�9[�7�|
e������m�v��X�[`�m�/�@#��*�r ,�n/���6�aE�>LEP�������p����ĵ\П��-]qt�+Ew�r��Nvs[���	�h��$�҃EʒP�S�a�!0�`�������t��Q�@�ţ.*������`.C��z��.+���?-ݡ��0^��^�r��\h��C��L6m�%���^�Bj��29r�T�H�8e����1t?��b�@2�^W��+(ܞ�t4Yo�!��"��$�3�����=%�
Ѹh����s����r�>)9�|&����Ek�A��9p��,_0��+�1e薉�Bt/���-�_^-�۾H"6��]��Z��lf�F�����l������+�����M���M���[@!��
b߉� ɪ���67��x���mf�ϣ��c�m�ۺ��e
�s�!�����<l6誻0;(��!֫y�&�񆶏
ǭ� #W�a�6��Â�X@K�o�EJtY^/3��T�m֑y�|���уYI4e�?���.��Wv��r�CXӧ��!��ZA��ȼ���3ޙ�Qݓ<�կ���J\�V��z/�|w�L�7ԡ����v92sYW;�^�%l[¯J6+�4�)a{�N�O.���,�h�%�M)b ��&"kat>�/��[�k׸��&�c�����g��PԨ�6�@{�5��!��m��8�pa<qQ��tP� w��v����a��r·�&Wh7�=^��.N���jV�a���H/pϝ�e�ڌ�D4�Й��C���kc�]����r��V�M0x��Lg�k:�� �Q'�K ���P�[����2vxyc�ɝ�7�����4������?Ġ�/��}���L��Lண�;��8���W��x����:	�2x�����ng����e�
�Pq� ��٭���)6JC�#N�
��@��F���5܃��~�b ��g��|��/|6/�Տ��j�h��Y���!ZV�!��9Xb���qcH#'�ڮU2�!���ؚϲ�$���D��|4κ6��c��Gid/��Aa�� �5I�P�m7�o���j ����)��N�2�'g� ��3�|6)�'2C�E��\�d	Z���Q�d�c����_ГD�ܯ��z��=����3@�ٲ�S�r�c������\Y^hU�n��e�ي�	�����P�b�Ä��6l� xO��<��=g��2MvG�4Wt�2��N��+`����y��?�k����{~^�Z��.̦-,�,�a�>�C 3�^�J���P^����aL6����]q�fp�{9>g� �&�4�x]'J�S�0�?����F�8�\���_>&Y��Kˌ9fnr�o�4D�s�[|er�/��\�	�Y\��l8l!FiNۙ�?M|�E�~�%�c��@Z�)mj�r�j"�&�/P�HW�����V�:Z�krs�;���7��?��h��9q�	�,�m�o'
t\'����j���U�j�4��
2D�q4�w��L��[Ղ5�׽8śx���x�fi ���T�u�4-�V��2�2u�(���t��/{�[>��Ĺ@�x_@q`�B�y�h�焘���� XS��8�{5?
�"�3����9 I��慿�h�p��V��8V�Y���}��u(��`ݪR>�oI%�/�t�%����:�)іq:�&�	?�f��;,�����"ǑД�RLO��o+VrA��|@#S5>��K���r8?��5$K���M6*��4CцB��.8�&Q��Ў��^rj݈FN�~���e��q�/G�g������Q���V�.�����iu��(�������s��ex�t�_����B����7��|Q���Ꝅ��ƣ�y�AUv0���B��K��Z�!�L��dA�$#��39�A�̲�h���H8��&Q�0�gq~,�`��BPz6t�N_�p�M=i.�c�,�ε�m�����2Ʀ��<���j6�D�<p�1�.�t"�����.h&4f���H��1�y*���"���d�+.�� �=�=n�*Oq|���V�/��'ixz��٪����~��q�	�#�w��ɰ�OzrH(8�$O�z��#r�lzE��.�*��,����B[��+!�Aۀ��zڞ���r�O�m�;�J_T_����x�˭�"&J�Ae���*����������03�X�V�b���WCd �cx�HΪ���W�pM����	�/�el̩�"Ѵ��x&�$`�#0�`��l9�����Ă�tu(&��9DX���:44��^�R�$Ã�ndŕB'������Y飤��Yzg�^
睬���eo��Z��n�'q"Ƣ�eހ�V�W��/sB�������W�?����3^_n�e��#!��x2zؓ:ި�qskR��Xq;��ӳ`?��5�Mv������l�fǁ��t�
=�Mm��NA���K#�����/���QE͊�@oo�c����s�	�t��Q�w�+��]'�-+�8��0'9,���i�" �JR����JZ���`$i'���&Hy�.�����V��j���UB	�h�F2�����Wq<�=q�j��/��J���b���gh-�l�٤s��C�t(܈x<Ԝ3`��R�U㟦��.Sh��H��p�S�i͒���wi��/M�'_�I�tR�y�=X��,�X��h��0�Dt���^��`0�5 ���%Us��d�O���(��T�pꫭ��<�[��Ɨ,0�p5k5kC5A�r�+)v�����')��7,%F*�w��?!�:Q�<���ھ�舙���O/�8ՙ�vW"�HӰ�N�����x���nS?�,�Cs��zu��pW@���-5s���ٯ�(K`�y��n�4���R�2&����C�	��MA����#]�������1�L�K�t��0Q���wAxށJ��b(*r��G��Q]v.�r��k�0ߏ|s�_�@�[���i�17�,��#�rX^T�f�Ž��>�m�<Պ�B$2�X� \X �.���J��
=�#0��(��X��E��܂�Sr������=TX �?�M�Cr�����U=G��6�($*��'u��y��y��t@(qx+�4n4/FҦ��sC�
*����r[u4�P�V��[�?��x������-̣&�˂79B���V���/+�~B�$2��p�4Y�+7C���"0Ig�l��9��-slO�<d�Dʜ�k�~� ��2�A���M��ݡt�t�WF��|0��@x�Q$��
�%����Eo╆�k_=�c��� ��%1^�˨^R��3c�8��?��Q&ͧ�����%;ђp~&~�.9	T~=�}�MQ5��	��\ܢA������y����n�N}��}g�E��%x;c᪤���&����JS	�h�<��[��|]��>Q3jUdq� `��6.0�#.��q*`�_C{��k�Fx%+�T�X40K�&��,����L��6|K��B%;f�DӉ���}X���g��K�*a��T���{��7�����AV��a)�e���1N�+Z����ۡ,�ǯ"��(�����k���P��/�L�46��[Q���m��i�Q	�B����oa��^�sɯ3����?~Z�]W��.��(n�	��?�$���&hJ�Ⱦ2��zy��{��칥�59X�Ed��t�iB]Kjxk�/�m�y�)�����$-���Q��7L�-�:��~�@�wU��#��1x�t��s)�6/'������F�S������be�5�H�
]v~c�Xhܞ��T��D���CV�o�&��o�ljG/~9������c�ƥ;ڇ��Y�4X�_E�(6v ���,ӏ�hu�*>�/�c��i8fNJF��w�樷��	@`��6�b�]�,�$Wμ�BG���"�p�SLe��i6���|:��v
)!�3��,D�ӜzerV���%�z�yk����1����y�_c<8�5��KpB3��C�k�=;7!qg�]����E��W�J=^�����m#��"�Y c�g�jL&��r�$׾�����Y��]��D�/p���(*��e�]-�^#���G���'Ua�J\Bh�X�@1�������K��Z����̼_������䪟�)��uH��Ӧ߇�p�<��7Qr[(���+},��J��
�P��*� �إ��i댥D��jNXtn��aO�b��U�o�x�U��E*�6����<�U��a.��%SW�~8^��CJiBǢr rk�/�boM,@�E���[fw�-���t�Pl�1�K�IA�0e7�-�p
�$����.�g�����m�/a�1!�I*a�1��#�Y' ���WO;,���E[X�!��n�����nWZ�ѱh!�"��o7���.3j����pc���4���&�Sæ%9�!R�͠Y����H8]���	��������$FP��e��XD��W�A'�M��e>吉�2$���2�N�Th�@���k�}�$�����1�`�O^滸��� ..�&���ҖY�^�M�ă�����hE!���X�t������H�g�t���T�f�[|�Ǳ\�Z�
�F�ç�j͂�I�1�~�)iJ�H揕�sU��}JER_^O�9B<GI�-�0�4�Ͼ���g�w����4^�"U�@���%��T2����=gc
�slJ�U������.�x��z�:M�+s�x�@|�dq�>0 ��z���}:�A�)~���\���{A��������Ϳ���5��pd�l�bm�\*�G��Q+��J�16@O���������3}2szn�Ȗ����vh����hS����F���:��v2>�6��z�Jv�c@�i���z��O�MsbQ�^D$X�/j��	�ub-�����XtU�ݦ�0�@6����oh��k��]�a}��^��"�i�5�-�1�t�En?!��"�a\������S�f��o�������t�����������mh��t���w�L�gۏWX���]���\�;n2��<Q�J�ʦ�u� 3t=��|�J���QzOAe��EK�lks!bb�5k\M
j���8�c��zO����_�$`\�7�thˎf}{�N���/Β��XL}�{�c���Y�eU��#C-��� 7Q*�)9�f��@D�A�5 ���U{�k�Lg@�lVևK@�"�?q�4�w fiXGio"WK�;�ڀӎK���c7\��x�F�)����̿��G�3��T<Jߍ���}�7Ø2f����=i�@�CN��a�o6�.�|��:sV�����k��>5#*C�G�c��꿏��e�x~W"̕7 �*6�B��TϠ������9��k`��i@���w�Ϸ�r�1e���[�]n�F�*���s$�?� ƎЖԕ}�"� ����������G�m��By��F��Oi�����-�%���Y����;/���*��c�mAE6�v�k�%2.X&�|����J��s{��ُ��9��R�fʥ���y��L6��<CI��=-�ٞC�a�l���P<� A�C3��;k�(��U���!��v|���euB�Q�e&���U7��0IhX�&�B	��Eާ�̊Tn�û�G�Y!��ĩ�����)������li��f2���#�q�
�0e��+k	�`���sb�k�F�������8 �Q�j�k��>^/���q6�t��ߕ�������b������� v0��#���D2�Ĉ�&jC�o�-A�^4�T�.�s�[�z4��S�B<_��Xr�u�ʫ�(C�a�sڬBAh��	�.��Q7�/��Ŵ5r �V�Q6�=����ZS1nZvo����$+/�7�K���2�W~Q^��R��
�1%����sL 
�
�h�=����,v|}��:{o�Z�k���3����0�nob�Q�oǁ�tV��b*��E��YSs�.�+�K��R(Y��vF�
&wj�h��\p�&��'�X$ȑ0q��y/��s��I-�������^�����Կ~�f���I��s��� }VdU��;��U�+]��$��l-[H�u��d�������aɧv}����f��/�G��;F��.7j���Sy��O)D�Y2��naap���WV� ���׿~
��rD{�&�U��E���_#�J�
�jsM%I�6a��S��m��vn��j�F�$O� #�Y8�i(T@�����r�C#�/�=�����2��=����0S��9
X_�-��;C�%�> /hO�38v5X��M�Y�I1aM:�xD�`p��vЮApu_���=(���2GӎDh�����"7uA�Ͽ��\��.9�ڒ���3���{��J3Seo�Z�{{��Cß?G+2���f���&�ъ�[��$r��֥��'�Bp�sni����2!��weed�s_o�:_�i����ih�r�#��j~�����M��+���6����hQ�J\S�#'jqm�#�y3T�)�f�3����l@��u(;�*plV��	d;Uoj�B��E�;R�g�1.���+�.6�iz����0נAQ2 ݔ»0�z�m���@�y9o��,�� �z4��q�����%���Q���M��A���� ��[G�] ?�)�Z���>W	�	���W��G��^��U�~�),&�����e�v�+��1 
�[߁�m�L�{.����I}�{��b�L�k�jy��Y�41X��!��{t���*��J�@h!9M^�F/Ya�,M��Ks�[D��� 02�{����Q#"7D�#����i���j���^u�[f��#r`ߣ��^��t�@{��2_��Y��.�d'ޫo��G�����h`?�����׬2�9�)��Q�+���n��:�*-�z��=?7:$�**�
��4�b'@���K�b�hC�ʭO�MG��&8^�c5/�%�G��r	N��~?�};Ml��ń�+���[�l������b9���Wbe��%1�gega�~������!\��P����Įˇ���_�HX_����Kđ�I�|?�[`IN9t!�O��������ߤ�E������mU�	M�1�!U�9�f�4�u�!g�5^��� �GH�X�Œ��0QnD�l?X����>��g�� ��%����פ�<�R	4:��Xз��𔯠
�5�͈��Ƈ����P�"��(;2]OCrI��|�`�,��}_�@�`(�~���cs|���:%�f7�l�9�5s3�՚2{Wd�-*7D�6�t�-�%���g�y��4�ڰ�9�QL�Z?u]�<�%��8?�	(��̴�/�A�q���&�Lf��b�����f�'��Ks�,�̞rs[�� <F��6���6�����h��q������JqK��	 
���R.�Z����7�̐���`�����8Dw��<`D �"&8������D�~�i�v�FB���V:�!�\Ld�+^���K�G�Fo�7P�Zp��� �{+��cp�j�`��U�l��U���Sڂ��0�����o�|p�3#3+�3�:{��H�J� і@`pS
ǿj���!>"�.��ծ�wXz �N��5� [����f��T��7�X�a-�t�ۈ$�}
�����M�9���2�E������L[��^C3��z�҇y%�ì�	<�$�t�$9Kz�/�]��-�W��ذx�=
�V�u�?G�N��\�<,����6��		�H������4ߌ2�p�#U�_~D�:���(�`�򺈹:��C�Iް���9��}O��t��r��ތ�m)p��A�_�<z(�����9�'}�J�$^��CW��1#����*��bN!�
+뇇<-�3إ�ޏ4��� zC�g8Z�FxNi8�t�6��g�e<
}�3�w�T�����i�e����g��u\g�Z�R�)33=�[�HP�����Z�M�8�o�	�x���]�_Md���$�P�GiC�b����jM>e��t�������[ҟ�ż[��z�*;�f��^�b��z�	I�mC��~����Rg"
��r�d�!��f?&��mq��C�3��
�]���r���!CUZ6�����Xލc[.�*;u$r�"�}KQ���w���ު]Jɝ�%�t�E�m�=[��@,9���Hr&G�#�0�(��Pj�>�gy�����n��t�s0�Z���&g��5ԥ4ع��a�$�q$u��]v-�X )�����?=,[st�Ռ�y���#/��N�
R�'�$����5頍����hM�yiiXOˎ�=I��a:B��""a��R���u:{d�Q(M�D@@�r�y�� q�u���j
�܊�G�R8�I�U�[j��D߼}�)�e�}����D�����~��yZܞ���T���E�3� ��=����F*�c�C����ő?��fv�ߩ�Lgr?�3�E��^"Mc$+�N��5m�̏v]���(}��)� ���wîI�+s��h�T�	�@���twz�tkqk�����*�5v���F��6^H��o��a;����*nCC�u�Ar��8޼?�H��$\�w.��61,�2J�a�3Ne��7�v���0��Ј�VZ� �ml���6;�� ?a�i`	�e�ȋ;h��	g�P��erþ��$�sMu��,xE�y��6�d���F7`�-�?$�|��t���&�W�F����aT�q�u�,��[�`Hϧ��5��#tb�� ��ç���De&��O�\�I�7�B-�L���������9_t&�Ӟ(�^��-���H_��Fp��&E�)��������;*����<���/W��n��6�Y�ϭ�b�fTky�V���<\�K�F��vv�n�W�o3�7;�%&�+ɂ-f��o�H��OhQ�{6ҒN���S��I�܃�>{���\3箶#B-��Ji9���_��U�R���&�2�C�NȻX��Q����u֑�Yc�Q��Q�0
�c�1������#�h��^�7��5	"�1���������'�O��SWG�§�x�S��Б<V�jo��Q��FG	�2���K�qDF�(#"��e,�9�S����q���f���M� ��g\�<I"�c�p�A��b�1n��`����BW%��b(\f4��k�4|7O�F�T�F�+���o�s v���?��6��"O�*N��O�/5'YW��6`Σ�D ƛ�JJ��5O���C¢����R�B��~���sck���/Z��w]�w#袯��������3��:U��Y �Ğۄ��ޟ*])�/��r��9#���&b {Ա,��q���#*�'=�t�ǁ�B��f����z�Z�aD����@2����jƫ��x@0�mH��7~ȵ�쿵��5Tp��g�S(ױ!5M�kП�a������z.���������q�OCp�����m�9�:я�^k���۳��o.��_�9D�6 d!e�EX�7K�P�|ܧ+
:�>��e�x�l�@�մ\b�����v���g�(��]֭p��[�x��s6���)���h�͇��.l=N��B�v�1����d���լj�g�ш�[h�l����i$/��JT>l[���\�ɾ��e`�Q��<��{g=�4o�cE������C:4�����J��WUs�N�9H]I2a$/e����>lG3����N�vbS|�	�/hV���2i�^d'DG�ߑ}�������1�	�����x<�w6��]�-)�Y�J�K��x^����'y7PD�e�p�P��W���Z� ��퐺���>�{1��2��.�Q�lt��]��%����˂�b�]:2�h�L�D$	xN?�>���iV�S?��x0O�!5�8�٪����-�	K����N@wUxQ��u'�����q�����t���4��k�0I�8Vo�Ca�ƿ��\�~�O���H��ͩ��VP�^u����WDԌ�H�/�ti*UY�� i���Ҽ�2W�����`ޅW�J�������X�-\ys���2нw���g8�i��KO��ZZ3�ϟQ�f:��v��i�ō;�9D
��a[5h~���a;���|> �Ψ�K���HYu@���NA_g+�\�p�|�$�}⌃;Q�v5�
z_�$Ϥ�XO��,�W�����܂l�}�2%t����8Ĳ��}k�K/��2|��i�<�^DY<����G���e�Z!a$VR 윰��K)c���7ƹ��;Wسdcюs'Z��BX�c�� �!G��F	�۟���Pa��6���R'�EA-�{�cOyT@L1�W����:!#�ؿb�����((���'!����}��N��ݲ�@��st֟x��"����b��5`�o�"�S�3�B0���)裰�)ι�;VG���R�� C5Ӟ��4��]sk�/2f�h?�{a(�&Rk���Í�=�9��A�I2�/��v=gaA�2�,BF��c',=�ny�3-� �t�� ���.2�Y�}O������
��m�����H��#���F���#eн��0��m���Π$���3&�,�Be�bM]�e�
�"H�!�b���c�dR�!���Ow)����%M��5;��}(�%�$��
B��OJ����Ldf !K�9��p��) L���W����� 2TN&)
{��Մ끢&�ɀ�y^[y������c�L�*0 ƴD!�m����yZ�������������������|��rV�gȍp��/�#�� V,��I��ϯ@P�d�f���LJM&w�Pd1b �_�g��5~�m�@I�����Fͬ�,�nXI;T5y�ISl�2�Ǡ1 H�><��zCQ���s���~�h�!i�x�e�Z�-Q��Ӑ�䀃Q�+��H�~�/�g&���f��B��g�ܴ����%��a��Ie�I��<M���<V����!B� �ciЭ};���q��v(�Q �͹��t��t�-�8�W�L[Df�|um߼��Ri�����-G�<�q|C���UB�'E�f�ϗ]�H�� �u܉���+�f���єe�~�a�j�!�8�pv�7&f1���H�Z�vy��i��wHn�?��1��t�̊�cs�?����6�A%wy-6��/di��k�֜�:BS���������O֯�IMMyfr%<ߤ��gsyQ�H�з;U"0�%������+X�+��0P�����Ax+�E��%�`-3j�+��h��J�xQ�5`����C�X�*<��r��h=Dt��Ԣ��s]J��=鿮j����2]t�&+&�O>�<��>�s`O�Q���`w�������H�F�q#��*Ho~>XB7V�<ԯc�6����7M2l$Rj5M���i�� �������+�Gv�Z]
��IB�S��P����f)$�կ*�K����ҒT@�'Vv�����������)�p��l�&���]
(K�]X���a�a�H��� 8�a��D�3*M�ى��-$�/�b�)�.�M�3Ă� ��u�����ud��=��q�����],xr����e1�4��߬GM�����L�D��|�U�<�P�djM�_m���mU��Tuc0|0�0�^)�2'�FK��e�s����샅^#��l���7����Z�(X�l ��<?L�1JC�(�7މՐ�i~�F{��B���i��s��s��p�/6�3}��;�W��q2�P�p�@e�ų�{��Ȫ��M������_����Q�����N(d��M��z�����\�\:��e�bv��q��A=)F=\���	��,v�YzK���7��9�Z֨_i+��TAG2�ı��d��-�
fCEs����{���Z���3t�Oa���R�|={nv����J5�HO�>C��!̊�g+rr,�L���#++aj2�AF1������WC��L��i�|!p5�a銅E��i~����z�*�F����9B��>aJ��hhE���b<uzx�3�*Q��r4Ƣ^& J�