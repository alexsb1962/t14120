��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^��������yD�^�o����p6s�5�s�PV�.�nQ#=wL]�F�~K��f�;��&6��G��?�E�ȿ ��;]��P;�n�A�����J���5�=���A{Y�*@����.R��ގ3���F��}���.�,X��զlC���2���k���tVx��9����X�2��������$"t��w��hRKo{�{�ƀ m\�pI9w�((��)�i�1sQb�U����}�j��3� �x7����(����f�}�}��o������%$��|,d���[2����~\�K%^�ȴ���4t���v�=z}Ժ�ѲIM�^'g�՟9�h%��c&G��;�>sO�s�uH����s�� �������� �������	k1�����H�Ohb��J�}�I��>+���z�%Qܗ8H.D��n��WcY��_��{��J#�E�2�.��o!�2F��L}�Ӻ�^w�b����� H+ԋ}����m�]19,��&@�;��:����J���5f ������<Iu�1@�'M>ᛩ$9�5�ϡ��E���BA�:ds�z���Zs�_b������f֭�,|
��ը�w;��z+|;��4o0+��s07�5_�����aŬx�+�v�����Ƣ�I �g�%$
��l�lS�:�?��<��2G���ͤ.��F��4�,u��J[��A�81���z�5�#6�o�]��Hɲ��w���j���l$���n�-$1�!�<�
�q⩬w�S�<!pX���R�ő��E_%�k�����&�?�٣�˟څF<ڎ���ze8�KL���Xbt��Q���C.�R���t��")U?<֪�
_3�pb2��Oc0c<)��ؚ�'�jd+-f؉�6O�����@��Y���� �HeEP[+;0����`���)R����DP��a��Fjn���
�f��P4��X5��w�U	�+D8B����i�_r��س@Ƽgs���tJ�.{[졊��Qc���T�#D��naV�&�I�4��[El�n�wdx:K*���~�T=6S���������dB�s?2lW'�����Ft	� #U�
��1~�'�f����\�"h!��1@�j�r���4�ۭ���}��6g]l�j��+	��n^Ͼ�Ѳ�&M��>�|Pi�x�^F1�,e��2i-"���I�l4���{��3Փ�ĄQ�����u��D���� ,�U�I3�[����	W�-RH:(c�{��M2�S�m�S��^��",}��c|��͙O>�Y��m�h��)�����o�4NM�z��ؚ�d ,����z 
����m�RZH(��+�[e��Pyu[0�:�s�*�O��:>/��Fr�U�ѭ5,@v4���'Ln�v�K��0]Ή�A���M{���C�`�յ���0C~����#ue|[��t�o� �	�d�JI���t��/��Z�(�)�oP����J�&�#�M��,L��`�#��T�'���Q=u{���禰8�
Mk4lC��4|�'�xr�
���/=�H�/�'��kT�0~�߯�(k�*��%%^t� �vt����Ʌ�X���V��yF\��A���5k����M�?{�V�_,��w������=����P�v7/<�k�ƍ��e{��tvfK���\�����v��_.R$턄i=�Eh��QW��:�x��O9���-��;k}�~iݎ�����T����I ]��m������-218ު�&��)�@E���:����v���q80e�P�OpE���N�&�t;ϸ����M���{a��-ꋡ��=�� �B����m[��	�'�Mm	��HY��ӱX�CC�����j��(��H��#��o8N�Y����h ~ɟ]�am���;�ڳn��G���G2͚�x��Y�����L;����8y��ʓ��r6�i[`��F.~H�ųQv�i�O�Ue�`��&+��kf�׊��"��L�	g\����������"�ŷ�ۖ�2���\mvr�8:ϖ�NT�G�߉�h`���jr���p��T-��b�2Nm���a*��c�pѲ�MX?��ߟfH���C1�CA���6�|��F��и�j��Т3�2y@A2�-��g̚��Bg�$I{H��z��_"��������7b'6���/�4��q�i�/E����`C�����&9��P����d�� Ѐ;��x�s��vԋ1"���<h�Q�_x����N8���HK�R�0���l���U԰q��D���l�"#��LI���{Q��̆���G/NZy������}C�zp��
�*��4-�,�O瀸@��e<}�:s+"�d
D�&]2_����&$d786�$�yH��(K��V��F^��7�	�ó�Q�J_??|�^rF	3��eG5oG~D~t���5Z��Q8���k��y6�T�Oc��Dc�uYu�����O�j��Z|�HFۢ�T���!\�[��N&�d�_<>@�O���E_Ǭ\��"����.gV���s@�|P�v�g(�C7O��-��l7�T{���֞	K�������p�s��[,sX+���R]�nLb���a�N�37��`m�i0�l��L�׷X�Ik������o���]1�� ɦ�z�nO�g��o
�Q�!��V�q\s���?���,�"*eGV����0�q���<is�o� ���	�\2��a'12 ��v�뗵|v��w�����g׀��l��g��l�w��s��`��Ua��0j'6�U��I8G9�{�*8+!��"AHq����4 �����+��k��!���¦4{�M�4JDB����$�Z����d�:�ܥO�s�It��e 9w�l(]��J��|/$�e�˪�j�*�Z�*3
�EV�m�>}TVAzB�X�Qpd�[����
@KH ��� /�ͅ6���t����x�%�}��&i���)�w]�!��jZ�����>���}�Q�u:���I�J���E�/(�����q��N��
�hn��Oy�:�j�#�q�%*sC������O��C����9Р��5�O�!Lah�a!���G��e 
.�q4�1���@�}�q�WH���[vϥ�DS�Nw�ʣZ^�	�rh ���wQjb�+��RZ�wH��-R�\]�lW�nz�'��Q�UuO��k\�2a4�av�+�*��ͼs�^�Vr��*���l�����|��]1�W`�5lq�@�����&{-����̣�����M�y"���j�s������2_����'�A�6���3QT]�d2�u�L_�3I`?��R6���y�eD����1% �P�~P�]����w0��^�G�� �=�%�5��|��U''.��Y&U��l�Pxn]N��s�q{���L��"4�t�1���ށ�{�:����l1�Q�G���b��)t�aO�!{�D�Z�H?���Ad��7��sD'�=�Ҿ�}�G=G����߄��+��Cd%i�;��H2Y�����'d�^��{��1*ŝ�͹�J�� �!�s��ɏ�د��>'*����o"�+�u��ؘ����,h�k]"�(���S�L�0�W���_{�c��N'�� K+X���L�L�Qئ����g�1xX�Sw�K��=kA�ѹ�ہ�a@�0�t��<��D���P���䥪�UČ٥3~�߼:{�tf�O@*|��ɑo���GP���׿�@��M����#�7sp�~X:z&��S���:��H�K��f��6(��d�x���ᣀ߸�V0"��a��M�U�}嘓�G�;ؿ %W���nc���&�h�K7ؠ��(~���%�34#m�kSs��3/���_ܐN\�()m���&�#�e�\F���YX�Fnmv�49����#)P/iC߀���k����l1�L7#�i����^�Z,"���E��%N��,��&Y7 ��%��I������/vRu�ɝݨ�I���LC�M�䎱������2�<� F�C�{� ������ ��M�M�rDW�����R��n���g�oX6M�� �T�}��!a�������2��ҷR�k���V�d�Jlk�#��*��3�1h�x��B�EN ;[��Gi�G�ʗ[>��	��w?)�kvE�M7��l�bʫm���k��q�<���I��� ���eu������]�����6C�A�&J��d`�U�C/a9��E�E�8G�qvk]�}�'P�S3v�+���4GD�$�����T�r�N	�V�	~k�4�˓Gg�<���uĜg�g��g��݀Á ����k0���)��6�.��0�^�7A(0��*K�xk��eu�9��b�������ST[�6`�#
5m���UZS���'o����j#DP���3��᫏����3�P��z����ȼ<y�����E����X�5`6���+0�x��ְm#�!�4H�	���R�ZK�!�Q�&�(W�a��0  �ʱH�{�&~c�%rb6�����s< <�bذ?�@c��.Kn�MP��8㰥;H��| �l����f�:j�7��6�dC%���wx���^�>���.��_*<�j�}2P܊m7�d�U���i"�Z���>ҙךt���5��]�6 ��-% g8��7���Ӯ �X?9�:
�	k^����޷�%�an񆲅���M򲓌_�fci��A�4'�?��1��weC�G<�\}�rf��b�b�އu~���v;~a(�N2ѿ��o:���ؘ�y�p�9�I�֦��G}c ن�a�E��ѕ[s��$��T��X�S�;8y�S��:��=L�c���6)��n��EI�~�2�i����(	�*?,�DE�{à(��A:8kw�;������'���AS�^��.�D���E�}��&�y�T���Q�������`�j6��F-<�;`'��⿌歕��F��^rp7�&ӧ"�|��!�����i6]����=�ӲQ;e�5S�����ݛ<��x{1�I'��aK2T������ ������٥�(g��~ZS<��̢�� ���9��#��s�H_];@����s�m�&���=E΢��±��Z���Х��>�I�E`&u�R�������Uw^��T9��83}0=:1����?�H����ҽ/Y\]Xw�~!N�H�Y%>	Ƹ�"����_�mxLm:x�8�}���/�i ��ۇ�����Pk��<U ��W�IB|\b�ʺ�>����x�z��D��)�C6# ���z�xø.���T�Sw�I�2�N/���T׹{jԓe��*5 kA
REn��*��k, }��y~t�\���\�~D�̗�(���P>|��iJ�5�z�^� >)�a�6�J��ǲ����2ꣷ$z��&�AIe�
@60�Y�]h�2�nk1=����ܰ�A�$+�C.[��l��Aq��?+�&�к��0�IU�:���9�8��i�<
-"�g�����<�j�W��V&��"����>
����ɉ3�ʄA��Ob��EB���e���2S�эhkfH��T�~%Q6ʆ��+)ި�ݠL�Q�F�5�=�������,���ŀ�m��D:�t�Z����i���E
"^7z�ףҖM�L3oz�Ƕ�N5�T��)#Ez�[��s1L' �\��i��AЄ#!�"ӗe�Y�-���>�Y+RawH$��!�%q���mD1v{R)�=u�6�d�~t
�c�̨P��(A�����X�/�\�ڠ<N�<S��E��B ���ǩE�Ħ����n��Dō�vl��0���b�\V;�S�r��@�6�j G�ŝ�*Vs\;�;���E���co�R����5�7p<���R=�������7�)��FU.G�C�yP�ptw�`[��6WORc��-��53���{/ץ֬����~5#B=!�%����t�Qܯ��'yAυ�<�����d�L���[[��Cy�_2��\��tzC�qvrV���W4�����0@�>0�`C��w��"�Dp��ʂ�L�����&�~�X�10O�K��Ο(�Z� ���ȗ���J#�T���l�X����>㌮����}-ׯPsF�m>�Ū����vh�r��f0NoY|k��_k�紲q}0���y�E��c7Wt#g�D��as�H��i�;�`�].�ʌ���N·mj����V�n>:Ϭ���ߍ�㾐Z�j׹ތ��2��L�M�� BA�4���#A"g�-���I@�s��{4Ş�u���/J�;�7��Z<h�盏��iI�KI醻º��~��D����!����#�'��A�1�q���S��+�� �xw�=�Qvay!a�t������l�4p� a�Bt���9Ao��>Eo �x��s��8)��Ȑ�^M��n/F�0�n�|��l-z#�e~�_�V�GRڏeb�N}K�i�+�ÜH��  ���Y���f��2$֪��ڞE)������j����f�E�nYs��I��R�1��z�_���T�����3�b����@�u���L��R����3�*`��Z��~Z��^��k-~cKt_b�]�c�F��̶��r7K�Q��V�pk329�B�2��8l$ٜ��!�E��;���0>C��٠\I?�����§S���ы���!��i���Xz"���h2�Gp�a�j��%q��tq&0�GV	󫙦`{{1���)���RHw��&m`U�6�c�Va�?uHO.�].� 1���c����W~SA�:�Y'�G�+��PS�!y��wA�BO��(P(S�.�������.;"X�C�U<�`1���H���ɶ`7�U�̘'>��ѥ1�
[����
z��]�ĩ8�,h�$T:4u]dX?9Mh4�Tb�~�_��J/D>23flAw�ģ*��t��SOY��.♂p�
�ÕD��lj;Íx�VNz�g"f���h�ʥ[*��s��S>����1�3Ł�I���~�`A��[A�+�R=E��Iz4XR�����w|�
T�q�Q7GMih�c@O���`r��U�O�"Xc�IZ����z���5�s{��ih)%�����+3��<U�kM�E	�+�Zr;�����u39�~�~V�>^�51,g���Nd/V�m���^]����M�����6d�=���.��/�	ˀk��M�\��&90��Ճ<�_=��>��vqI_!f=<)�n�W�w�nv�hpB�,4�ym���Y��2
Q��Y{Gi?��X�5���h�g�JX Z���UirhU�-L�'v����3M�a��)c�;�B.�n`��lQ=t_�B1Jt廋jQ��|~EC�^�ەç��G���־�;�4�oR�32[�O#@��#`�JsK�`X�,�#���}��s���8�y�����˼kj#�fL�	�Ͳ����T&Wx�?M��jvz=����@=�(������P����r�.yaQ�T�;Q<ji����B2FD�.���^C�NO"��m��-�8hCat�3��w?F�.�-���΄?��9�xjgUI	�]#�ܩ���I�j��r#Ⱥ@�ŉZ��?\AS´����X\�q�N��#i���Z{�6��A}ȢJ�Z���)��m��1b

=��c��h�f�gD�Ҥsg�%RKLh�^m1׃c��;��!��Ô�ZҼ���L:�1Irţ��K�7��z�w*��W�!�?��Nc��.�dvg=���3`��Ǜ0#<h[�g�������;�'��o���9�D�Qa��y�+,�����c��'���@��T���Gg��������޸1n����%�������6��_ν2IS+Ma�$D:|@s��4�R�R�������L���fzx
֝���M���8��/	*:5{\�p����$��.�(Mn�Z��@�R��b�������B8�+�lʠw'���L�c�V����tG���_h3i"�!��φ%�Po���6�&�>)�ms��u;0�pē�QE��[�S��a"j���DF�ɘ�
�E�z&O?�+�#��΍�+�GԜݩ����p�����\�������%�5.mÑ[k";�&��:0�W��P9���n�e_F]�4�$׶]�	_e8Y�_��� 6���m��^ÇR�a0�ک����ir 2�����ə|%<�i /n&���*{�hxĀ
<	ؾ�6i �]#��[A�Z���b�B��K���@�,��D�z��Cr"�a\�t-��i7 6�&0�[\�uj��i�����7���-�D�/��F��n�+�gw�Yz=}Z�M�I�9�4-"أ�Ux]���?>�V��v��F�	VK4
R��D���!����vBF��7�/��C��k��������o�ϒ�<-ni� !��T-��F�Ҽ;1��خ�2���i�e�f-��V�-Z��l�V��@�o��c6�|R�q�P��q-�� �P
�W��e ���,��p|�/�����g�2}�n)6D�v��Ő����/	��ԸU<ȍ�y��4