��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�.�&ʺr����$l}��V�W��]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUPc�k�u�}�|Ѽ�r�ν��e��eG�I�?g�f�SL�<.w[!�� Q鹯e)�Op$���j$��N�w	*D���y&�f��+K��[y��ڂ�1aY���~j5���N^�/lt�3� P�;��1�-���f񻲗��~o��:���F�q�\�>Mg3iǭ�lbڎ�Qַd?�X������t�켻�S���c,��# � �bRw�����IL�+�{Dr[��I�.j�r[��f%%e��gg�AՓ�'������L#u�#�5˗�B���	���
��M!�nz��m��+F��8�ĭ��{0��d#�t�  ",�N<��;���u��w)�SU��T�d�\Y>;�>9t���$��Cؓ����9����E�@�ͺ��t�����<(�e�aO*NQ�iF J�Tފ�WItL�5�5.h9�Q���:f��%m�!=�y����h�}�BK9�H��K�|�Ű<=K��:���U�)�c�0u��
;+�$@�9FYg�]�ڽ��_�-G�1��o���sp%II�~�>")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}|
\T s�=&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[nS5H�j.F�6�Z��'i��6�g�m��+Y#_WӇ�s8[ZΑ� �}E+�vl3�������7���	���q���Z&��i1�F�\��ۧ孡4������rYd�ea�;y� a8�����@���rah7Ӿ�?w��K�L�&(�DV$g^��O�>�详 �@��&}�����7��"ꤱ�Ȱ^W�%-C��og$iVdW�E�}�?c�oZ�x��N��2e���m`����[��}L��,��.� U�Ol�#a���j^�O���W�]_��.�O*��i���*.�@gW�%-C��o�.��2�i�Ƿ����5+���J]��$~��U�J�쀴'�뽣e΋*���-������uS�(!(�_��U`c�P�4��o����C�H�
��������+ކBD�B,�dnE��k~x������Wqz^�	�����rYu��1u����@_���P^Z�V��'�e����ʺ�;[��\�v�W����ĮfA��x�%�ܐ�ʟ�]�AZ��:I�"_��V����p{���,�#������s�0F�2�^���=���8��/��m�����W���9�GW���!��������F�┠�Gj���X��XM��d:p{�imlK:�� +@���0X�K�9D���o�j�0�J�vt�OF��������g2Uo�H�0�{�?Nt�!�ei�P�?��'&�s��Ia�|���+,�)��R�ᑧv0-�(4��AYp/ܷ�Kj�.�J�����;*OZ3$�" ���;%x�6��y�g<.���3Q[����c8?-+eN7��c��;��\�v��x����
L(\Ӧ��!�x�!v��v�4�oK���-��%M�rs�i��UQA$��5�%]���a(􆿳����^���2jɸ�����5	���]���c�A�L'�������W��_�ړ8���/��f�VHF��Q�#<4^���|g�Y�'���Xw�E�i�m}6	��	Mk�r��|g�Y�'���Xw��������lԇ�-{���|g�Y�'���Xw�4��}�<�D�o�&�����
L'���Xw�j�7����'�e����>�֔�u8��,�-����#u���arG�n�����KY�ʃ���"����>P�2-i_���F�� �yz��$6��1Wb;T̐����&��4����U�̺��{�U����׈�Ψ��F=e��i��nš|I�&yy�KT�őż�K3����µ?,���t�`�S�S���aB��$�9_��C����A�HvY3���G������߼
�d�,v�M�����ݫ�Q�����6��-�=q�:�x�@u���h���D��uqIUe�JHn��z�c�����<�W�C%����_Wr��;���EWrb������L�j_ R�ϱg#���]b�"x��b9����@<�{1�bYu�c6L���@������LI�.��4uB����x`��:�	1�Y�R�6 q��`_�˜` uqIUe�{H�3)-.�c�&��h�X~��6�='����R��4uB���='fL��ˊ���� �(�V�ܼ��Y�"x�	t�y�9�3����6���@�5��V;T_8`+*��A��}Å�S��P�>����|K�{ߝ��|b0�$3<�H_k.'C���Y�V������p�0ty�P���Պ�`^��3�J��\�v�w�?�b�>޼�\�vų�N�Y�e��D�#�[�����Q����s��'n�^0o,���D�6}�8&x��ߜ��}����J���ɶ�j����+�5[\],�E�ߥq���L�5�e�C�;�[�?��;
V�;���EWr��U�L��Z��\�vř��Q(����j=��T�\ ��)�mZ5#�Y��x�&�F�]:��='����R��`�Z����_�,����0���t���{H�3)-��l���Z\9Ecv���+�&i������Vw�\~^5�C�2Z�<����z�+��p*���Ŕ!P�E����$Y�@��.�c�&��h�X~��6�='����R�J�1���۪	�}a�����.ĳy�"�V��q&=�a�7j���;��D2
�]��x�}Å�S�c��`a��
�?�6j۴�i������D��ܒ:m:C81[��V����X�ޑa������%4�{"�p��of��[�4�u_��+L/w�b2:6�B������B~M~���^y�@5�
pr�����Ac-�Ƨ[���f���_�>c��E�6|�%�(E������D�N���; ,@�� �2�^�~�6����k�G�K�}�k��>\�Gu�����M����e��f�r�X��A-��t��M�+4n���Ek��^���-o��`���;��@�%�e�8��0�uu+��Fz��k���.�)�Hi���i�-�[W]Z�>� -�u�tI��'�{�"��}g�����zL͊�q��io2�&H��ݫ�Q�����6���'�e���ъ����K(�
�cc�V��.�8�T no#��٠R�^Ƒ�Ӣg�w�ԙF��M�����%��/q|M��lU �Ac�N�A�6~��:����{/���kS�h}�L00:�g��U-�e�/CَA�2
�]��x�}Å�S��_��Hv�j×�C�c8?-+eN7���� u�Ů���zPt� ���2(t��4l��'n�^0o,���D�6}�8&x��ߜ��}�/p���xCa��v.kr��(��1ra�"Ɖ�E��T�
�rW��]<���,Y#A�b9����'0Ѵ��V����aU���!�f���ł�!r����|D�$3<�H_D�3U�C�W& s����J'�!�[�#'���ƪ.Rs;���[!W�T^���c_����+#��.X���*"v%)��é�G���cY�~�s<��MR�������c�A�L'�Q��
���lC��U�T�\ ��<��3�
�K�N���IQנF�����F����>п�p=	�˳͠m�xW�J�H�[��'n�^0o�<:�W�_ĵn(���˧�0z�cUL�ݵj�<oU��֜��3�T�\ ��<��3�
�K��¡Ȇ%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7���c8?-+eN��`�6#�6�_��f���K�Q�+�4�i iJa��������ܖA���ol��t�c~C�|��m=�L|Dt �PW��a��K�TR"K�g��U-�e(��w��x�ȳ�5�(�T�\ ���|.�Tӏ7U We��1�pxU����FR���'S/�_wπ>@ �R��P�9J\�e
`�q���ʭ�O7}�»����Ck�MN�3�Q�D��̣����F�z�C���#�^�&F��C�s��e�������hM��1o�l�P��~l|����N���IQנF���ϸ�U��?���D|	�õ��Mn�;��c���XyR�b!����`y���pzl��a겟��`5��}-�п� W��$0���>����:NP�=��N���%Ɩh�����<���,Y#A�_�=�����w�_�2��K�TR"K�g��U-�e5��e6²Cz���\��؀ǏU�e��FR���'S/�_wπ>���9J\�e
`�}R�򳄸�U��?��]�W�m��õ��Mn�;��c���X�`�K-��`y���pzl��a�8���SY�N iJa��������ܖAA/���G�c~C�|��m=�L|Dt����U�#y �Ac�N�A���1#%�"MN�3��cSS�b�(Q6D����z�C�����DP֞ �&��b���O��+�7阒|�6�"�� �J��-��U���T�\ ���|.�TӏpR��������*(�X)󿥠&���Z02{�"��}�u4��d�bR�wX����K�Q+�uB;yUid�4.`�]`�?���� ����C �Q��Y����Qs����j�����{����E����FZ鎬�������(������aU˙����W��T�\ ���|.�Tӏ�`z�_���'���yc����+�J��Y�{'%s=ͱu��� �Ac�N�An��톕����`y���pzl��a�8ݚ���ZMf���9���q���U�ԡ/�f�<�5��G��%�;�$�v�?��w�6l&W݃��S;��c���X����J`%�?�d���&��p��%u֐�U��)���Pa�L����N����w�b�i�j� ���Abs��2[�a��o��� �jf�+��@ Tߌ�\�����aU˙����Wѫ���Uh1�b_X�XV�b�z'hۉ)��R���*qA����6\�4�@�� �-j�1m�I�
Z{�Ck_���'����Ut�\��8�|P�nk�Bzo���h}�L00:C?�Q䨈硙�t�\ڱA�e!�.ؑ�A䧔�Wá.��a(􆿳�^~>��m���F��O��N��b]�f.*A��)�߸��S�Ȍ;`�y�&�c�����M�~�-\��5#Z�he�C�HC��w�;�uh����Wfza�y`+]�3{<�Yo.���y�B?̬N���Z��D��LnP�}R��s��9�;��%YMYo.���y�B?̬N���Z��7��"�,k韸�b�T���Ӫ!�xkx U�_@�N�C��� iJa��������ܖAA/���G���K�)�rW��]<���,Y#A)�/����Cҷ��e�WaU����.oױ9$[{^\�4h�f��꺄��m��'A>�g��U-�eP������e!�
ܯ�Z��pAS��4V`�{CE���'!msR�����נp�Qe�L��}w"�5O7}�»l2�_�V��T�\ �ͭ��t��P�u�.�p��m�۶-�Ez�?���e���l��c8?-+eN��`�6#'�c��=�t*V�M��nDŻ�&ǥ��?�d���&�fTpgZ���jp�6G�k.9Z����t�h��E�&�y+D��䑝nj}�C���&��vt������m`%e�I��m��'A>��"X��[�-�Vb� �D��䑝nj}�C���&��vt�*��]�3ྯ�;ܙ�c8?-+eN�CyW�f�tR�wX��*���?�HKM�1��n��FR���'S/�_wπ>jzT�;D���,e"75�E��W��_�ړ8���/���y��BQ@M�1��n��FR���'S/�_wπ> ��XҴO�6 5��;�¬pX��g��U-�e�2Ex�#V��	��y�`�V���%p�*Ȏ;��|B>6s�i_E���m����e?�d���&��
��Z���7���ɜ��6h���v�䩲$���5�R�̺l��vC�|1,'����0�zG��"Όd)����Q6>"��iMUI�![V��M*;��c���X���%���@��V��� Ac�dXQ6���j�M'�4��r?j����K�TR"K{H�3)-�N�C��� iJa��������ܖA���ol��t;N�09h\dN�<@Iv��nt=:�Z �I�ӦC�s��e�������hM��1o�l�P�u�)�'�m�b�vA`vK7͍��|��W&":#k�˟ܒ�P��f������̀mfF�5.]���^�����p�@��F�KD�Vr[/}>5��0jJ�_/�+�d=i��_��8��GMX��WG ��5��{�3�H��<�C=��~���cO7}�»ԯ�J'>cI��@%B��qĖ7v��\���D��P�)���i���,��V�.o)D��䑝nj}�C���&��vt�*��]�3�@Dx?I�+�4�i iJa��������ܖAA/���G�*5o]E��~�1�|27�Y\�� =N;]%z���5��Z"!�%2��N�� ���E���*5���@*`Dg�8�Hk��|��m�d�6���:Vg��Iقgt��ufb��K���L����6�<Z)��o�B���/X*F��c�D&����\��H��$�)�vx��h�����i�N���8c� \����&��a�C�e��7~���*Y0ht������4nh�����nt��Q\���.@�w��o��un��G�\P��ZY��D���J��8���/���#|�d��5�e��	�)�.�i1��Olkg�^�:����U��֜��3�T�\ �ͧ�����.
Lq�5�p��dߓ����7/��{U��c١�#pl;��K���y�\��F����F3��#�m��}�x��U��";��YCV�Fz�:I~L�U4��\��P�f�e�B��؈a������l���Z\��C �R�x�kyhw�U�1�he�C�Hc�|��g;�X��WG ���i1n�6P��4,�Q����W��'�)�Բcf�x�HZ�, ���q3HL�1p/-��}-���NHRxF� lƔ��M�c��M'�b�	�)�.�ij0���!{�"��}n�m!t%qa(􆿳��ύ�>� ']v1�_ُ�&��b���/Q����ߝ��v�Y/�ܜ�������#oM.�����a�x���Jq�Y���y-T�OB �4�r6�h}�L00:� ^M'��k/��m#'�a[μ3z<�_�_֛��pP�i�a�sirs�"��=l&�c%=�)�a�x���2�b=��������W�6?���Ө��'�hiC���i����  w��_z�X
3kZ��<GHj-�_i9���xQ�m�۶<��%��������O%W��ł�!r��Qטg�u2��R�xbzbM ?Z����rW��]��C ����X8��8���/����$������aٔ^?w9Z� 0��}w"�5 �Ac�N�AO%^�p�c�g��U-�e��pʆ�)�x�.���:��KY׏�����M� �U�O��/tD7Ijl��6J����!���c�A�L'����eq��".S�i~����'9tT/K��_�&���j-���aB�����rn�����P�7� ��.�[ ٓ��r_��m��"(��l�)й�e�Ɵ�s���%�z�J��Ϻ"t�Z;��6J��(���27:����aٔ^?�����zyN5���P�L�1p/-��}-���NHRxF� lƔ��M�c��M'�b�	�)�.�i91����E]v1�_ُ�&��b����ɮ��؝�b�Bϱ���Jq�Y�����q��k��\�v�07�����B�R���>_d���T��jsrCm�k(%�ar�s8��b�Bϱ���2�b=�������AԢ�a\�	PcM�9S����q��k��\�vŅ��J���_M�<TC�}�����:(���27:����aٔ^?���w:&��ˮ�t�s�'�)�Բc*�r#�ӑ���?O�y	�)�x�.���:��KY׏�����M'Ƶ�s]0{ɽ��&k@C�Ɨ0z�cUL��.�^�,��K�$�z�X
3kZ�ڱA�e!�.��t�>/�u��,P���_Wōd>A�T�g�v��o
���^��5ߧE4��
��T���x�;	㯰�$�)�vx)�K���'�#�c����ҷ�R�Ճ������-��U���u霴ԭg���NBq�`c�!1 ��Ktf*�gLYR!�rE�j��8�b���=+��<��](�!���`���\{ف(�7���n��T����C ����P����=�WK=Z�R�ڠa�r�"�R㬽�mV2i��h}�L00:�^Y�`��O7}�»Z}�R+�!�'��أͽgF"?LO��M|�sPn&��|�"���>� ����G�e� U_9^���\�}����� ��$A"u��p$(���%����H���=磡��{��1Y�[�2(���($�|�*��=| �����a��Y� ��|����:�����A�A�C��-eh�/�Lg�4����&D�)>B:�Z�m�۶t�����D�P�E6�n)Pf�� '���Xw�j�7��֏j��[���_��*`Dg�8�Hk��|�օ��x�����M���ߝ��vԩ �E�p��"X��[˹�H٫!qĝ�&���w9Z� 0��}w"�5O7}�»p�[k����Cҷ��e̷_��yC��S8�k��m�ݧ�/\t}-�п� W��$0���>�����qD�{��/���k��Q�D������X8��8���/��NjX�U�6j�"Hs�󌘓S/�3�	����;;��M2��<LC9s��� �*$��x�9��_ڟr��GP���*�N�^���\�}����� ��$A"u��p$(���%����H���=磡��{��1Y�[�2(���($�|�*��=| �����a��Y� ��|����:�����r����TH�&��b���/Q����ߝ��vԩ �E�p�g��U-�e"�A��"�Y�{'%s�.W�jb��w�I����''�|7�=N;]%z���5��Z"!�%2��N���}�Xv�9$[{^6�nX�7>�a(􆿳��@�A����������j�>���/���k��Q�D���R�%ǝ�rN��t"O]��!���c�A�L' 	���ȹ� �tw iJa��������ܖA���ol��t���K�)�rW��]<���,Y#A� ^M'��k/��m#�ݾ-/�;��|Bφ�=�cc���)�p�#O":S�����X��)Am.#qf��2Lp�����cSS�b�ь'��5�6<���,Y#A�}}���*�/�J�0&[z�k<�%'tF��;�I3Ǟ|Qz��������Dm-�="D�f�ͨ�1Y��e�\�*@��ا�D��Z?����=d-B���K�TR"K^�kO`,�cSS�b垊*���-U���� ��h���1;��|B;���<A� �Ac�N�As����,��Q�D�䀟ju��Sk4����&D�E���s��U��֜��3�T�\ �͊�51�X�c�rs�i��]S���D[�l��a[�S���h��P$ iJa��������ܖA���ol��t����aUF�7'HR9q�}w"�5O7}�»l�2vh�1�{�Y��a(􆿳��˜T�Ԕ�m��'A>g4�����������j�>���c8?-+eN��`�6#�-�Vb� �Z鎬�������(��� ?�8���n�F���5�mb��k�OM�1��n��FR���'S/�_wπ>;>��^J�:U=[[���!�=�ߝ��v�R�OE�#��Q�D�䀈b��r�
M��ٌ�AmY�f�k
�K0h��A�J�XY�5��uXC+�>��mW'�J�5u�����(y|1��UU�w1ϯ�|��^��S��+�����hf�Ҋ!J��4���Lȕ��'�B�#�
�2�l�w��#�gŻ�&ǥ��?�d���&�,!r�*�}cc���)�p�#O"
�D�V�` ф�A�xX���b�.�V�F���A^#����6c�+�����RИ�ա���ߖ^�wp���u�����
�r-����\~��$	D���l�^��� n��R)��'/�bD�<%��}�'<LC9s��Fs��u8�RX7���#g�k��qĝ�&������w:&�����*��|>����n�T�K�^d��]�!��	Ǹ�y85���]��^������.'�L����^��''�|7�=N;]%z���5��Z"�'��G�<���,Y#A	u�e�2�?�m�۶�so����O7}�»�QNȮ���k/��m#�J'�!���=�@qI�A�5��黦��레%4�G�1�/��D���J��8���/�&k@C�Ɨ0z�cUL?��[[��,'�*;kO��u��"�C�˂j}�C���&��vt�*��]�3���p+���b"u2��O�/���k��Q�D�䀭�ĭ��Xw��l(�i�g��U-�e@�0Iݥ�Mj�(ȅ��Z������ܓ���'Ս��"���<'X�|��I~�v�(�>�{��D�h\�J���/�hD({ՒD�jט~���@�5�^R�[ZD���Sd�o�#���Ik�m�Q�<��W�2�ý����,�ǰL�[��V�����J�u;��|BI��r�{׳-�b���2��Ȅ&N+e���ٿLv�$�`K�'$vr�����&�j�^*zV�}zj>gm�$�kT
���ۚʦ�9b	J?QW����h}�L00:;��|B����ɺ��K�A�'�rW��]��C I7z^�e��A�T�g�v��5S��f�`�80>,?��Jh��� �~�9rF�؀ǏU�e��FR���'S/�_wπ>��֩mh}�L00:��YJ�;�rW��]��C ����X8��8���/�۪	�}a?�d���&��E��(�D���G�/R{-z�}h}�L00:;��|B����ɺ��K�A�'�rW��]��C I7z^�e��A�T�g�v��5S��f�`�80>,?��Jh��� �~�9rF�؀ǏU�e��FR���'S/�_wπ>;>��^Jh}�L00:��YJ�;�rW��]��C ����X8��8���/�۪	�}a?�d���&�u�܃s.N��!Όg&W�w��fD��SfC"�1��n�G[������o��_�,���� �Ac�N�A Ҳ́p��y��K�ݽKJ���� 
~�F���r?j��h}�L00:;��|Bj��!(�#���^xJ�$K��A^���\�}/��/��ڳU>�f&��'!msR�����נp�Qe�L��}w"�5 �Ac�N�A�a�sL�g��U-�e;d9ךp��4,�Q����}�Xv�9$[{^G�\1�����"X��[�`�L�iցc�����M�~��������9��L�%��x�-
�΁#g�k����ξ�|��U>�f&��'!msR�����נp�Qe�L�����*����6��	���Cҷ��e�|��*��U>�f&��'!msR�����׽��9\�	Z���/:���lC��U�T�\ �ͭNjX�U�6j�"Hs�x�ʤ�^m1�H���W�w��fDP������@[�_zβrQ�ͼ����b�A`�Ҭ����5A���t�T��S�,9!:-I/B޾Pk���e��q�w~��A(�c���_G��Hb�ñ ��3�JJݾ�'�\{ف(�7��<�h�#���C �AƖX�y���?~f|��d�����w�⽒�;��c���XL;jy"k�{H�3)-)��m���� iJa��������ܖA���ol��t;N�09h\dN�<@Iv��nt=:ྵp�!����&^��b5�sw��
�(�V�ܼ�.�%Υb3S6 -�&���^a�nu4Bޗ��jw�	��-��@�%rk�,l����M?��y�NM���������[V��M*;��c���X�8vw��^C\E�'����f	������"O����n��T����C ���Ǭ����RO�?��~]l�*`Dg�8�Hk��|��!�x�����_|���N�[��|������hM��1o�l�P��~R��b��N*�95��{b��vW'��}�D�Tu�^?�&^��9�׍�����u���?�)����^�{"}W;��ܐ�}�۪�G���_��e0�@\}p