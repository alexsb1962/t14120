��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����Q�c_�}h_�"�A�[f�.�%a���f���zxETQ��o7��������r�m�@�'�Q��l�+v"گ��E,�29[t_y�{��)��a;ʮ��yt�JO<7��c��Ʃ/�;���l������2�1��b�<}��n�^�L@���P�Q��P5l���=
T�n�y��2�Wz�Ԟ��fa������ފ��m���(J�)�g�ڷ02Dy���3�����oC�AE�ey��v5վ
�+*B��k}z�ڏ7�7��H���ɣa]�EV�<œH�m}�"R�0�*�آ'�]R����>����+B��Vt������kd��>)�Qo���:c�85���s�+���� �~Z�=�2�5�k�Q���1�?Dk�@�����O�i+LQC�i/V7��O��d�����R3�gFB�~�)~�Fh���)^�V�F��"���
�Я�3�򰦫v��^�*pЗ��h�_��o�M�a����Pȣ�^H@������S-R0�D5�)-��1L��ֲT�%��Ƽ��w�k���̲G3}�~��>?w
muw�>�������]w/J[e
��>��]����G�ZZ˙x�:����ה�7���f����ؔJx�`��Ş�P��pU��\���f�ۈ�%��tݚk�iО�u�A�[@M�^��X\xv#[��r���u�9os�t�)3�O�BQ�mכ���a"���Pƍ
�2g3[0��9���������Ͷ�$~-����8y��v�1!ޫ�|zBq��|���2�n�R���@ꃭ��c�c;V�=�R��t��=��%��C��YO����1݀�R"�J�7)�Ġ�'�`.;��Ox�dM��]pk���A�.'�c��ZIg��y���Q��0��S�_ ��Dh8�p�)�h���i?�/~:M��?�vA��x��RDq:r�N:~(�e���z�C�X�/���_]�.�;ބ5ώ���?�
99F�ڤ9��𘒍�jmx<Ó֔��D�j"����xu��C8X} S��Ϣ3��"zue��Y'�:�t}����ѹ�ܽ�81�ve���p�b\)���L��@�-�Q̏���R�ڈ���U;@�2
|�HD��1�ɟnp �7'{|O5�O�;�~�jބS|R��N�ʕ���,��V����M�~�6�ק�V��ɷ!U�[����G���b����F���Q��ȱ�ln�=�|��n׎{q��0��h��Z�@ �En���*{���G/_���3`x��`.=5i���i`e�VS:4#���F���&��q�F�aL� \�&hU�r�}���Q"��P�HK\��%Q@� K����8q��5����{�������_�t1���?~�D�����֙x������G�����u�F���Xw9�ǧ�Ƕ�|fJ�XQ����(�W!��*�����&�����da��7&�7z�X���`�g�,�K..CL����h�M�c�
��