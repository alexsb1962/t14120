��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aЫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α��wԊ�6�a�3� G��λ�:~7 !�v sh��~��P�'|#��x�C�[�~���{-چ��!�:���)�#aE�C�;� ���&�'��c�w|�:�)��$��Sއ�Y�K��N�4uFLN��6n���)G�Kh\��V��Bm��ĠJ�k��!�Ll�!R��Ѕ"���8Z�ɼ�	B��o���Z5T�Y#m���og�x]���S߮_�g�@8O٘00�.�wJL����]��A�Ej�N7�:d��zE��~}������I5��;��0:W�'�)T�WAP�LV`���Z�)��Vu3z�	`.Rz�lLtmśKN��6�i�ǯ#H/u�Gl���3׋]�	��J�9��Z]+�����3��t���\V]�#��ܙ�}�9M?���Z����᝸ž�U��d�:�H�/髝�c��2�e�_��%Y(m�E���b�cU�KA�@RgސY�/lͫ-��?��ޅ�UE:}�M ��{�VL��B�_:�S�(J��<XR;��]Ƅ݊���K���hp�T���'�O�f{u����e�"�7�i�Li
[��)�z���?F�`�R`i9?,��%� ��e�|�>c�׏�"/'7�,�i�Wx����`#��	���K��Y�#oMIW�V�j�xtkE��8�j!�O���"��\m�Y9�i
�/V�
z��H/4�\��J��f6��iFL�'�_��*�3x�H�T
�`-��'=�Q�#\q~�E�U+�6L�����a�ox�`�_�HҜ�
�uC��>�_W��]�bY8=�Pw��W<�AC4�7jJ���f���X�8���
�ի$~A���n����a����o҈��v��ٹLC3�y�X`Y��L�KzP��r���22�l��ۏ��80����kNy�.�K{i:m��k	���rm�v�d ��0@`֦����*���F�u��������Ķ��]}b���z�f������2l頣���|�AUehJli��A�n���L�~
�+����U;F/닅W!�sk�_�L�1��*������V/��uGk�`�	��0ʜ]�j��)�꯮���k����l6�\���,�_��Z��.E)�fo=��p}򍷃�7S�?��mrE)�} �r��@� L�n%Hv&��s�!��o������D���-�EEc���9&�QS�G�f�y�o��y�����Z�ѭ���������9���@���IjY?k�iR	R,�͜��&�VOwl����ae)@&��f�˞	�����c��5%��cA-!Ev�M��xـȹ��Uu�Bq��E�K���6�y��
1цVç���K��Ϲ����	\%�dj�p�ޣ�]9�jݣ�y��1��Κ��y�����ױ=��M'BD��X/"�Ztnu�P�\�������uKΦ��0��Y�NM��2�2�����_�&3K�
��Dg_v�7�b��n���6��ȭ��&.ӭ�"��_�.����ɵ��{#YB:���w�=wƱ���F�L'�K*W���r{�H�/2jV_�b���c5�A��ֽ��`;o�.�K� c�V-�B��=Fr @Hn�n�@}z��DM�������%��8�6����IB��,�8�X�)�N"�6�W�3��Q���+~���sqx@����Ie���q ��+�@�%υ��T'��Lp����������P�+����c��?eۆ��P4�t�q��%��0R�:f\H�D ��o��Wg����oG�A9�b��A�6�y�3���t��<r�l�o��S%[�!����\�K���3��J��j5����D��%Od;�����?����m��aگ���@I��.��/ᒵf���n՟�c#��_T�q��}Ey��D��	�^�~�4�2��5��M���vT� z�Ȏܿ^ _K�����+���Vr-�)�Zbh���o@Ž����yeMb����:�G�ӃŖq:	P�WM�x��8a�̈́+Uц�8�h��\��y1"n]7W�$f5,��v�FTX��7����LW$�`��SqK�X�%5ѣKB��_�[ ���z5�wy�Йw��5v�)�W{Y�K<�3
����3�TE�7�ŭ��x`6\�֊���.��	�?WP�<����phdI}�i2�'^�蕑w>us������R4K��\�2ٺ)�_���(�_l+�2�`m�AR�/�Y�F�)#���e1���	��:��S�*M��^�T��6�a����_s--ވ���S�;�l#O�.�p�N��V�XO4����	�%I�h�"�C��FW�+��Zw����ܝ��4��R������C�}��"z�y S�;�����"�c�} �d؎/W~���!L�bFn��*�����[aZ�x0�8����ao=�f5�j�-t�rY�-�6�](
J�Ȁ��x�Q���򣎡l�j��{e�0��8�;�����?����҇D���rlg�W*Ln)��� ?����)~FoG��L)<�;$LE�D�>*v=�2ч��[{��zmCƩ[���Qֆ{��ؿ�������Tu�<��#r%F������$�v� c�|��f��%�޴��l0��!��^�����p4�4�#%��YE�c$����$ƃ!X��~wv�8y�V�a�� �97��Y�j�������Ҥmm4��C�v�K����uK�>�v�/s����3�e�KqKC~�aC�A�a�6kY��i3��k�m�}�=���W�'��V�k;�ڃ-��Ɉ��o�'�r{�-��*�I�@G��O)�|~��W*S�Ɖ~��ⲛ-&� 
öX�����Ϙ҈��Q[����za��G\k�^�-�H�9Ų��ջW������,�%ք��ߖb�k��ڌ�06^�F��]*��n۷A���_��Bz�=��]3��l6�Kvp^�ث��;��>MqЉA j<��۟��7�ը�ē i�M��$E�v��?� ui�Du���%ϒ��������I��@�R����!����b3�a{����eB�j��D߱/t��7zsv^C�;A<#�<�\���.f���