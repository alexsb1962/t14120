��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������LX��a��?;%l=UX�ƲZs���4�
P�û����v�ܩEut����S+��������S�Žtb͕�!�`��!�ۂ5�VF���\�gC���T�/s�|�Mu\�s #�˺V�HI��(�.%��$I�a����ь�G�V��&Ҙqs�?���]!׉������Zdβ0m+��K[�,>���	��n1����쫗JWI�]�84�9�u���q�'�H�.HC��A��|L!��d����ˈ ��\��t�͕���ei��
(�~I�2�}�)�"�f�,p��Ǜ���e"�¦,�uϤvEpX*Yv��G^� ,���?0�0��[ԍZ��f�߃ց�Q�3���2
�љ�'��}��`ҁ?�pP`��i�f���Խ�&����}��Ln@�Wi6ފ˻F\U�/�n�WK򣺜���x��Sm�0'a:t�:�S�B3��G�����W����͌��"�$�7Nh���.��˼���@�u3Ead���"M��o�fq;˛=��-�uB^�4�5ɴ�YK�/�!�f(㥗]P���|0��&���'�Vwg�ˣ5zm=K"�h�\�����K���&»����cG����	(�͕O�J�l[���#�&�@*��\�mV�
�e�Gː�@wۡ軷��{�ߡ�`�3���I�St�?���I��� %���{H������6�O�
~��3�8�����������w ��ۙ�-pC1w͇���冷P����am���ҞK�}���Khڷ� G0!N0I�P�8��qO脃p��jM�e[����iɶXE[��4���ӥ�Q��3N*�xX�FݻVͲ�oڐow��T�>��M�4�i�@�6ړ�ȗ����~[�`�����_�����͎��v4 ��>�[�=�h=x8e��f���(�9���}\p� ���65CW|WO��}R���d���������G�( �3��p�E�d7�)�Mb�oO}����ΰ�H	L�D��?���}k|z��T�(g���諭�t��_+�|���m��5-_�q�a�X@�UE�6ͻ"3��])��#BHIk�-ӒM)��I__� �Σn�pa�^րUs��~G�}�[7�Jd�1�U�� �[+�U�rś��Z��);e���db����r�zB��X�n�´E��M�	�QoL�'���M�B�[hnV��\����������rSFX-8�-�����z�:*�}�?Ed�Jc��Q�i٩��O�j*W[�r�L�c����M>7w�S��u��5�yR�.i��Z�o��I�Bj;�