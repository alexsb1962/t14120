��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������,��r�'��l����O�$���i��;�[�^pr�*1ժ���K��FD\���7������׺9/���� �1�nT2gvf؏�=�?����&��. ��Ox�!���W�uF�����q�:���or:g��؈ѫ����ܹ҃��`jY0��m��fd,
A���Ǫ ���l���M�Y%�+�]tkZ_xz�*�]K�I�{��Ǻ9��#�֊���X�^깘)��i�������4�-��d8��jo13C��\p��Ԫ�-A�D�����D�޲5���bG��Ƙ�Ɯa�z�pc�r�f=��@�Y���,
y\S�1C���ϛ�x>�N�ٽ����>+���su$��m��n4\#
�k5ԺԎ�b�.r�NM�6z���)�CN�gm�]Fx@�;��M-�L�:�RIA�$f�0��>����u���}*sJ
����ȵV���N�m" �v�
��q�?Q�V�<G�%�o�������ؼ����@&;�(���\����5��z�Z	D�&c��4�~3	�,|�l�#�F8�W��o���ͭMdR��vBR�)ig�U?{��6{����]���lm`$�:�$����D�?C�T��`�X]5aLƇt�p�F���IWodB��|Qz۰���U����*e�0�x��X�y�b�⺞�yCzbv�t��DKAz֚`�k�����#ǧF۰���w�.p�>�[�59��4lJx]����c��9b#c<���/�g({�h6���5�ɗ_i�";zl���IT�s�����P��h�އYѴն��b���`���H���}���Jp��N~<e61��9��ucP�#���]����w����Y0�3�|�.J6�T7��@cMM�v�Ӆ
#b��z�B������J�L�1����7��yB���B�an7�n��(;�&Yj���n����%�r�
�/Vᤂ�Ve���~��Aȳ��?�:q���|�|�9��fʼ�/���K�>�b�pu�v%y�|oW�c�4�9b]�(Q�W����8a�����3g���5p.�����H4���6�􊓎\}PBa9� �*��lmRoQY/����}��Pk�y���(3ƜFlה�Zn�l�v�)��*���3��Vc�l�eF,>���^���3ِѱ |{�����a�w�U@���Uu8@�z���]QÀ���^l�7��.�r��/��x�|y�|���p��K[Ǚ�/)��*���-ɂ�b����n�=�Ϸ�郈-�ۥAv�bi5�R�I, 52`����zn�ihБaV�_'X�X܁Y=1��PʷX,�8���
����1{�^u��QS�r�.��8�3�Hq�*�oL�AU��M&���k/�ߡaf���^�j��`��Ã�szJ�~l���-k�!c�>'Z�B=�Y;����/U�!<�"ur�\��*d��A&�g����`���Q@���ҏ+
"#�����v�Mf�{"�)x%��ؐS�`����ڛj&�^�iTp��F�Iѫ�SlF�E���̄�5�6tr*�|Rھ"a�'�7�d��A�/���������L�H&�x@� U,�Uڣ9Á��j���w�7�I���8��q�,�L� c�\-ngPf���=d�85O����g��M%I/r6_7��%�	�T��&hϙ�ͼ�F2njZ�(�u��gN����EL1��ߣL�w%�~���4E<J�Z���|�&�F]|��qx�/�e����)>��Zo-}�H��Wyh�XWh.FYu&В�3�6y�-wu��9X�]�rq�J��ybt7ȚU�� rpV zY�h��e7����X�C���e_�_)@�,ɬ��+�Hsy��W��#U�S�%����-�K�>���E�}�.]�w��,o�K7���]O�S�k_�#\��{��$Γ�)7)�v�9a�ֿ���%�@5r�u��-	�ָ� �r��9=�p!��N �/$��^@H����b��
gT:�GN�z7\��׵��84�� C�������d �?��0g�����a�(ē�G�7�L4��c,K��^W���yI��& R"š�v��3��D.v�����a��Tg�WMc�eU��b��I���E�њ���zuh��N�vN�B�#��D�ۢoI�$�g�f
�g����w�b�D��������o^ecZP�?n#���#U��t�60��A�^��`�;l��D~���(Z����I&�@�d*[;>���	8kft�+b����ʖБ�dP�V5X�l'�id���:	-)�Ib�+RʃC/J�n���C[g%ZP�A:�C�����)7gs���g�lb��Qr�����ۦ�?^���WsS}!.�9��<���28��N1�3e���5�q��u��'�/ ��X��k�'���|��Z&L��G;�l7��$�+7��u� �Ϳ�`|Քk�"��Ս9%��*��Ś>���n'?#������J��i�������/�3k����fz2)]��Gק�4���ze�$&�� �w�K��������eN�l��ݧ���?�0����:1��Ȣ���L}Z,���T���n��#J����RH���i.o�
R�����̐Nm[��5*�/[�m��ð7�+���#sV:�����f����/U��m&i�g�J�O�v�ײ{!RJ}��m���x;t]'�2x��h/��Hx���ܤ\6��խ��e�X��l�fJ�b�*���#�t�T����F��Μ5煭/4���z�g˹@�Ǌu!�n�⌃©��5�N��.Qik�h��1���Y���l��Ta���)��K�k�&�4�8v�"����
71c���(:`.���߮�)���3&�'�����z��n)x��~�
� ��s������LUõKB����>q��FZ��>X}�)��_߉�4y���)+bK�b���1�3OFVa�I%������Sb?dV�,��m�ɺOt���$w�`k �h���x7��Y?N�#���O��%�g�2T�ʤ�A4�0��H���m����Q�mݫ>?��o�3_s�D��IZ�k�v>�dk�;ޭ�Ԁ�����7S�[��q]@,�r0�t������\ 3N�F�#�$�䃈�UF�3M��%�^���#�It�3�t��&;�8���1d`m�p��8����n)���������;�*��5��h�Bѽ�?2��FƢ|ݷ[N�=f�ײ?�e��rٯ�1xd�?��)x���d�KO�w��A�,�C�62%��__��/�f��Q'���r���5�δ��M�~��q���WŖ��u\9|�".��	�O��i�.�郇�X:M�bDP���:H	��7�He��~%��oi�e�:3QLN����h��]\��b;��XϙT5Ȝ�>
eUٟkj�:����d�_C�1h�mm�m� A����Ә�1=�J�X_��.��܅d�p� ��V���ͬ��
ϖڴ��.���ly �W+5AM1�\����o		x�`	z?_o��Y�ٳp�'3���.C��÷x�G�Uvp��#�J@��Mݮw��l�G����P�ukl��9���-�Hk�H3�C9���g5���"N���y�><�(����]�D"&��uWO3`$m�'�}���b�>t��=�\c��� ��G�9��0���&��x���L���֑��W���Ir�0��s�'��Gބaz�1�!P�
�^�%ͥE�NG�֜��t�$P�%-3u�v@u��S\�uhX���wcB�g�b��FcK�/�AS�u�Ia�>�KƶR{���;��*�j>�%��^��A	����D�O^�w��B�7�ȋ���Ζ�K��b�zM@`Bq"T�A��j����f^i�8y�>��u���x)ũNѧZ>�z�YD���%�.�ۗ;w��2uDN^�cO�ZD6��}�j,cgOie���oǹ����u���.��'�n�iѩT�	{���
��\�q9���ݼ�M�$�4��Yၢ����{r
�|���{��]!��A:���Rc8�L�=G��Nv(b���_6mj�1�� �+J m�6��`����1q�4c1�)����~�F� R��oP��&)_$�s]w3����딡�,-�o��JM�
!�~��r�n�[2�ьGȲU"S��{��[���> 9/�6u7�9<���9�c�'�O�a)�Sxɔի�S$��������t`f��6L |E��>�t�3p�Pqs:/҃a��Jw+�pS�/﷞���?d��P@�9��
5nbގa���7������.g��1֙��=���v�%�����~F�>Clfg�mV]�1�; �Q	p�����x`��O8���8+�Y�S�c�C�H<ѹ�^�ţ2�v&�Y���P皫�.p��4�|A �wMF�?\�KΪF�7 }<.x��!��+7(=P';I�z|n}*+��n�X�l�,�"��4�Ȳ�̈́���07�1��<V�N��z�*ڤר�ۯL
ׯK��'����J4Ⴅ�f�ʍ!��D�T
� ��/�Kآ�W�M�*��NG�e+ô*�����_���-|�0Lu��n��P.7��L��L��WN���S��~\��[��B@��$�VQu@ �y>�qer��Ն�gs�.� dip����?x�<��޾�$[T�����/�U��Z�ۤ$��Q��j5v�p\ש��Vܜ|0B
UE6�:�|�ڄ�d�PѰ�6;c~q=�MI���6å�uz���Q2��`�7��X�p�Zh�b�dI�?:�7��0/^�#u��XN +w(�Wl��6�fv��ѡ��`���]��z9�p
*ߵ`�a������yU��QƁ�T;;;�2�ʆ`/����g?{{��:�䈳�Zu�N��"�	��X�/	�J��?K������������ú+�?,��s�B?�G��[�b�K[Ex�4��d�g��5�����G|�E�����r�Z�&�p�ړ
!��z�Ύ�2"I ��
�P�Z�7��!{�%���)����6(»1���n�3�ﵪ&1l,�V"��KD���]���A��:=:�z�Ќ#Z����z8���AY�b�1*���I	N������N�m��(�o]� ���H�,��U�ׯ��?%v��d ��������|k��$���yi�&1F����I��
�	iu	�Y�Wr�1��l�P�]O����M�ZP�rժ*�l���UFK(��zį�| }����35 ֩��vѨ�����V���ev?����A��sŋ�k<"3�<	ĳ��帙�j4�b�7��Ќ+|�.�� x�=$��k�b�} �F��l�/S�\���LY
�~k�"�pm�:�SB��-��&8i߀i��_�L���C�R�z�&���$l21ɥU_E��B�(T��^"�S`���3:oK4��bf�`T��f���]>Ly-�ޅ��M�*D;�KO����`�/�`�/t����n��X�g���5�5��g�l����J�#�I���b����vu`<��wӽ���7�/�:�G�-�R�KG��߃�/O��	�)6�#�5�����9�s�߷Qh]�������,�O��E�UVB���Li�����jmsa��G��ܰ�p��xj�%���'S���>�=,>��
s��9ً���ELE��Bv�+�xvJx���C׻9p����A\FqZ�V (J�g�)�d�>'��ԭR��)kY�>'���c�48��m��RYCZM���ys>H˨�Ї����������B���	����k���i�F93�P�
&�J����3!C�'��d��f��o���^b�x��LU���x;k	n�7�#_R~�%\���&��8G�B�$�*3�]}2�A�������K����h��=�\߄<�tѫ�ޒ@�X�+�1�.�9�K+)��SV"��x�����{F����4Գ�S##�-���@�ߎ"6���l�����(������9#3�2te����5�){i��xxUȳ><�Ɖw�lo������O�7�)��Ȥؙŕ�EQc6i�	�A�WD�]�$�>��)p�z'⃸��3H-)˨�Cm���ifVi���7�(�6_�� ��J(+s�Y��ƕ�v�����#svR��d���]uo3��������i]`"��dP�j�����O8�Q���q���kz�?� v,���L�/1���#����߅����8)���S�w���Y8���acϢ�#�ʜ�	�ug�没�XzBM��ef9{��Y0�Ai�+�B����}�CM�Õ�8��k�Ä4b�V\1�H��Wb�p���@�.�E�)�s*�
Y$�ۇ���~��U�������}�]��餔ማ/%�v�_��Hj�}O��,@�^���Xrt����0^�r�o�6	�V'�O~��0�i�4�+y��е�^��{���dk1) u��%�{������Yܜ���1><=eq�#�|���5��w2|�l��"u�� ��o<���T4�C�Xƕ�|0<�]4�������7�̗�z����ű���� ��3$���,B�ZPx�/�~j1�4Ct�1q��:&%-��-A�Οp��wv��ޥ~���� oC_w�Pԥ�1�Ͳ%�T,w�D��7o�K��n99s��k��-� ��J�S�&7���[�DU9���E�9����@�{���E�(]Qu��l_����]�Ǌg��E��O��4E����k@T�;�4/�*����D�$yczf}���<���%MG5�gQ_ۺ�Wπ�JT�%�fX�Aʬ�mi���mƬ��:�KQm�2�:Q�=B���[��W���|�"5[�5���D���r�<� MM� ��,V��'nf��sD��>����;���5� �q�ݜ��؟�b��#9�kotNCƤ��S����9�a� o�0;�)D�=V=p�L3doZ�	I�<�-�g��mkW2��v�CXb]�+l@�D��4q�P��f���S��rm��9�/��S�!u�P�ڰ+g7g�_�ĿCY����u/�}�u����oφ,\�ߨ��Û{�3=�C�{����T!xro�%����� �˻X?�{���C����"�7�{.i#P����:a���q�S�?�3-�h5d����f[X�,c���-*W����"�'*����0KͰ�1u���@�b�X���H�z�ܖz�q�{�<B��o�����Z���!m�毉���+.Q�|����]$�+�&+ԷR���5y�͸�$U�R��ɂ�KHR�|=쨤�W�_�l� إ�lSh�A��VS,�����>���	������OQ5= �v�B�]3�p�W��bO�;��+<����_@9q�~�C�-� -oHO]�}��e����6����}S��M�g� ���]厹�y�,�����OcfB81�`*Qc9Kߐp�v��$�彤�8o���b�z��@w_e���i�QE�� �x1�`_q&�4%����Ö=9
�q����mٜϥu����K�d��g6b[ܻ=kw�k��bb���7�S�b�.�ꌗ���RL��>�v���Vc�� U{AE;�]!O��3��_WD%T���N�M��)�1�`���=��0D��>�k�y�F�?�������n�I��pYw�q�d����ᜟ=Y9���v��*����\�>��>=��G{F7�/MP��P};��u-�J,}�C�X�ti$�ѕTk��=��F�f�:�駔*��0��P"hR݌����!�����*�/XR���̞0���/�#㽁���n�e�Vcߛ��'��u��7"����F-����(d����9�-� �*��lR&��4>0��!�˸��x��U-a�ј�}��3��N\A�3"�&K!�P��0���"��]���{�g{� ۤ������$�t��_ۑ�Y���a�-�[f"\��Y�}��0g�k2DR��#He|���Z�)gW�Ly��+r��]�l�ڜtb�'��!X� ad]���xj�M����7�|��5S�,v��m��iN��gˠ䵒��/�yݩ��{��8ή	�Z�����������2��`�՘��Q9n����K�c�`����,\������v��3uG��m�lpr˸IN���T���@mGE�(��n��Z�(����+�wxƢ����7�| ѻ�q�Eb����ޢ������7&9�L"љj�=�`9�ȉ�@�|P���XK1�Q�a�@K�?��ܪ�]ޒ�U;����N��b��J�⺤�8��N۳�!����{>�fgl5}?P��lރ:��������W�^͋��e�D�%�~f6^d�p���Os�Ls��~ƊBJ�t��=��6)�t@�����e8Q4)�Z���0X%;�����I2a5�&	���J�U��R��!
��Ͻ%[�KᏃ�����i�:]�Ռ�ig�po�z�d/��뉞 ��#|'���(O�������|Z���Lpˈ���SL&����m�i��ޯ�PK�B΂�=T�����NO<��1q@~����H�7KЇ�X�OlĈ��Im2�v �F�r�x�1��"S;�d�B���t�(Oz��r���%�?l��lJ$E'\�������>�:d��i���,���&�ea��� HX0�K,��:5�Kt�⿲�.5Cd�;�	�����/���U?{�LC��Py���| )���jʎ-��$l�����G��JD�I�=�޶@�{T��ۤE8/=8"�J佾tz'����Uz�t�s�����n�5�)��C:L1^�%�0wD;luI�<���e����o�~Aia\=r8Kt��nQ�����`�Oz�'W0f-^�8 �i�]��L֋,mN��>�˨�:Z��M�;m�*&L?&^d�r��Bo
{��/?�Pgn�(��a��Dٗ�  f��Dڛ�� 䇙Dbi?�X]�Jڄh�����vU�)��N{��8���4Zӊ�����^PЪ��ߍ]��֕u��q�._I�id�� �Äp�&���ME�Y��K�gք\D�]c���iB el��b��y���K��#m�k ����pi~�>	��BP����;�28�G٪��Z1\A9����~iŢY�u���'��\zc�3����Οk��9[��T��/'�A�9���t��b�L�:#5c+�Y�}�����\_EK��w4�P�|��b�E�Id�v!$��$`�Sx�9+�ީRf������g�(�c�ar��I�y!<cU�P��3��QHi��em���9�,�ҟA����K�4�3�ӽ�4�f�xH�Gy�6 �!�I�M�;��j*gT��ſ�7�<R�D����������ڕ�U{�k�jd�D#N?)E����ρ`�%;��׀������}U|TM�X,R�#�Í�;Z�sK&.届4�1΀�����F�Q{J ���gm��A���r�$�@��M��@�h'{BLQ��L����6b�����'A�R6)xxA{4]���E(%�;��Z`�e ?~����R�˺�=t*�E�w/a@�!�D��0���h�w��s0Z�IŶ�����ΘżL�A�;x�c��!�ϭG��ֿb�v9{M�`,�]�����D�>`�����x����x�Z� :Ӿ2�
��_IJ̒���:HaL�ܺAH=��7S*O�	���a+:� w2u�L6R�K`��4��,�d��6�~ ��P%>s���61�G|�7�=��_�O;����5�u7���h�Гݲ���c�h-/E*�x�*Dr��w�~ U�0��Y�}� ػ��R�ec�ڋ���q�h����G��z#����@h�EQΗN�Fƥ
�r�����;ft��Ka�hܢ�3W55|f�9� �l,QO�Q�i��iݵ�����D�$�Ї=; ��?��@|��F���R་B9 &s	j|6ZVooI$�V[�f�K.��I�x��ƾ���sh��b���N;Ta�p %{��ߣ��|��:�o�����`�����0�v��ť�_֠0?��Wqt;�f�.��r�{�aXFm�����Bs|o�>���|�BT��y&n��J���B�AD�����Y�]2��EZ��3Y"��@wJ>���j��(�I*�-׏�C�ூ2zX�4��֘~���i��ǔ�� X�u!�rGJo6ʓ)�R��sX���-5�2���8�Es?!ӟ^�e�vg�r��i��[��ԿF��N�7��h���Y�0N����Ã���qp�Q%�~�DeŮ+�O�Qji8����G��
+Eu_j�}���a�Ҩ���ڐ݊�@�\I�,[���G��Z�%Ӟ;�O�e�;,��EШN�!�Cm�e�ub��u���\6Z*�cm���Ⱦ��-ol���c����;�����������#3�ʙe����H�9��l�V���k�� oǅ�f]IXO�8�%(>܏Z.]�2}F�5�����z�>Q��¼�*$,���o�>�D�va0Ԕ*��J�:h�0��*�n��%�&^�Sk�>����D;�6e�CH�l�7_,�sL�V��s2PF�c�S�-�~�{�aA���
oD���"�¥�1IWo����ES���}�UYtn����p�Ɲ�����>l�7yf����q�����Զ,n�&[q����zT6��VanxF��)��U-T�jj�l��D��{�`�*�Om��^m�ӗ�*Y,Y 7,�4h�,Q���Ճi��F�i<_E[�es���z_d95Z ���B�4�r�ҏ"��f�qۏ����vT�7{�~[v� ���`�J��t|�aeU;�=����^&��V����/���!������e�p3�W�l[����5y��A$tZ:Sj���(���i�\����UGO�eBuD�Q��y?�tX���%�m"?|9�h���^Nm��Jm�"��d�T�3XگHq6:p���<�#�G�\��7�o�ts&�(�N9�7ӡ&˴jo�K��Pj���j �i�'DbD��+
;����,����&�����q$��n�m�  =�[r<ER�H��r��	���������Y�1�wD�&�(d��o��}���2��Ji^�c�͂����V@�� ����;�U�������ed= ��.���;W��Q�5R�bS�����/2� �T#Nn���i�~�8�C�G`�Zֶ���1����3P��]9�)�n�������҇����G91���d,����^���a2���$�Nh�A�%|��x��{�V��n9��;����Fl�i�h���"S	�)Y��s3H]'Q�R�B�y+��B4���q,@Ɯ�}�EYE������#,q�[.�WϢ���8�]��xO�eH7?