��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������LX���>O�.:Ɨ!�}�9���4��`���ĩ>5*�rY�4-B�:����9��:�S�R��	S�u�$A'|ܼ8�22��Vk��)Z'iL��i�9��c�[7��9J�Zݜ�y�C�Af�1�7u��%�����ț�Gm�.���F�e,bW�K�{��S4x&��������	F�����|��QؔAuf��[ �ž4��%�B�sH'b݆n̹����BY�$do�N��_	���zj�,��f�U򱋍�ܤFk�=�l��s\���cK�������,�%4��~wJ�� ����֞n�89|�X������D��_u�1*�#���<8��dzd���~ڦȅ�T�ҍ(��0너w���1��IkoE�Z�7��Y�[?X3
����B�<�.]��Y��b<y�O�e���o�h�s,ue����zC+JAa��0=�#�.	g�츿�uH�l�1h�o�eJ��(:'�D3�uA���sv3j�(�:$�1;Cb��R��1%����w!��'��nU�c�<am�>V�4��PÉ�����!�����#|�������x7`s�G�l�ց�1�x��D�0?���U�ʩ��C�3�҅��$�v����B+��k	� ȳ�Znw�ϊ��$FJfY!��Q�E~E�p�>�-���^�c�90{�G���6����~�������Ƹ�#������w{��q��i$�Ʀ��mx
E�������S	"����)�A�{��(�P`�	�_In�Uؘ�D�xXjT��)��*�����<DbQ�e�d)M�M�&�s�Y�����b���nݪ���Q-b���]����
;���5�B����ĘxZ�M#L�0����eJGN���GV;�"D�V��\�����[���_�@���j-����\��V]����]La���C�/%��XrZ?%���U�?n'\�F3��(����Po�n�PyǑt8�yP-	��yחf���Rɬ��S�pW����R��#ӆ^c��}�e>��QpK�[X��~:d�z���s����KN���w�ۭ���7�?�mH�F����
�c�+���/�a�o4�_��X$c5�n�`�+��� |P�J���yEY#�b�6�5`�*����E���5O���ʍ�
���@<0��)��W$Ko���_^J�x�1AJ~�f�����fc�Q������c�Dw���g�݀.w;'��
������Bs�Y��K��*w��L{1�-�ܹk���7*�I��,��Z% ��\�h�)�_�t��z&��(�Z���
fҏt�u4�w��Pց�;^�x���c:ya2��J����`��ހ�2��,F����f���K���˾��Lj�چCn�f]/R�?�!ѝ,�҆�Q^V���5�����)9ޅ�B���:#mm�M}9�QC�c|��Ýc����yR���+�a"��`4$�i���� �3i�s�����>)�Ԛ��x~r�é�Xqz*xg�6t�pb��~s#���r~w������ڄ��ro�T�zK��S