��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q������5Ij@�fK��s�8�Pm;�̘���������RzF��c	�^K�[ߤ���p(�b��:��Ɯf����?1�gؖ�7W�uJEF$'l�q^l\wَf�ͩ[.��6��+�����3��
I���4>�h�|L���Λ0j��a���o'������o�G.J�o'&P��Ӫ� �����9,�8�;z!����Q��~���s�pפ 3�XR����-NY����.[T�����#�gzJ�qыn	�B��JY1���4R'~��-`|`p�%�BM�5
�������q6���"6a�������s&������mAz�Vv�¢��jo��g�xi�Rȹ�0�|�O�\ �í�R�).ȳ�}�X���x�����bK�0�y,��P��8S��� ��\r��!n�3|�Q�:�I����c�r���T�q߹Ḟ&���*��[��uA�3�M>�)��F�S��V��}�j,������UpĂ;�Pz9���@��|'��M��vŨi�XO 61[=d�W(h��I�X���ь�a����{Y�ͽ�:%���6�1g�uE�w�o��[p�1ވ��Z���I�RKH��J	�l���nc�
p$�W0�-Ei@uӁD�8v����-E��RH���}�Z��bpkmw����	��>���:�t�2��۞�OݾP5����@�vH�#]��C�p�P�,��bOiӓ��}˝dw�$]0kJ4)��bF�����\�?�8���V�t�# :m�a��03{��똄|�:>|�L����J��u�t��J����.mb&iw08�L�@�3�:I7�ա�N&&�g"q|��:؉0)��GK�T��'�u('1���������1�|�7\n����R\����^\o	ok�5��ݢe��N4YX��w�Q��mLo��強����q��[��T�])�V��Y%��	/�Ifت��}B�����Ic���A�G����a#������P��Z�t[-�1����� �?�,�\�˒s�Y��$<��
��'|t\��b�vb0��j#p��EX\��-�F�:��XL�O��xw�܅bh㽒W��	i���y�ƛ���
9��Q�_}���� n� �
o���@�__����XK;6zaO0����W��z$��:������uI���R�X��nb��W�8�{r7�#�de�&�WF�=cYƣ������tse���X�U4�q�@f#<z��6�ۢÓ;��₈�i{^��|0��\w,+wkrJ�I�j�9e؜i�'\��+y�o�#Iv���$ۆ�Y0��������]i�:�Ʌ]I6I~�UZڌ@�oq��t�MKp�Z��G4{]ۇܡ��>A#�v��.5\�~��0qB�;z(^���;�?���[%��B']�َ���pSWEL���tsZK���_pa<��X����'-I��߲������5^�� �䆹�2�z�}Q��mB�EFl�����K�LZ!Rrn����c����@f?�O���[[ID#�B�*4���d�	vl�co5"MM��(m� [\Y���?�!ď�L��ˋb�ۊD���?t�S�1�Ta�)�@�3��3��4r��-�f�j��T���_��͋���]���`�r�v�OYZ�k�D,n@cC���U�Ɠ��B������[�5ǂH�fj��Xh��4�����[�ġ�Ȳ��tOhI��C�=G�D�T����2u��ŉ���d����'kl�ѱ���20���,�eB�)zSo�a,L�V{���d ��.iS��;ū���^���ҖCN��<.(�#�ꮴ����"ވ�3A�QyCs�Pd����Fw��I�%bj��6�.��>�E|`%E%�RGxWרϵdm�Yb�8�G;����׉�,j��]�ط�/Q$�-����и�ɏd����]���B/�����ō֍ ��Px#u|���/9�����7�v����Cqrb�Y���*�,���9k�*��>+!��D~(4��c�Z�Ѷ�i���['#X��'�đ��f��1�}]�NT�5d�p����=�%������֗eʒ�J�K���B�b���q�%�ꭰ %�b�����D�W�hB@����^����J[���tI���yl�8i���E�I���j�ڋ�A�I"ʙJjH,][֤�#�wY�5l8�`�݂M|?��c��PY��CK\��#��J
�k!ɃF����G�d��<�Vt'��?�ж������{ͪ�Yǯa����K����x�����@*�$�A)��˰o��R�!�4t�K����Z9#x��۱�**�k�������R˪�>n����@�Q��s�xY�v��o�J>w/���lC�Aw�|�ҝV�1+�3^�MP��%�����MF2�cYadf�?SY6�e�+Z�#�O�R��^��F�˄���Н�pؾ(�F����2�Ò/�|.p�D.�"~�߲B�:��� ������<��lWI��"�6^-����l�% ��o������G(����*�i- �!.��RN�!��� j��Ge8���K �@�(���ͷ���#��/=�����b3��P��tU4�ɺmN.UQ�l�~��E9�hQi�zO��B=Guj!$8��T��i�2�	GW��	5jvnS��J�ը��{ ��L�v�\��"# ؟3�y�N�~[B�i�g�t�.������l�,.ʤ���le�.�{JK�;d�h��b�����_� ���2͓4:�e� �Ճc�9��=@\�N7�<�:�C��1�;7�����b�F+?4V��4V3SW�"�����>;�[�wRg}����Ӄ'��C�=��u�:������ZD�{ O��(�z�t�B��n�Yu�uJ�FÉ�A���ٳ5��t�a_iN�<2��\�	v8���~xђ}����-�����kE��j�^z4K"��d����O?��6[�H��
�
������[�=���s�s�b�ؾ�*����8k���i���w�f&�?�c�2�6�����=�ʍL��n�<(�hC>x�K�E���pЄ[خ1�aTg���	��9�i�����M{4Q.~EWAyCfﯭγ,�<��!=����u�M�A�Z������Y�l��:�e{X�� ©W+���I�z��b�vX&��v_��@+_�g]s��1�0],���c�7�)���#���)��ܝz�uC�~�x[�����m�d�u�Դ)?!�^�1��0�*�l%Ɛy�h*�ҥ��q�q��U�Z��GQ�#��������f��M>��������}r������u�O%6_3���~["<Y?pڽ̿�_�#V?!�9��ŽړN�y�X&��D�Y�J�q{�i`�{�ـ���5��j�	���e�������o��u���᫹ҏ�ߝ�>�R�;������{�c���̞>j0C5�B���+Y��Y��t*�f�SjN���;C,w�(�K~u�x�Cܘ1
LvO���2q�V��v CS�͘���ĽP�&��FH���".?����UUܻ7I��Z2��[b��R5�;q��k�Pk�Cٓ���qĠqJk��/���Қ{t�ϿTu��H��i�̛����^�G��[h���FP��fw�˔����ެ�D��xXks	|���-8A�4R��h��b�:\��GƲM������n0(�B�D��
Λ�,�����6=+Z�"w9�'F#�$�����	��Dݖ�M����o�c��HZ1���N���'D����@��	��{@����ԄG�o5*���c���K�� 	��4�w���G���`Ѝ�4/n˛.]2��D���{O�u89�̥�tu�|h��nɿ�ť��ܓ)N��_ Ŏd�Mv�A���L~����d�%a�y$�rà�:*�(G�9������w�pc��մ��󦑘>F+�-��T�ry�����7lխӪSu�O��0������d�?�a�E���2l��wPeP��󋇮ꉂ�|�l�^��k��3ό�5��O�6�"���h;X�}U���˛D6adoْ�#G�y-��E��P���rC=�z	8so�2�;��f�dӇ#��Q�'d�-X���;��K}"v����Ď>�;�we���Mu�Wfy�|��z�Db����%�C�ʾ�� <�<��BR��}��3�P�y����Hk{�;LD͙ȺY.����L����FO7.�ч�@܎�T��)1��s�ZDn}k���@"`�d���=tl�ν��Ä9n����N&]�;�8�u�Oy�Ԁ���gR*e�÷HwC���q�'�d>C,?Tv"���ho7�@B.������BַM�R͞�;�k�XZk�	CM1GkQP�*ۍ��.v��2,ꝷ�����ǡ�%<7�e�:Q����'�-?N�ȇ�0��_�'k_�Ͱ.�XT8�.���J[t:������� �U�����x<���}`0��?y��8�n��������kp)��Q�2G�_xk%>����Դ��/���'*a�C�μU�wBn�<u�8�A�k��o��Hez�2�꧄�6�цTŖ�������f6<L��6.]�ၗ{EO�^����Ja�����j���!R�����6�-o䎶��)��;j��a����L�XFs�oo�GץMQ�����0c37ܓ�'(h�%�B\|�x�'ԩ#=֟Dѷ�ORM�~���07+c9�R��_����h8U�Z����ou4� ��2��xB�����g62��RѧG^H���i}(�4 ɇN���ƣ�������TзM���h)��.�(6��!�<3a%��A���C�'�>_������c���\lm�����̯r����H��C��Ժ�?�>���PDRr,Kj�| `�L��E���VBH�Ԟ���v���N*UL�`����h��
� ԝ�E�x�AT�C:+X{����?�ߺ�WI\��p	Ts�r�I�/�8���Ѵ ?�&G�����c�B�M$Hp;Ԗ�p��_�V�`~/H�8u��C�D7
;��pT�r,_�c�d�n.K�У��"{��{�L��ƪG_��cZ3�K��!xXѯ�3����a����1Q��܌�蠩yTxh��CE!E+�V��3��c��&Xv2Hh�!�x���p:�%�C���r�N=��Q$&cܥ����v<�}JR�P/:���t��Z�)��� ��qW[2A]��-Zs�р�t&
��9v���C»��μ��b�p�ߤ�D"�-�B8j��*V!9�e���gLR9 �ɀ&9=�[�nN�c�X�������"����0�X�C`�A��հ-`�sb�(���b�٧Bq��f7/��4�W���2��[1����%�}�yv��W�2f���xs�p)��}�l$��Ј[֌^�-�F`	<݋oN���4�:���R�}{D?�[6�6'���㌴$��a�?�;�R��3���[�l����.
��!vf=m\��+�V�ձ���5���̟�V�X������� m'�R���)P:%i��&����`u����C�f�aS��Z��lƁ8������:w΄~�r�e7��bvN�kt�C�j`D��/`��S]��u�����J��WW��'ߺ���t菂K\i�?e�����8RkBa;�����
��(�#l/��~�x���o�ѝ�s�k�v�[!/N�x�i@����\H|9?&��-g�!x�n�>��*iYJ����T�5��N��,��q�r��^
�*Ϲ��s"�,
f�k,��2��sJ�㌝�eޖSM��1L^�&����6�uVuqt��R��:�M,p��eMz" �����ٚ� ����t/
�a3a<p�P�N;	�|}4V����kO��ݙ��+'S��|�M�	�kT���('>]�b$�۴xbF8>��C���
�e����P�&�W��`�]��oFrqgB$��-|����;��k��op5���X.��h����`c�P�T�ǝ�]Y4b6�*�Y��%��N����r�w��%��A�y�	��Zȷ_h�L �Xxr��Y���s¢&�ۍQr���
F�}VOm�t���Zܔ���"�zT����J�Zn�=��k�pYU��mӟ�N�>��[����HH�{��-�jtt���?��f��	i�Ķ�޸�lad�W���y�sH���V�4��I�3�<�F���⅜o�1��2\'w���{�@��Y�}KR�޺��)p��|� g4��=�}r$5�p�}��lY�oM3A����I��>���8`�Ś%�P&Z��k�E�_��qMEOe�S��n�1��<b�DU�D�A�%�Y4T3�o8�"	Ɨ��)�D>����f�4���K��C`��m�!_�/<dY���psY[���Lҽ#D�Q4c�d�����ځ�����-{+3.ɯ�&P�^'Kp|5_�b�8z�;@;��wfi�ji�!�i�D�&_d�M�/�+�a��W&��r�^���$N�:Z�hÞ������>�2e�Ό�ij$�l;q�I1x�m�C�����k}�m�� �/\&��ۛ�3u3�YG����!qR��Y��)C�Gҕ��0c��.�86�a㕂�ZX���0������m�v�,�D;G���Pz۠��h��)����궟J�)�� �Uv� l	���� Ğf��f��9��C��A'�-ˆf�A���g��K��a�l�-��M+j0AB}D��/{�q$3��FVD_M@��Xʶ�+=#�Kt�TB�``�c&�<� ��(��7LU]������ci��.���j�&"���W�2Pp����:.�wk
a��0��sˤu)#('�T��;�G�wZ%�H�O�'��ύ	��S
��j)���Zm缼�@,�a�RK7�V��9/����kU%p��b�z��1\�h8�P!�j��s�ݽ����D.y.=�Wk�j�����F�;U'�t4��6�#xS�ὡ}N�!���tcK�8�a���kg,7dOi�cR��U#	~ h�>�[B�	���L]��v�U3���%�RL{��By���<�A���Ù�\ -�D&&h��4{�y�/�(���Yd����x3K� ��&~#U��&>ϓ3M�ʔ×o���2��!<��"Si)����ke�l�X��b�0��a^f�&�$���5=y*��� V��涵��T}Q��1"�J�,�+*�����Lv�|���I��V(bMh<�6߼	��]�6�򁊨H�0���rb8I�2�!�4���4�|/t�����0GϾwH�]�a��}Kd�,���c��ȑd���,k�X�!����Nӎ�?qൕ�'qԉD�mw4��ȯ��Ce[�D�敏�^�$����^[8��4=��9>Wz�MAL	nE��>Nm�/Y���B́ʞ[��.�5Vz����σ�$=9�O�|�!ql��M���+�ଥ<歾@CD�Ѣ`r�6�^}��M�c����=݊�f�/�Z�R��x�6x�<�!���o��؊?�!KȩI��N���Vzh+�����"��^Fȉ�/�d:��H�iظ�햑�Lw���	M