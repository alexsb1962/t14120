��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^��������?II��c+\S�F-8Rv�]�����տ���)E�%�Ah"�C�8�����������q��Խb�%����w@N[�5��j!��w)%����8����lk4��lt�,P��'�i��yI嵮�x�i��ڀ�%$���ќ�,ތ���/�@�?x�aqIS>����L��Fi�R�xN-�U"�4�����M��%U���Ҁ�����~5�'җ����Pn���5W@�1���z8pVsPv<� ;��Y5t�R�rHM��a:�����d��eT~]�R��1�Ƥ
.oD��<^EV0�C�&����D%2��� O�![���4#<p�)�+b�s�RTկ(�ـ��Ĝ9���9q�;��kPz��%Z�<P��������(��^.�Ȕ�����l5C��ߌ3݂N0�$�3(r��G�Q�H���EЦ�u��K&���b�p`���YO��7a�`���30��d}��*��BG����8S�����K��_@��"7��.9<1��j����u�f�e�1�+�fq?��3O�VL���NHq�M��_B��<O��˒;�|��f�ʒ	�᝗�i�P������k
ƅ������ҡӶ�(bH>x��m��{crnM����� �����q&�����ґDj�q�B�p�sСTY�η-�u��6�x���>��|B$Md0&�2����n���*P1�K�l�j�V��I����g.�=�ěo8{�?��4pzd3p?�*J����U��S_@@?&�%��2�/X ޯW���P��9(SK�IW�Z�� G�MG8\���#7��[�E�<�E��#nD����x���z��~�=}d�l�0˟U߻�ˏ�~��?�/s���h|��ܕ5#�W�Ӈ�d4�^�!�j�A�(���l�LJ6��l��ϯ�O���~��koW���*���=s��"ed�%�6�n5ܒ�`v��~BV� O( 
[r���s(��zF$�n�ȷ��r�I��-ΜsF]��(�!|��{��41��H>;Ic�^n.�uE+q4Ҥ�~FL�r�CD�\�Aھ}ˆ��n�Ho/�l��O�!r�m���� ;�?����]L�7�A!_�I*�D��.��dF}G�{I��f��������#aƺ��κe�@����: ֛���FAd�p^1��!���p�&v�&Yb��\�A����";�.WP�5Ɓ��6�-��ίo�\�ѓ!������ME�~�;x� (<Wl��+i�/X�[e�B�����;�ԙA���Ta�G�سNtu�o��4Z������B�U��f~o��A�x�,H������Q�#�����xt���[m	[lTV���H%ܴ����,D���D�ѣ�R@��F��~	�&(F��!��,���yqK�ϲQ%W�����Ñ�{�(�z£!N`7� �q�$;|K1��M/L�W�e�.G�˜�ڛ�=FljNl�\g������e���2>á��D��	T֯ʜEޕOSv5u='XZb�H��	>q�-�ɓ�C�ήd���eܔ�n�8�P$��J�DZ�;7��b�H���ű��uԎ:�V{�����B�2#�O]��KZ��d����Y��Y[[� �v�f�X⧤jN�ƨ�uӴ[og���zV��Z��!]�r6��Ϛ�yV��ed#R�{Ǝ�]����#����T,<U�>z�Sp�QϠhI���5|�/;���m�#�v���9B�E��*1F�O�G����fz]]��:�q�õ�q����`a�({��>�oC�݁�Sіwg:��q����0GT�˾�(��w�7�d������KQ�U�^͎��x���8/ۡԼ%�Kޥ��X�oD��Ag�j[CKޅQ��VR�hj���N�N:Zy���qc�������N=�ƕ:|=���R�� d�Z��Q����^2e$ˇ���Ŀ�r����T!G�,&�9�|�x��&s�tQ�Upwe����dm��W���)Z�iDa+�>В�t�O�� }C���o���0�j�7s�B��RK��+*&Q��nȉ��*j�����Z����xǇ��n��T�̮*��0CSc���|HZ�B!<�.|��4� |i���
�8�]lѷ�^k��T���Q>%�<H�4\p�o�����ck��ke�Q(<���O�;5��P�Y��Z4�*d�-#��	��͢2YN
[��/j���f.�M��D�5��l"�w&V*��J��U6Dyoj�?�#տ�g+�a�S��c�����f`�;[(a�n��_�77,8ϣKD۠'������y��$��x8���N��%��(?�w[�F��S�a`9�D�#��Mr�%ZT����X�v���S\T�R%����1��`uW �\��IT��fYa7�ngLK�1S���I�>e���^��#�c���F3@/!W�\pl1M��<�)���Zjl����9G!��f}Z�v}?�:ȅ+�&W[���3�B_,Fck>�`�Ppz�$ԯa9{ޫ�U�q}k{�.�|��!���L��ʭ��ʭ�$���	��84z/���9���o<X��gP�ߐ�N+�TS�OF���bɧ׋���u��3$�X�>^lY)w��#�sK��0ei�u͵ B	v�������m�b3v�Ao��Ä=jH(/��h�S�]!���j����Z�Pk�,�jM�mDZ��,�h=a|:ʝ�*��bـ���Z)k$j4ƛ�g�� ����~�@ �(yZ 	�s�1�2���<=>{�x@��?6�D����Zr
7�V ������#��(�ږޕ����;'ϓn�Tע�Rc��ՎuF��kT�A��`���p��߅)��A��3��4��oޣ ^L8Ç��ש�9DJ��lb�]��|쾠���V�]��4g��#v�O�!m���l��I�H�m����d䶉�bX��lܲ�Ј�r�2wi+Ԫ0�!l�Љ��G����z�ܙ�q�<����ڌ<�����bYbF�x 1D���H���IUg fs�)�_��>����OՐ	y^ Ǭ�$P2�^�\._���ʂ%�J6uѧ��.�����Re�����a��*��o������j���]� ������5yg�������_�����JcG��}e���6o?�_�B�E�^����2aR|oN�W�(�,#jqm$�#>�&�`\��ݞYv4H�i1��s���Iϧ��AUGih�|U���8\5��T��a��J�ƼZI�g?��Ϗ�N��/���q�ԫ��t$��k2�!�lpt��R;�fvH�o~�Ey�[�"á�k�~f���7�?�R�9���Uk�'m�E�?�X�c��g�ψ�����,#N��-A~o�gmw�iZ�s���A#�%
�$��r��/Ŕ	�%��D�c�B/b:ĩI�8��9򤉙Q_�e>������C�[Wq���p��^��3�)�>Ft%`��O k������@�����lW�3X��b��,G���U(��nP�`�|�A�O��OU�=�gjS��6�2�����9�d�_nrV[�6�m]�t����z1K�e�>�Z��b����F޵(2S���^F�q �5�3ܔ�L��_!ȵ�DH⺈��(��jg��y�2M:mM��F�WG��
r�C߾��6]�9���dh-#�Da��n����S��|c-JIݶ���Y-�i� Y"��������7w�*,��Պ�{G��"Vb`}���`�J��ͧ|��F�*BާG�zP�g��4MK��W`Ҩ�(�AX8i	F������h�F�V,SI��Z8N]�8�
i."���7�"�eYy//Ҕ��}�Y{ i�~�v����r����;|�m��DW2����'Dh���_�,��S|�͙W��އ������H��>c������#��vD�:���oy�x��V����pz��I��ϧ4�wݤ粏��A��,�j�@TF�ے@��o�sEC�_���Z�#l�=�[�x&@�!]�5��N��m�X�(n����, p���1W�� ?��:������$uL�|_��O�-��R�� #�ax���`���怬�]��F:Q��f?j���N=��|z�?���Ǘ|���u�m�-0��=��_a �0,;
m\Mϝ����+����j�˜�K��<��.I�8}˴(Rf���i�D���$(i3� g�ˆE��P�4�;�X��wN��	�bW������H��i�s.��X�,Wb�;E� RM)IZ(�r�ܕ�NXϸGuz��//����ɰA�R��c
Yt���������|�t�x�C�&I���*?m�����%�^��%��=.�p�D����ME匚�Q@�bu5��nauo�ns��Ny ��3P�/���ɶ���ᗃ131��y�
.�e�@q[pO��Q�)�5�I�nkb$͕r��g ���(|C���R3�^dX\Գ&mB2��K1ɁpY��{a��=B_6�L�"�A�I�A&��Q^eO������I9��̗�6�5�� u֝}s�r����6}c�G6�_���`]�X�L��E��T�Oh�>[?87W6��1��BZ��,�6�P �EV�>�(��;�kC��B<��=�N�oR_�0^�Am�<Nu�s_v���������%��XI� 8N{�b7��G�VJ�K(O�䜀���)|Bs�����n\��� ��:��V[�+\c���T{�����[8�LR\#O�J�஢������ch�����}�C?� ��P�)�f��O,�)sv���H8�:��������M8g��Q/����8�������ߨ_Z��w�/'unYxm�$����d����~�4�?	����LM��M�]U:h�LH�jp|I��O	�b�������(���;z���e�Q���ʽ�֡��k@>\6�宄nrj+��Z�>@q�NNb�R��!��BBgW�僝��YW�aJE/^��X�y���5/� Z>�퇺�%��`�m��£��R�5�AC�G������r8L�Q�ܝ�w��?(�I�!H����H3c�9��Yف6��J�{�p���w�0�ܭ�'`�^�s�E�G��i*�{�SM<�k��q�5۫�`��$�l�^Վ����pu�K������S׼sY���&rl�MjS��֊�Q/'��R�j;MR
�u%����V���ŝf���NiM)}��p��*���ف��<��i��/�)6��Ký8g��v���x|<�0OL�E.3�FB�^��3�t=gX"o����_�/���L�Q��l����m���U�wk����?�m�ɲ�dd�Lￆ=�~T���p��@��`�7v�#X�*�~�_�x����Z�c=L��ⳬ5ZZ|@�]L�W�)�*�d�R9�m�(�]����_��D��-п���5W�x���wJ5��7��/6���`N�U�nPwG�ʻ�:�T�	ĭ��;�/`V�vȣ���a�,��#��ԖbI�Iފ4�p��h�)Trj0��>x��0�/��9�ҍ�|.�/��pk_c~]�:��F�&���M��/��P|��Bi���m�*k@��/��#E����76Z�rX_7���8,�S�rΒȍ�Y{�[��x5[��Q�ba���~��/��l8O�aV��2_�o$(Cĕ�<�����e��!kC��O,��K����&��-�����ى����4��T���o�8k���g$�;"�Df��趥 � ��ܹ����A���V�@�5�M`� pzH+>%��H%�+���;�o��:�v����&�΍(0�D%�[`���)"k�s�s�#����u`���؛��V�KX�}Q�2d���9�Y�X����^͞���VI]��^G�դ�(��j*��)�L-kD�eG\�/�ZA��'�
9������h9��#`-�&���������\@a�UP�ה<�� ��
<_葇�D*}Y�� {����[HOp,�.��lºm��!��O��MyB���T{ �A��-�Y���T� Z��d!f6�Pn���xȱ=�{�z�u۸�IO|Ż�b�U�`�
��Д��Pe�H,QzՆ@���O�������c��dL����[�N0���Ş7�=	��D'C�ܠ ^8���o�;@���Ȯʶ�H����өʙ��ny��/<7�rq<�o�:��i¾�_����C�BzD���)wH1����緹�'�4^/��J5{f@�	�_��)�L��/�[���;	y��Yo�����:�� ��Q\-6L4�����Ń�{�� ��Z�iklZ�Mh�a����l��+�iGל��:�[��2��qJo�l�
�?�>[��J#5gA��y�N��kE��,ڀ�J� �v����L�-;�-�+����P�R��1#BV ����zݗ#ة[��������ir�8��oac�Kt�v��>��:�M
S�fb#�g��7>����=L�J��j{`��|�-u�}�N#�0G�Ěs��uMu����+P�خ�s����+�v����2@Ώ�.W2��m@!h6c6pk�Ŗ19\^q�b`"<�7:��-	T]��_���D}���LjM>�J��Wm��%g��;������)S��P>��V�ַ���^piw+���H��v�����RM	��֧�hKէ�<����}��4�T$"��]BZW�'�!��n
�[������}��ֺ���1�
5��,܀�1}�H*����R��!�>1�Zʝ$��Dޙ<�,[b,W�z�#fv����7����w��6�we�܄0�1�U���j����˝��L�$�Jv��a̧M�w�����$�A�`�+WT�1K��ҳ�{ �y��Z�����Rju�&C�}d�\\�"����9�a҈;'�2���]���̟z-+�Dzlb���8]j�hrr���8h�������"ٵV�Սh��탺('�6�U����f�+I�4}���� �boq?Q�d/<;�M�1�u��^/}=a1tyE:�s���no���r�=4_�a>�֤�;Y�p�h��[�_��l�r9@�Vis���yO	�`�s|�l[���F���V����x�t':��5��x�7�W5*��]�\�]��|yK����${������-=R�k�N�㳐��g�������q�F������8=D��Y[���GM��& z]<��!�1ݲ�HB�.���ҪG�M�`:!���,�>��1�9����1]Zqg���������>�.�B�{`2Iq7h�<�r�\Y�em��A��<쌆�d��2Ӟ �X�X�TN&@��")��o�B�8"���)?���貞��
�{M��=~��s0�?��Ƣ��ޖo�G7�fVB���W5�_���XݕF��6{��/mk��,����ԩl�[��0D]����̘�n�g?�:)JWw#q9�@HdEO��҇�'���%{� �?۟TR�|�h���t�M��GN���� p�d�Cw�B�����
Be�Ċ��7?��T�$�1F%hj�K���#��]��XY51�0zٞ �����b�n���Ж$,��WC��h��#{��=�E���:��6`��G�����g[J��C]��TE�'�%��h�*��7�$�)x��43�Q�<�v�Bf�
TǷ�BZ�M%��''��⒨BGF ��/�w �~C�#��ϑR�3���+*����9���[��"�
F>:B�?Z�s����obOm�Ys�����v�~�Ϡ8WP2�mŹ��-I�[��X;B}��/��@<���̰��o��@���d�}�i�t����ng�o=�@Y�ou�����RQA���W�����r�ԝx�� �!5�ɩFI#11�P�p�$�3�^�(�r��ޏ)�|������ 6-6Y�0X�@ț/�V���.�)�2���2=��HyM��FY�޺E��1�����3�\�Z����.�I��>�-_��gL��/+ #�R�ۑ]����S��ǯ�:��og4��ͷ��$Q��Ap֫�j��}{٩���l2"r�J���h[����b3Į�<���(�!��Sf?:�!�O��Y�J�$P���hO�����3��4���D�w��:�|(�AŨ�� *�X�]qZ�X�K�"�W]�;�����i�94��n1�Z��w��iֳc�y���%�=��k���k�3�5|2]��_F~�y�zrCrٍ��*yvAxa���pɪX� KN����1�̈́fTM���Ժ	�ۏ���q+'����NK�-�(�7V����`��Z{����VK`��ıΏ�skA���!����i��p8�����;1�)-����	�
(��z(��s�Ǘ؁��l�l����)jBw$�$��g!/��5-�1�1��(������V�fm:��7�;����J>�`\��m��9�(�_���%�}�&-��BEd����x�%�gҏ�����,��3�α[�G�4_�M�\ˆ2����:t#3�!��k��"@�>�k+R�gҠK��VE_l�4��3�YY�Ofe��,+��[�E`��u�.��<bԋg�6\}^A
fA-ɿ䁷X�F�o���on��Q��*�ĉ��*B�u�zD((%�3�,����F�^�e���NۂX9�Y�,�WKψȍg*���;-��d��-��4XӁe�5;'��AY�����X����~��J��i��M��a�z�f�"Vr�����Ֆ����L/�EC�I�*e#S��	~N�Ɲ����`��r���ί�"I��Y{YQ��tF[�#�]�\K��+C���#sƗ��L��� .>f�7�����X�tL��J�)tKl7)�/�s�m_�MN�p�
	���$�s��&�x�^��ٛXe�ϐ���� |�	r�����l(HK>��hF(I��[�F�$����{N\J��4����Inp��Pԁ=�l=���ʙe�m�V��Zp���#��] �T^b�df���,>��!`f_k#�<F��`_��Ŷ��P�~u|�aTd����"N͞�_���q"��୊�E��`����L���>�D*�(>����K��Xɑ�:�nPk���3G#�($�X�!0o�T�<`�e�VB��OIu�5QO_�����,���J�p�q;�ũ��,�'>H_+�1��/��,t��I���a�����.2�ڗ@��?a#��,� "�������7��=���o��Y�20�WII�7�FB��18� �C�h�y�Z�g.�ܜ��t�P"+�"��R,Ԓ�Gᦄ�0{Z��I�� ��1I�H+ٻν�	�C��غ�G:�FKRfdy��Ȩ��2������mk��CQJ�v�M{�++4��"�s���o2�}睞q�t�"��!��÷.@:��ж��"����V\ȴ�$�gK�.J�ʜ���FtH	JQu>#�x(�%w�!f:e���])H�-���1��6_�|BE����Wu��d�����]V��)�4��x��,����_z�_E�{��pi�p��@�Duc�-�5ሣ#�|N�� D�^n�Xe��#�6�s O&p5��*��d��|�,�"#cQ���0��d�;v3V*�P:�rՑ��]x�Ѵ��\S�P�l�^=*g�	�{�'ǒ/�4;ir��v���F���ζ��T.q�<�(�.�{z+HQ��i�wotu#�w\,��:���p��*����#-��'�`�P9K�n}�|Y�͓w��6J���������C�szY��l¡ L�����Xa��d�_ɨ���%�|E�n���øګ�nP<o����5n1���@V����:��q��o��%n�do<sy�\b&�$�Տ�.Clb�c��e�ç�Ǣ��$������.:)���ʛ�����#_��9b�2�����������G� �q)��=�"v�[��V�cR��!1��^�O����ˑ��7,b�R%b�l�BY�a��w8� � h�]L�l�yz:À�[���C8Qq>���.��?���?�pF��	ѷ� D!F(��1K��F�g�Q��ں\���(��9�؄S���[�Ic�!4i�_�Ҙ����3i���չ1Kf��W�>������b��9�
:��Hf�����fu���Ĥ��_�{��������r){�?|�=]Z�͕Â�Ĳ`�c����!�*r
Q��Lڼ&j.ol��ʍC�D5��">A"�3N�v���nC�ea<�voQ�ˠ����1��@����91"/���۩ʒ�Һ��_���� oY=��yy^�],^yƕ�Ͻ�Q�� � dՁ�`�#���}w��1 `i�gn���:	O�I\�6�j�ڵ G��u�m80�0�u1�g4��$&G�Pt19ֽ�Ek{N{!�F�l�ȋ���\��᫫��rq��I63��D���d�m� �L3A=��=�2>�˛cIF&�ad��-�
_u"�x��C��UX��X����Kf/ݭ��w�uq>�g��0���ɱ�Ʌ��W�X����!��S;��h7��H�A���N}�z���c{<F�	tR$X��9��ܟz�ְo*��d������p�Gu��p�^�-L���44^�5�{��!�L��6�c�i���b�ܺ��=��Q^���o��e6���Fo?GAYNݒ�b��/݄�1\F��i��
�����E�T'���WP��aH����/�	��S�oӥ�������FD7iHj�<ť7`F}R��$���`
u��!.�+Z+BWEC����jvk7{��G��>K��Bq���ķZ�����@k�����2:V�:��ic�ס�������ֻ���7	�pe���O�0$�h��K�%�::�����UG�&�Eg�<Ku�;d�s�j)J>d5����V$�wd�M�)�f:1��%y�AQ������$ с��)V)�y ��������j���L���\hQ�o���-1�-$M�U��4EI?E�o�F�T��Di��	#Z��X>ֈ5�KA��9�ʭ����ש����Z:�R����nM{�N�ޢ�x��3��?��R�׸F�=p� =�����Ǽ�`Jz�3S���T��x���?������<KO���.z����sq@Wt��SL�\��t�-�u�X.-���s�(�K4�)H���ƀ:Mk�lW_�t����	}:��o��	�K-k�S(���R��7Χ'����.?BXf�j��l���t�[�C��;�D{
�X��Ǩ�D��qGʞ��N��\�x	%N3=���y��܁�����Ƿr��d�����B^�=��yw�X)(B���_�r��譛�������O���y���-���sGm 5�,��
8޷8���E�.�&�c{��*6�,QÂ�4��%�M�R�8mM�� 
haholX��1�ǀ�/<B��Af�1����'��%�pNvmuۇ`t�P�`���-?�\,Nܐ7Gm����^�k~�_��IF#�?;��F�r��HC�j��F�s�+�P^[e��|4/}m:���i���܀�m�&�:��iEqX�N�u�r¤0��3eV��O�����h�1�]��<
m5�q_x: ��eZa����?1�1�>��h���0�H�#�WR� ��G�R���M� -"�$/��!y��� �m�cЭ]�75���>��"��4{e]S���;��d?H5.��ģ����*nҚ�]��?՟��¹�V���*��$���v��o�*��ӊ ҉ՠ�07��k�r��aDr�ޏ�ۑ��@撅���)�sOb/������h`��A��#�f�\^8����]�Ak1����:�B��klfלgP]�����fL��k�lC����IlՔ'�oHHo[Dɐ��e}��W���hZ�F6���d�	vրN2���l������*�vm���D���.�t#��98�ā���H����A�)�&�EOc�	�H�v�'軦��g<N�w��A�1B��OY�U9�gH�>��JA"��Q�-�;:�V�>���Ů�9p(��+�?ک0jB1����z=��d��b�fһ0LS����נf}�ȩn�/Y3��H���থa��U%Te�;"g���	~���Hw~yG���uY�i9D7\�\�	&����K�v�$E��HG�&�K��$~��9�L��g����?M�8��7��z��&vQ�|78T�
:�i
�P}�y؝�bl;��{�ryM�\�N.&��?���3�f�39Z�����}����q܈ٔi=��x�É�]�b�b�)��b&Yx��Eg�}��Qi0}sָ�%�%;�R�8���ۢ3�'d���q��HC�g��m�_<xs.�`J��7'��%وp��==�+\e����p$��x��q���w�z�0Ӝ3Xw����P�	��B�Q�qY�maW\����E�ڌ��2��=iQ�t�f������'~T��2Cؖ�(���G��.����i�JRiڨl��\&�{Ͳ���J�:{�)��B���A��������h*�4������oDĒ;�ZC6�eT�%s�^�FO��{����2���)�尡�ز��:��a�f2K����3F�#?�}&�S��琾o*׺�Tku�U�l�3O��QWc����� s�j9�AP�s�Ǌ�6�,�&O;���E�s�S)�E�{2{�r����A�Ju�������TEb#�D�;��Q+(�e҉:�%�����r*�]�΍$�Ê��� ��B �#�����}Y�h?�>��C�xD(ǂ���~�y�i��7��"��0���Uhx������ ��JP���Kw&���)�c�����5����HY�e��ڢ�n��$�8Q`DWA�b�4�]��G�z��;os���)4��@N�����3��L?�M������+�kS��Tݔ�/�٬@^9%��f�l��k9'��dF^`t�K�n���Q0{��f��?1���I�A�A*
�^�ۮ�j7��H����÷ϔz���qd�GN��Xωl�x'�8;(�C!�SQHQ>�×�����:rl�i ����>�"�ꆭ�|N|I�73��>DTs���fY�������q��Q �	��/��� ���u�����՟kǉ��y5�<�4�?�!�({����X?7�Y �7�KI85PYע��@�ǅ�����w;����#����+@I���mp�-%���+��l���j�S�����A����c6K7�j��ol*��PV��Q0�䥂�b��Q�rӆܾ⟳�U��6�1������8M��;��G�?�><kS4�������e\h��7G��̮�Q$[=%$Q�ϡ�i)����d�)��n7+�|I�ܢ���z��]V���Z*����i�/�Z[::���M_*f��^z�zВ�w����Ώ�G�ȝ����0=`|� q~�~ ��1�Z�C�wŦ�_���`�	�!��噿]�~:w�b['�J�'T_1���4��[Yt�	�S�ü-���@�����JJ���rS��9�䝵�ߝfZ�[�C����*�,��9eY.[vx��ln��C68��;�.<fS�[1�j�'k�mh	p;'��Ņ"%�c�݊MMcJ ��'Yq���l���ۨ�ja���~'_��N~�{A����D�>):��ЃeL*�X\���Y�H�F�hj;腌}P�F���`R��PP?]�.(��2hARu��Sj�	(�q{��Z~�CS�|�hzq�����&?�O��[�u<�_9�R��,y�KD!ra��/3�$hX��ȱl��go�y�,L[2���s[�x(Fcͳi����7R|x/�L_ծ��־᪢m[-��4��Cei��A�l
�M�4�!�l[�C�ó���Zc5�x�x�q�����QFq�I�j׮a�Z@L��������-Ta�Ԅ�S���7����`�����Z�	:�*�gG�͏L!�o�pG�;�x?�����Q�.���%s&]�A��!���2SK�6�0S4���AO���Z��t���E��r�+S��W*@�!�����t2!!a	�X�b�|��
#�%D�&�b[����� B~at��x'�Ȅ�Q��!z�m��#�¥G���OY}�nNi���J�>�>��F�K�M��??���D:8���`G���D/R,��LU�S��N6RԨQ��PSo��WQ�'�uUr���p��0> [C��gO(X�����S0�4v��{��T��|��C5�,�f�O����(���K�3N�-�/9b���n�U#(�W�QMX�b%�����|�^�j�ol��R{m����b	̹�T�.��qCB��	�ԭ�t�å%,]EƷ�4_�&R�#�7V�,0���/5��-h��+~XX�*�3�*a2~�FL��Y[֩���ah���b����A܃��i���:W�y��nm?�p[�&�G�d�`��8�b�����P���ب���d�MA��/�<�"��g�K�*kl��u)�')VmU"�ƂA�vEI��y�^�H�
�����v��(��G�߃w딸 {��^A�Zƽ�s���I��K�̟aK�tM�7O�Ǯ�J&�܎Ƨ��U$	@���K�dWg≹K�vxb�|�+Ӵ���&ˋVN�^�B1�acPu㧩.eyϖ���aT���B�ƚ��7Zh0V�J��7��0}�;(�����D�nK�D�;wD�X�/I���x�fڃ�	]�Z!�J���a�mWFb��6^�	���צ���!�vG˅�����'��`LW���T�{���4�l���_A�ξ-�bf��or���Ҧ��yIp8�y�# �𜓁���Y�<��yy䡳�iM"�\x���R$�=�}���7�u%��ǿSm��!M
v�b/�$tޣN���P��$���h�z�s�en���C�t�6^=6چ��x[�C�ި�^�c/�Y֤����~ *��X����dqh��o����	�I����~�J9	�Y��Ǌ��.K���j9�	>%�����$Q8.�'P�P1�F���ۑѡ�f`v�������~�LÐ��v� mS��ß��+�Jg�ǉo 5���WW��W����a���+xmY�aY)ݮ��}����ʰe�&ȂR�>��1c�����h����?R�*���ٲ|Y`��C�1y���%O*`��?lib��;IѶZ�Z��}lA4�It� U�����m�ɏc

�!DHi���A�!��'���-���J6C���e�lN��s%���toL��)�1	�x�P�J@M�o%v�TK��z��b<�7�7����<���(_�l�)��c��?(�2k�E�f> ��{L>�!��N�֞�F�a�v@�����!A�c����Q=���t�e ?�^|O��#��Z��L�Nц��L��1�i�ލ`�F�O�W��܈/F�!�{���{���_�� wM�;	'6>�g���ԕbY��2J��K������؍��ݳ�0�ċg�,���^�!lbA�m:�Ej9���QZ��o%��H5����esD�xz񇧻��M��;`K�����8<�D��N�!؞�ܩ	�d�)�;W�*�i�:s,��k�/����,�� �Yn�I��75Oed��\��`�&&֩;�d���	��$�6-��xF�'e�<5�W��K�?�?q�E����8Umҏ�x�x.��5KTɠv�����^����<c��(���to|m:���
�bK�4-
A@�ŷ�W�$�E#������)t�o"�G���[�v�8)}�X�3������><m,q6>�囡����0��@[����(���"�݀[7w$������� %I���"]�T �-����$�����0��<���ĶE��Q�K�]�v�FGl�7�0	s�����j�T��<|�k�أ�Q%Єq�=	@W�E�+��J����x#:v�ʼk�B<N�z),�Dd��Y�!�bz��w
����w����
r�xo0�X�mT~WZ�ǅM��]b-&��Ee�̬�3�B6ѸG�rMg��f�ڃ�Zr>C2���h�N�qĂ�p����� �L��n���'�s5�I��C4:���z<����������S�����'
~�k����/4�g|��)+��g�Nq�1��ie-���>�����ײ����A���4S_7kh�#�l�/��+P�����;\q��!�1�����M{��*��Wu�˰.W�0&����(g�
肯O$�v+:�*�����&��Cc�� ��@�Dv{��2+/�D���A]2j���7 b��3ֿ2B� ��2K�H �\��Pt��s,����{���6G����J�IR���(yv@�q�se��lꙿ,&�}I��A�GG�4�
��Q̭M��ާt�)���Z��"�����Q��Y��~��+i(� ��gS[��54�-s��Or���-ĩ���A������P?�m�1�O
`�O��O�[��2�Y7܆���!�ח����Bq�;E¾}�P 
�$!o^���F)Ք"2�h�8��^+���p��zr(Mm�d��mg*�l�o�h���3u���k�7�5�������lK���c{��Z��bR�B��.�]
j�O`�i=x?	��������V!Bɺ���Y�q�_yC���Ӕ��*D [�����TH�Z�����7��d��Zޤqgc�v1�ed��%�%�	@=*1 4# ^^�+�����~f��R��'��*�T�8���u�R'�[]_��.ۺf�Y��Jg�ˬ��jx&�1�/�j��<�}^�
LY�&+Q�]��Ȥ��D;v�=���k�*o%�s�G�j���mFL�9���=�^a�3�Ո�� ��ӛ��c��*��D��Z��ɯ*0(q쇴�嗖u���ۊb�;x�\"nC& �LOx��}�s�5cg�d�bYgrݰm�C���β��;�`z�A�Y\���v�[_��y�`�ދ�����h�i�23z��D=B�l=�t��C�UB��/8�+a��������9L&�Q(ed7�w&H�� ��rq��<�x����H�U����zݽ�k��ѠLT?Ι��R�q�3���F�"�N�Tc���a���r�u��fu'������b�!B�~����&%��=�A���n[�����BR��}}��]$Tj`o�&&f�	Ҳ� Mļ�-?c������ 7g� �iN�ڴ^�&�ק-/����vC�1{� n�/�OV���|���L�����l����3+�W@�T�;�����FD�����_ +���9�(��4��D3V_l��h �C�#���=���v;BL���*���Nx�)���M2����V-J�yq��z��e����N�^�x\��n�X_y�y �:{���Oי�3Sd�:H��΄�q�s@}ڹ읶�v�x���J�
0{��2�bJ!8�+w��
��P�ʟK�&#{eX
�̱"�!Kl]k����9�ҝ��{ɔ*��p�Z�#t�F���s��?���~v³� v�Uٌ##^����9+�5������5~�V�L��a�BD�a���7[�"��E%�6:N~�
5t9�Ab�4ѱc�9d��o0 �{�<xv]�!�����KՀ/�|�������h�K�x������UZP��t�{%�O�ߐ�o��z�N!�����o�J*)�,}*e�X�J����e�S��)3���0#Z�|u��u�︍�N���
=����r$cn���h�#��ܔp��)�:HU�n�P��Ú���kz�yr�r�zB"'KPz�T	^Sr<��Xg��s�/�-����݅Zধ���ꅘ�k�.��.m�� PH�䚐n�#��D�,�Nf,����|�drÌqZt�R���z�����*$��E�����"Cs�=�x��/���[1�G%p^��-�B͆��G������d�0�����T��i��,]Wg��b&�^?6�ڑW��2��kg4��o�6Jcݮ��dY��� ;����sx�P� �5���?�4���� 39�M�8���*X�qAPVޫ?)��������W��>�_R�Lo�6;��<Q�#��Ȣ66���ߓ&�\�<��'l�B�4��K���Eu\D�m��MP��|_!�G��q�ڕ��g~�@{ݖB��j���5Ճ�*Vm�vq7{&����6���/z�(��5Pգ���|�|:M�d +�pr�w���{�O�$�ls��;���
�ާ?���Ȍ�>i,��=;�	||���Q/�����VP{,��IOIӊ>�M������!�»i����|������}�VstN������-K8�ό+T�[�m}��An(��+Q�0d�\5�*�iX��ߐ� ���2���%,M����^�-|��O�#Hv'�UfS�L-Ĉ�Hu�B��E?�c#�o����/.�,��a[�h����`Dt����@e�%��Qe�8SĎQ|,xM/զ��b
�ga�;�܌����	�8¾ׯ��F���!s�����_�H�~�8������[� ����N�wRb��V4Nr�NqC�>��)傩�1�)�^��,�����,ӥb,$����M	#��D��k���PZ<y�L�Hp��y�*?�<T��epڭbb�%"IQV�pڴ��%Ո�"rWb���)��bw���g��M�m��]k�3��T���^z`#�];�rh�*�֠�}�+ ۮb�Xi��M���� �
����2H(�g��~m�Q�+���,0���@t������O���D�Z���g�������
5τIP��s�pL�i�x���c�uxY�$ô:�m�vo��y�Wb�JM��%HkywM,��W�Տ�m7����E�y6O�:8ӽ���a6	z%/l�~d3��::�N݀j9HXF�_��8�ԗ�cc�!"`����W���	|e�
����ݦv��tsX�)I��IK�x�|���=�3�|�l�*�QW]P0D)<�Z�](�f�n��9H�����6(�[����~��Z����n*���G��'V�VI�ת[�_���������@����Ι��}xit̆ʠ�E��$|�u	��7gx�`d�ǐ��mX�>��Cl�
�"j.�L���|���`$�s�Ո�7�b���K���Ъ�=��M���wʙaT�o�}w+�e�ա�B�������0
#Nſ�+Qm�K =Z�n�=�9�Wa1����pMd���igZ�D�5����\đ�z3Յ)����*]�Fk��ܛ� ��ٱ�"H!$,���x�=����Xnж�u����wm�[���Ѷ��rs�	'��wŗ�
~���s��a*�;�j��JZ��M��=`s� D��Ey�,���7��ͫ���6��b+
`E�*�}��,��)����=� j97�].b� J3Z	���f���_A�mH˃���5dZ�p;g�{S련���n��cȶO.{4M��6�$gVq�E_|�>�t���FϢ&� _�r������Y7A>18S����-?���{C���ʔ���xh���H�y�S�|
��?��i���؄�+��4���Y�@L�[F>�"�ꄠ!��8w�"/�&pn���B��������_�o2�J�#\���9O�)nf�W���T��_�w�A�im�^��Zx;=����G��n%��+;FpT
�����{�ow�Lc�{[6�����˾���(�5v�v�'F����t�����`�қ�d�p�Q�,�4�C�3ѯ�HWH<��Bra�|�Pùh��2VUbg~�=/x�u�{	�W�p�BK�
s*��O�������V{V��j�X�bKi�Y�렾$����e�@j�t�h�0MK��],�*15:���Hk;Z�3E#i��_1�3!f{"��47����I~�a��*0_�I��3�� ���-�=U�~X-� ��b$b�K"�,:��_IOʏ�;�bE�=�h�QQi��$[?����&��דl����1e��4��Z_y�P]�ϼ��`��U�B��ċ���na����q䎖�__P�B�r��j���H�\}e�uM*y�J�}ɶכ�� xhfC�;����	�z�׹	X�"/�b��J���o-����j��#I��	M,��~��M�{^�ZsIgq���3ޥ5y��E!Y��8���y�G�I N:)	��ӀU���Й��՘Ll�9j��{��8;*�e\S�6K[u��F���ncO�Iʼ2��%o�5���ՒO/��<z͓�l
F5`��=���;'hb�|3zb$�(����pE�F���D��!�y�Z��峿%R΄
�o>�߆ŰK�h��O�{��ԩ�����@�@f��5�=B �ѝ��ָ x{J}G��s��;��e*�t(
FӠ����p���UG����*��M;��O��"#D�n��/�I�n~ԒY���J:(��yf)R]b��(�6Q�P+.aҗ���״4���7�W_�s�^gd)�C��Ee�7��v�����ij+$����j��c5N���Nq<��d�d1;e�?2��Ǘ��DV/C�2?�������p���.�ᰄ���Tڌ�8cŲ.!�I��M��+?q�?q��{7��9N���M�nHy,o�Ğ� ��_G��-Z!JD�W���I�-bd�ѭ�Kdı�9���aH^J2����D�jt8�;�z3"��?�kr��_���,�'.���A�����I�>N�j��lcʘ"�s�,f�V�<����93.tSL��
����&����������ZY�/���hDa���0�(-�k��l��W��9'Ń��!���r�>"��
�o����������]�����jfZU
�%�3�]�R'�0��̽�E��k1�e��M|ܰG�5�����%q�~h��9�$�|�a(�XG�K�#nA_.d:��L�`���?a�u	2y�%,ֶ��i���gd׍c[Y�S�*�,�L��S�8D�����yLt�P�h�۲3�2�:��ƏwJi�/�Ut^ԑqïo������M�3�O̍1�7���(2	C�{:7�>�ё^Qc_gK�6��2R�h(1�އ������lv����>��P�!�,���yu;���<��mj����k�<�_^#g�e翦��o�}��y�s�o,��w�����PP'(V�\�0տ&�f~C}S���s��(MJI��3�D�r#��^fM	��f(�� �
Y�o�����X��7��ƨH�v�+�$����>��43�|�MP�xu��|�y���o����*��>�5��Y)R�o͞��Y������~�Q��i�Qё�
��.�wX���>ڍq}�;Yk�ϳFNs8X �ƈG2�l8���
Q���$�nN0���E����6��q��l���%N����N�g^��qeE�dY�r�)���S4K z�-W��=7뒕��f��مV�l�P��?�)��Q�2u� ��9>@������M�B��)��{���:�+1�\x��<���X�'Z�T��S�qmh�0�v�������}���+7��!��Y�т�o2t8u|�g�lZF'd����������~r��8b[��m���7u���yS�'K��_@y�,��"�� H��	0@�<M���	<���: �n7��=���t��}+ŜSs]�b�Of�K.�-���t~�B*١R�x��6O.���}�K��&����M��i;3/�-�p�/�`��?������)J�� ��	��?�	��.���#H�;q�w�	ʣ�A6�F�+^�y$���d,f��&܈�Z-�n��76���:�W���"{�2���Gؙ_[�F�-Ae$��!���L�M���&pR�i`����h��k��z{�fB!�9�L�z�8?�s��k9��V�H��&f#d�;�]�e�עY<(���K	�҆��N35ۛpW�������d�Ls��ҧ)J{����Uȩ��9�{¡��G���o�onk-���4��t0���ٌG�pyԹpF*��}Ѻu@����|���[��#�y��q���)h�A\��g0�2�_j}Y�#�lԟ"H_��ᗵ���L��L�k�F��X����K�u�:��BV�cl̠6(����R�'uI��g䰂xr���Y-�L��*ُ��8�e��a%�^J�D[TR!��C�ɠ
����`���oz�)�;�	����Ő"�?3��d�K��uD[R���q�5u3G���c��[�<GtW����\x�x��ś�gb{�kr�=�W��=;Q��l#�Թ� ��՛�������D
bGs��a��W�ݙO]op��kгV_eN��"KwWpm��~י|-�FE�<)��I���?B�l�JN��#w.� ����)YU�����%� tKwi,��*߬�K�g7�`�t�E�@*>��J9ҧ�t *9ʮ��jb(`�
d�����Z���ҽ��I�/���e,��/��j$W.�ET+g���˘r����%2��I���@*�w_L�9]T�}�e��TX�εk�^̌Z��)y�I�Ŗ����1Q�`ޤrn��դٻA��LM�9(W`�i��+������?ahKip(yT�:K� ����,�����0��'Lk�Tc�ܺqܛ�?����{�u4 I�gW9��PZ�h����n9����g�	p
L��ie���1���y��h�}�����L�����(/6����7���M�����w-Llʡ#���Y}��l�
̙�?pmkHՃ����b��J�$�
x�ه�t��K�܇�~�܌wr�s�7���%�	,m���:�
����%��h~����j�`㬢L�G(��?3���JdO�����)�);/FK�M�^� ����޻V�}}�_�@������&(3x����7қz�ݲ�߾�Z�E r�h-�|��}�
�M���ٔy�Н�����P6��t;*�r�1s�ož_� ��O�+��qz��MS�p�A[<?�B��
H#33���;b���q�D�iG��<���]�{���!)�h�ʥ�e�R@D%3�{"�^k�}���_dYc{%�R[ltv��ߢ]��' �mʌ�:#-�cms���0l�G��鯟�L����߾1�+�TP�8a���c�\��0d�"/�e&M:�=��,H��0�7��V#�\�x�m#�O[<�����w!t�~	
Pyl�LUWE
��o(�ӑ��B��E�]�&������?.�9τ�njvFu�ǎKY�5�U��m�̏�罙��ٛ��t�G��Q�+����*�9=��tGR<����tZ�?$�_�so���C[��|��̷��l�?K_���Z�}���}�L�{aCC��&'Y@�$��5ç�qh����g�����D���A&�O�<��T4vY�}��|E�q�e��3;��YI�֝�ڶ)�w
��ǹ�1���B���\S��y���n���Mk�����4g6�	[`npd�����S���UǨT\��xE���Ǡ���ӱ۬�_���b�{�����DY�'.ʭ»�p�}���( {�-���*N���}�Eq�`(�8��5�r��zO��9LΣ����k8��i��@hx0�_�JB8
���mv	S)"�+���.#�==u�6a�Y0�s�\/G��	)6>p�+@4JR$D��8���}O�7r"�SE|�ݞ R�ܩd�'Ld��EQp%,��A�~4	�q>���4�DgCL��U��o*�����]a
�3��Z��v���#��Kcvp	��>�z:�e��ǖU����+8�:w�݄(�c�
yߥ����e�huK��AN�� ���;��H���7�^)�3�r���y�����W�YMa�����^ᘯE��÷�����dc�`�l�����q�y����Ɔ�&�iL��-���0ݻQ�r(�r�v��k	3$��Q� �TaB�з�J�c�`�ʀ�Z*��\�1�A)��<��h��.�<K
�׻-����'��3��R����аg����[��ڇ�h"���n=6앵�<.%��8�Y�D�IT�U.=�n@�]L�L�4�(�&�rn���*��D/�Ax(�%�k#�_�;��i+�8����F��|O�s�/���]���.�w�[<	Q|��T�
-3�/=������ڤ�e��!�|x��~Ӄ'()Z��[~��(�����!�����u�+��v��L�H�!��&9�"K�3d��4��؞��-/��1���p��r���r"a_~<F��P+-2�턢�{~'�Y&ɛ?Zz���������:fx8������:�~_�秆�l��B�%P~ڭ���%�t��H��p��&hc	b���t�ڪ%�@��|L-<(ﺯ�M'{�y�p7[�b����� ���dB�d}�������Y�#�}i��p嘄&V�j����� a]:�u�j�;p��H�� '��h6Pk��ܔ��{��9q#���ˏ�l��Ź�l��H�)C�H.hb�6��uF��}���(���Ȯ�*��TDs�|��6�F�l8I���b���Dʘme�vJ�'M(�1�|�eLV�d�V
���R�u��x�Tv��X��|���P�Z(|�e�(�>�/xe�L����� �-������4�E�w�pv �lp����s?����K��@s���4W�;���:;FR]��B>�P��Ҹ�r�y��x���q�	��\�$ہ�d����}� B!wr���S�y��[D%1�`^�i�ʅ&�ݞ�1K�t!,�[B=���2I��"��
�9,!loM���4c�m))�T-8#u{d�>�i�L�:pl]�qE~m�*�b	����:��y^t�5�*Iim�ck��SIX��x.r��ˍ5�#�_���t�d�N���=:��9p�]է��ʍ�_�㕼�r�ߙ#���ZGp���GF/�t�ݰ��~�ߴ��	��P8@��;5���:��u���B~��{+&r���#O��a�	�~
d�H�N�{�R3��g4���ј�	�ca�A�l�Q�O�w�A��1�8���p�o4W��W�K��+�����~�&��ֺ�+�)��]�W9�8�g9�����3	��|�s͊��V�H8JC6�3�M�'��W��AS2l$.�@�UD��FA����o(�lV�7�j7��N`p�����ݣ�{~��]�SD�PZ����ņ�*��^!��T��xYT��wL/R��DK���Ɲ5^R��\dJE~
��o�����gz��Xnj�m�+2�ZrX��W��νsB�ٕg�;Zo`Im�W� �&��{0j�:��,�.�Y~��'�b�<�M�%�g����0���P�qdJC<Bnԛ�QyD0�0�?��4�ϳ9�mn�E��ʺ&�MV�����2�Ι(%�RnoC�1x���y& �>����2��t/+A���Ae ����]*?�^���W���,�Qp�z�s��CS�`��	W��x�f>��d3�O�08�5ώ&�?F&���1+��.ȣ	���XzF�ڷ�\��E�!��'Kี�|�!ab����d�E�(��Ķ����u,�Hj�b���ku��K�l
3���5p�Tn.��,��I�وꤒtv[�5%=�!%�3ؿ�ܽ#;6�)����3n���'�!�!�V�^D"����� $���:�L�R-�仓�c/'��V^d��mZ a	&��D��0Я�vۉSe?]��z��̗ڄrG��+��;������)�-��E�3N�\"6�'s������p���:�?�P�|&�]��x��q'����U�u�"ۄ�fe�Ϳ��H�-�����DoD�	D���\[��l$��-}�1}�:��q�;����<��eQL��	�!3�˅=b�Od��Lt��=,�<���Ɨ�� Q���M�&�B�E��.�i�^X 1�%S����`v?l�ȯ�f�m2z&X��fm�=q�_p"�q�k�iv
79�މK�ytm� ��	����r���m;>�ñ�ӦI�-��mV�������|�J���Q��P$�z�|L������\A{2�7�/Ĉ�$���5d�S����Z��5�l�D�&�g�`O ��楦{z�YҎ�G����+�bL���M$Μ��R��ik*��T�p;ݨ\� x�͍��:�>5���'.�y����l����z_�W�:����.f�.�߷�'!DR�'Ga_VY
�)d�2��WS ���B7������t�ҩ��r�����p����-�����vkKH�M��KLO4I5� MkB�e��P��q��7G��h1-b� �Y�����j�cߵC'h��x��n1j+��S{|��E�3@5�yϷ�ӵ�\CUrwm�� J�9����̼E$3�X�-��d%8�0*QJ�CU�}3�Qr�����}��|җ�ᬜn��g�؍��I�kL�e���~lT��z��bܘ,#�8g�|:R��ِ�Rȵ��r1��ʗ{Q�=���8��c�W��Q`�ݱY]%�i��`t�I$Ci��<���#9� <��='s�d;�#!���ؙC�ot�]� Ct}	�����I)y01}'�3ꂝ�>���]�+���iG�z@�:�Y?'X�мAr�W��fo�1�<M>�J��vP�#�v�SiGA�w�f��qGTp��9���|6�>�T.f4����`Y#��ݓ�4�2����Hw�O�8K	���R�z��62��}�U�L�oi��T��rwq��[���H6`'�Jݐ�u�ݿ� u��� ��Ŀ�}_N-��PI��[�[dbXUzZ}�!l�����b��N���+�`a�3� ���3�Ā��P_�$&	�,u�ɋ���llUe��<�b	�x��~r/ƫ�l���ft��`���*F_H�&�`�O��,\���M|�UT]$����+��0��*�ǁ��)�	��H#�����(��6�*��@V����;���[���1V�	���'"#��G],rI��W�����?�z(?�uv�� )�"�1>,���Nd���al�
_��HX4����II����Ā��tR�Y��G���"���+�To_��X@��$F]	[=�i'"l��\��C�[7�7���!���l�QVf�}� y�NU�K "İL���qO����� �T�q�:5y�g�.wى�uqI����ߋ����I�
���H�VaiA�w���:�U���v�$m�7��S��`E)`р��/��q���v~n�3C ڝ���_G uL�L���>�j���lףb:ۿd����!�|���K >�]愈����\�>M�å'>ډp8�&x�']��j�d�>���I� I�����	%��?���H:`�[_����B5�Ec�����y�&��DO�oS�/a����a�����"W{Ⱥ�}�4�I%Q�*�����	����B=bp�Q�bcP�C5���b�|�#������������Bnz�TC}�Q�l���+���������&�/�h�:��Gt�-oRu`M�z�^?��f�tT|�̰�A��V�C�k���~�kD����_�x�0x啯K�p�Q�+֗��$/�q�&���',�������z&d;G(}x�o3E_d�>uq�����!@����\JR���� ��4h$z���D�eIx^�5�Sã}����gT&�H��ko�'��,rv�Y��sd��u�/8���c��v�kC?� (ǟ����Dp��x5tjT0�k���g�����y�v¶����pj�4�ܼq㪘���=܈�����p:�����=9N���)$�d>��`��n'���z+�Ƨ5��_�\B�W(`@~{�� wT,]>8T,��~Ϥ��ۘ�P���k%B����E_.�,��� ȉ��m�t$x"_�5���vғ�$���#c�� 7���sw(�t)��<��F���*e8Yk3����R%�	�eL�lv��&
$���0j �(�Njm�q���e��SA�>�S��&���n���hV�ܙ8k�ӷ�e	Y�O��r�7b�~���d���+Yů���H���ǯRl6�=fŬ��P��i|��N�x���}�ء3�՘�7(SV�V�0�S
�e�w[b���'�8ߌv
�|[MD&ͩ�~V��~>���X������-L�� [?Ή[ �+���> PO�G҈~�f��ւL�Q�'ڻ�Ϭ������f��`8��y�c1r��ي5�S^u��׉\� �Q�$Y�k�ѹ�v04������J7��⹘!��K��.�x�36x�ˡޢ��7��GȚK�MN$a�;#2�B;���ώ��O�b%k-��Х{�#B=Ķj�d�KG��M`�-N; ��{ٍ,��0B��'�f�f�'�n5���G��O.B�y�V��7�X�U�o]ح�>�*��G���ԙb��gq��Д�Y`5�f:���׸����%�N^��Av����1�_�5�%��u|�����8Wo3l�����ODM�H!x�_��q�,4�ևБgjW�mE�΋J��y����ᄟ�p��1���<ؤ�{]%�>;�_���~����q3�/06A�*����+P��=-�&=TB�֏�]8�:��V?�n%�_y�s5%O�'���o��G+���������o-�1
9W�Ji�^�t��L1���C�1(A\w�s�
�Y��%(
��nCGCoxd������w]�k��K�h����<��-p��yr�:!s�H���!S�dbFX���C{O�Ggx�LbYM ��ptB��L�UR�b�5��Mp���&���_L�i�� �R�p�W��n���O����+-���թ?S�dD:*�	k�^������ɯ<een�x �/!�����"8׎�Ù�%IPa8A̘84O��`���(��0��]|^��F����ĺ��� ��4��!.�`P��{��i��?��;�y�S�0�oե�=�������S�K1��S��:�x���ؚ�X+�k,�d�L�1@��S�L+��dG�:0J8Vh���'��(Ubd �$��@�yr��(�H4�q�|�5)��N�pfH��h�NV�+�x-���~i���i���cM�_RIn���^��rS�pt�0�C�M�v�N�cTH�9��z�(G�P!"��s���My��Z�_Q3y���R�Y�B�ь��Kv��}�s׷�<L�KM���q�R�!���QV��Qyθ^	Q���W'n!ۨВh`����+#_�l��Rk켲��':�i��$s���vu�q��OO��]����k!g?��(�.	0����1���N1,msP�X+v����2����c�o2/8 -*]��۶�Z*��m��<�P����QK�)	$��vN��b�U'�L�<��g�S�z1�B5B��������>���(�@K�y�|ڼ��e>%I4��y����2��U��M)% ����5�2�>g!d	�7�m���*�ǡ;\
�^��R�y���E
6�0��p4D�I ���ɑ$j���Hk߉��ɴ����8k��b�0[�}ggb��[�.aɞ[%+���XZnS��р�4X��c�+Y;6w�<T E�]L$r��5��MW��خ���<���p�
���K�	`S��e "���N*���rg�c�Zn<T����[�-L:���4������9s�=��֡�IA9�,��#�z٤����g�S�чA�@Euů��2|c/���(�?We��N�����.�̬dk��e�yע��5m�inFq�j#�^n؟eE��m�����Unn��I����m�u�;;�������Z�z	,�V�)6q���
n�!���BV5b�_����x�]gsF�W���E���+��R�ER�qa_��3}��֢�/F�wR���(�@����J;@@%E�2T]yh�X��l��9i�¼���$�f2W�u)J�4�!�
��W�X����r�S��v��4U;��{���]� ÕqG,`��e@��(�Z{�Ҭ����2/n�XM�mgo�k�H�,� k߻�H�]��leI������;�����F�km#VmW4C6��T���KUGZy&*;^�~�A������V�*6���x��	�XJ�.P곍�!�1�Y�`�~rTNӟ���}��D��3���/�황[������O��C�z&ϯ n����7N���FO���F��j�1�g�f�y�U�a��q,O�MQ!����٦0u�	K>��`�I0�'=�v|u-z4�B]oι���5�k��5��<�J��p��;J�W_�g�'�$��:�!6�2�`�������o�v\6 �	x>4[��5��'Kø~��|3��ӟ�WR�	��^yo�[����u���K�{MP��q�3�*��-���tQcm��^:2�̣H�AI���}
d���FF�3��P��������T%d6�@ �6J.�/��8Q3)�*u��2o�亂 ���I�6���E�
��օ:/g]q�p�az�$Rb���!�9�ѨKԂQ��X�+C���VS�e�g��a�
O�:�b���pp7��6�	����QI�m"�b(ײv]��S'D(��liL�������\(�T��8�,�(O֒��ғ%�s=;��cgә�#���^c(�I�}���K�[��Xz+��?j�uDvEZ�0��/�;��/|�d�:y!��.i��J<Ӿ@�)RQ_T�K~d����scN�q����B�D	����S<�ض~ '�O�;&����C?@��(3��2��3��NXO��5�N��U8Td�C��j�CT��>�FT ��c͕���"�Ju���`�?����ا���`*[��:4���.�PmJ��NN��,��r!;Au��'��4(���~�}����e�d{���²j��L��Y��k����yO���w6@*H9�?.\Uǆ2!�f2�������nü�j����xdLƋ��p���o�s��D�<��D$Te�Db�PeP��}��ץ�O�h�X�!҃�)uE1���6�D?�PΕP}!lp
*#Y����yy��,��d<I�,y��������M1ܹ:D��1gi���>�P���e���
D	VKr�8v���:�Aȕ��Zh�Ȗ�25�z�'B<7�}@��%o���i�&V�ģP�ܲ�F�߳�=}��u_��*
Й�p�c�������g�����r�݇K���D�mJC�쀗�ƋG�{�0����7��X�.SZ+Ƨ��0����D�L������'��#�̶��?r�ڢ��¬�u�K��%�i���ŗtYô@F�h���	i�OD�e�f�0{� ��.���ѱ���gI�U�x�r�]�]ja��?�/S3)(��b���P(�v���R��2��W$�x2��O�������Z����V�����)fU��a�t����7+��	8KE0�l�CAa�\�h��4��X����]oz��N;��B�%�!�wn��Q�L�g.4�3�dw#�G<�c�z�-� �ʠU��h�1��M\�B�<��=��iLo�b�kC�5硶��|YK.��β�L�L(]\6�p����;��+a�v��pAV��C��4�����:�@Qz;��<��d�'�;��<q�byq>�J�IH�7���-��v�(Ծ�B��u�:���v9щ�o�]q�,>:��o xC�� �0��:�[��-��K%҈���~0E��[��������$�q�S����%�zaJ(�/Y���r�</��t�:X���|��&�zo���3�<R��,���	te!��H�h��~�?3�I�v��W����%آNN�l�^��Vu8�zrR}�i�5�0��{��v*��z�r��g���uG��5�-js�)&���~,/L^YMaG�8��"�i���`�`.ջ�C�R1�-�B�xT(��^W�(_l�>-�I~T��W��~_x.O}�%i�C�M#�7���`Q�j����2U�,��g!�C��??�I'��2mI�<z��+U^�/��ɪ��_����Es }�$aǆ��V��爆���co:���2_����N��������z�%юw!՛}��>λJ����6��N������n�94xP2z��`4�9��>m�Ndx�׷/�='��9�nH:�ڐ���u�#��uͽ����.辰o|V�Z5�p��]���T��ٞ\��M���(^>O�&:��/�����}�v���E�B���!= G3'�B��ݺ#���ІI�77�_;��w�!�n=̪p��|2Zb%�4��9Lܚ�X����}֏�C��}���w�D��� {�	Ӆ�G=oqr����"��h�e����f?Q�@c/*�-5F��v�[q�<���vb�O�',����D��Aa�#Y�Y|"k��d?�B�XA�:t�w��x�"�!���.���W�O2 �x�Ui�n{�pjl[�N�M�`4 �,.1���{=n-pI�5D���D0"˶�V�0����h�R"����=;m�q�-�S0���^��Y��gI��V^�Ԧ����1��$�0�%�6�1s�\�s��`��p����_v��3_�����j�ǎ�y�N<x��q5*�N;�>���Y"$/T��?�D ��;�k	���ÄζCz޼��X����
>C�.��~�4���^W�;����],�`��l���5 ���̈���N����
�U��"��b|��C#)���<:�l'KZX~v��]�	���p<�<ԝaO�u�̥ )s�>I0xG���.���Q����%��E!�|�?���$�B���U��;�5}�����E(z��.�SFMY�zaU'	%Ǚa���p��r�[�=5�e)e%٨�s<(Ӻ����y���$`<��"�#e�7&'&<6|d��o@l`a��n���W�i�ٟ�
�<5V�!��*Ms��@)������A�sp���:2�̋!����*�I{��ȇ֨�{����c�RK^��V�	L�!QŅ��S{����"6�Y�5(��p���ʌ�Ɨ�|�t��J'�zNLύ,��a��_���l��Qّ��+�ޗ� UGD�~a�#��'���o�_�Lv���r��_�/���� �\2��R�)�nC���ąO�.�Q��o��Y���&V,���MGJX0KB�8�{x����4�f�Ʌ.���\��Dc�.��D�x�t�ڂ�.2a]~r�?MN�ՄW\�]�˓H�4��P��Hi�_R��\�pc� =V�8�Dk4C�i��`��.\ɟ�4�o��$�nm���.��#b�9`h`�6�_��&r��щ:�=�$s�=.�/��ۊr��6Ul$L�-y�
�j�d���:�B����#-�Ak],�\-��XMG�i��i2�9��S�I'�i(��o����i�Ĭ]���_����[�$�__6��֯L�t��!���@w�C�?e���}�뙝(���@�(�-�eI�A������QU�P�p���_(Y(V�����ϠB3}>_}���I((�iu-)��P.p�5�Hw6� ��g8W^�U�TeE$Wf��܌F�I�/�߶��ϕ��wWtܥ�������vj�{��̮s*4�x*;�ݖ�1NA�E�z�Hc��,�0l�`>�y���#�-wq���z�6��1��$
>�qп`V���8ao�a�1�qJ���PGɽC��:}J-(��h��_�~ɡB�	VӐ�껍�]�niC���ּ�.�!ڋTӚgĝ�r!0#�v���M2Y�<z�7����EnK�6��wk{A������h�t޲q����F�|Q�`k�� �=k����V��2j��tzʉr�n�j�i�������;V�q~)��F���
�!~OE�[b�L��G�0g��=܃��X�j�mӤ �cڍ3��=��p���\~Y\[?E��٩n�$���L>�C2ȍy��	Z}�)�?���=չ���踒f3��,��]j�s��$���P��!��p" m�z���1��Nk|�i�uẫ۶R�'GWF���h��%E`��+p��h%1*9 ���˛`D��@P�����kp1r�]mw���N�mfJ�+�&C����}_�������Z���ڊ[�uн-��l���7� Q�33=��ڵ��U�� �����M�����BZ*T��I�v��Q%�&���
X�������yژ<��玍{�S��s����C2�E��D��s���2x��aD,�*�Ws1��;�*n?ǳ��S6��1�o���Fkλ7�b3��?�{�Y����Js�������i��E���i��+(��l��	�5�ry��P1R>�z�}�������,��٨4�8 ��=9�2���Y
�Y�m|���4��h�5��ҟ�q�nk������R~ �* �#βd�f�/��2&gʊai����V���V����X���PO�<Y�8���	^�����H�UD1�b���n��$�c���E�g�;iRy꜁��5mb�	v�}lpW@>p:��=�:�%��.�ydĢ;�y6�)Ђ6�zz��U3I,�wg�@����a� $��+����1�ih�.p��w�WDG+���x!Sh"���t�=�M	,d�^��,�J;+9�bF�x_���%� &$f$��W�&ĒeO�%?Jg�Cw�\��-e��ڴP���.κ�,��ʙENiS�p�� 3�P�圔�
K���{��4��"%lpt�rU�*���B�)��~X�,���+,���m�ý���b\�!_'7�7��M�D��M��Uu�nHt.�Irp)�{�E��N���aT���N{h��X�u^c�i��r��(�=��da&�n#�I:Iūx�6�9���KT��ݒ���ocJ_�U.�o^�A��Ycg�߭V�/��ߐ�hm O���\�ٕhd�N��T��y���xׂ��*�ُ	�KF�#�8ߗj;=��`o�B���"�+u�X�\�atYKEp+�������1	�{�S�^��5�\��g�-v�����U�=��#�;
f��##8�Ss����|F���O8�rmxڟ(f�I݅��� �S����>]��?���_����ƠI���]��G"{�D�G
n�(�R���E����%/�T�j""q��<��M��0`��g��D�l�I"�V4�r�)R��,���d�M*0��o}�Cr\Hb8l����(Sܒ���m�=G�zy�F,_��q�p��Ob8��)�-� �9��x��Y��4W�̿v����!B�#f��5'� ~7�xix0����|�opU��!�pj#;U�!�kV�\ �:V[g�_��ep��
�K��M u+��п�^���l0�hW�돌�1�ȇ�
���=K�B1�$��\̐�ȣ��%�n]+V��;�I��u~�D+�i=wK�)*#~6��&ݾh��%�|�cDn�L��M��$���:8G���<��`�,$��G��\����{�O���Sib�n���^����B E�1�A�K|�s�@�FekC�;K�,M.h����F�7) �'N0�6,X�h;eF�̂���� �Ɣ{�/'J�]��yڨa-��� -�WS��_UQ��՝����h$�k���L�;C�=�7�>CH�� &!h�q�&�kcFZm��g�r79�%��͜�w�׆��b\�����n�^�����5/'y�r����u���S"ˬ2x��m��ٝ;�DqA;x����T��l��-Cr��D�8%�����镴���vj�5�t�S�XSǴ���̺��[�n�m��3U�c>��N0��~Ψ2m�zjmcj�jV�@����`)�sO#4�qs]Qv�u��#��W��������͢ܮ'��z��sş�auRР<an��.2g�F�����~gW�:-�h�TJ�~ҙӴ&�N��hF����ND�]S�z�m���֬����E�5�5׮�uV�Ͻ��H{��
��������`�I�m���p��\�PzP���,���80Sj̐{���i9�q�0���Dyjٓf&��R�ofA��ͣn�a��r0���\�����Ԇ��g��o�%���N{��d{(���D��I'��l�������R�W�v���|��F(F˫h�y���9��F�V�1�I��,�R ����B�y2 ��#��f�2���y��5ڍ��l��V�/u��&�YJ�*ro���N�#å�ג�ڎ��mW���AO�"�;��`ģE$<m�d����П�>�/��d��\B�0`���y�E��CI�ߙ.Ɋ�JF	�?pp��������2<č9�"�u��3�d��_lH�xX���F�	���=�|B ��=�u�.�U�iȊ�o�V@��I��x6�(��}�G�әD�c>g`AS&ܘ@vT����u��l���E��L�E��@�]�Vl+.��R����U�
^#(�A�8��g���^U&{y��ܿ%�M��F
kt�����_����Bu@v�P2��փ^i��B�{��������A���5Y�F��aC��!Z���j�iR�-����V4b�9E��-���q��Z�p�K�8�b����^��!&6c=@��7���U�[�S�ٲ��<M��&b׶<7�5�[5�T����$'8o�=O4����bMX���q*���>��r�t��]i���!]�u5��b��ׇd&)�
`g�q��+�2����x����C�
�<�q?�K�A�#�_yR�\��\��������a�k�n;�:�B*�E&3F���y�^����cu8�X��[�����z���������~At����xS��]��n�)�"�
�y�Sگ�w+0�������t��;��l�%�vA��ܣP%���@��1�:EXж��m�Y���$t��a�)*�������r���1�r��vdh`jW�Mm�ա�# L�c	tO}T>t
}�r��c �S�(b�
V=����B<�j�e۳��3���~�&�;�-Y%�wH����|m��Z��[.�sin��c��3��j[P����k��Z+�g�M�Y��ο����ѵ�F%��
��~{>Xm&�঳¨
5r+ALo�>x��?\Lɗ��~(�D{VoЌF�N��5�m�dJ6Vj,�O7̦ХC�J�vR$ᷮ�T���[>���QR$tA���Rjz;�Zz���p5�o����X�b�����<����O�����r����B�,��3<.��9/b��P~=8�?�K�o�	{+����fA�9�"ܐEx�|�vA��)����+2����aF���č\�����2D�T����z�X��e#�$zRm.�!?�o��l�������w.�X�2#ʹx����~o��*���+��R��55����`&�C�-��2wny)�*����r qg���?9��d��|��J�/p��QF�仯�w=`�4<(�a���u�*��2x �wh��-t��:~ܟ�Y�D�<����"ۙ:�m������Iv�
�(��0)��[���g�@A�	��h����x��`���6Ӆ%�i��X��9��a^>!�芪8���}��%�����=�רlr�)��б�|�L�"�H��t|A��N�z�|��Bw#��岯�/�N�{ؾ�����H^|!f�C��K���|�<�d���E�J���7]�,ZE^�Rtؒ�}���,��Lq߶"nd�w�s�Y>���M'�G�PIm�w��3+��dϻ����gFCtIӪ�	8���(tD!�K��38%��?E��3�W$K�[�ӫժ���m�l��ou�6���2�|N��]��)a/��?/����}��8�a�� �3�+_���?B��:Z�S�_ �<=���6A��o|�gF��f��X4�l�\����}� ����2T.{x�67�0�6M�{��zհ�s}\�A� &�Z�l�f�yBI�v%H��1�*�*	��P���ߠlڽ7=��tu�0f�|q3�^}
��QJ g<;~dGk"�����p���w�BB�M2K�[���7��o�؋��8X?+R:��N%���N���?;�	�"��]N`�ph�/����:���iе�z tL	��U�	r%��t'0C� ��sP����������E��3�H�7�r\ �.]���\�<_4��V�[������zFP1���'���Đ�3ʤ˃�
$��x����y���H�=�2��m��W�A�5��J��A;Ê�ڻ�?.�>R*_��_L�P���K!~�2��hQ�}8H�<$������q�u�F���@�����U��6�̩��;L�$H�Y�*���x�/�ܒa��e�h�XO@U����qg)yUm��wSY�)ՉLnL`����S�ZBor��E�͊B��V9���3^b� P��}��}eOZv��|�Ŀ҄æ���+{9]��J#��Փ�* ?�o���5�w�U7��/�D}�TkE��9X���Cո��lN�߆Bt�jk�L4�n�>+��kY�L�6��Z��E���<C����Gn��ނaZVҩB���_���>�������c��R�c"��x��͌���V���d�0Ԟƶ누�Ş���n͘� ��8�{��C�T����~��~��}��淿�<v�A��c��J���F+��<?0e �͹�R�
�E/F��
�+����=��7es��#���\��L��^[����+�GykH[�wBY�!��璨`��s�:
ҶI�A��c��8:j�y�>�U�������M-��LU��yH|"|`�0���ߟ{����z���V�� ��I+�0���e,���g3M����ܰj�����3[y}�^��{�	_q�fbi�'X���t�׻SA
c O��'��Sf8�=x�t�_|v���7)@�ޠ�8���
�I�U����38*�yxb��Ji��kU��-b������!��ճ��3�0����dkY�:��xR�!�4���]-�3���L�-X��y���)���T2W!�-	շ=�� ���K�w��!�D����;�^j�ޒ�s����D1e?c"��,�C�+��{���e����s�㐜�T;<!C����}���Sw6���k*2TX�2�=,t�Q�x�U�|@��T����.�f�D`mP7ͳ�i6�$�� �ܾ��Sra�\�u�LZ2�t�D�rX/Q����W[A��~?]�m��4�޲��y�.+���l��_uXP�A��$���� ���Ҿ�`���V��&v!ݑqM����#,i�4�
bϦӭ�c�,�H{�EXHd�<��T���.D�j�6��ޓ9Z[��Ƈ�TW��f�v���Դk�@S���u/.3��[Uj���C�/�)`O��;�Gp��c�9�[z�KIX�]�oV���>�PM�z��C�	��8�=��3$c5��LIf�yP�Z�S���ˋ^�+�Y�h�����:�;%��Q*����:��'�c�41X?�5Xw�ב�$P�Vk����dW����j�J:�7��CY꾖\n���P��ȅ�� N{�͉��H�qz�ZK�#c�f��i+���*h�Gci�(�l����/�h��nm�(������-
�u�Cu�����-��S.�G��9$o�o�+��G��ʓ�6(R�#��$��о�% 6��v6��A0ܚoV�5tF�q��1��)��b)�@�s}NS`c^z4�HÂ�*�j�����E]�S
7M1����N�)����� �7��N����4�V�9�Tp,d�'SSUФ�C}S���Y]�9�\߉�����/8ڞD|4-EN2@R�9&�0�c��^Ǟ�ࢰ��7a�|�_����Jw��� dr~��(<�k� >����}U������p�)!.�ݫwU� �gH[�aqZG(�V���J]2 �Z|viߤS����D�FR��x���NWI`٭	+����v��:Qt��E�Y��<ua�{��~ѳ�O�L�ߧ��Uvg���}�~��voR"7ÅD�V�����d�c	��h������`���)Q���c�l�K��"�f[�7�v�(N|U)�F��d��F@
?�|�bbȪ��l�{W���P�v��W�d�4P��6�-�%g�$r����-|��|C�E@��ik��q�󮡩�q���-Wk��N�����IL4We����L�.�]t��bW`����=Iٵח#�&'t�����
��G>��/�7Ӥ�T~�6��jy\�6\&m}��Wŏn�b��8Ik�	rY�&�AO�$w�2Ώ�3��I�Es�?M�z[CH��w�{��^-��$�wN ��Bb[i��;s�|��f ,���d��G�ӎ��EC����=jӶ2��Bdq� �Au7�|rn- ����(�ݧ �N��鸑� �+}=|�O�n�S��]7k��ȳ��&�˂"Y�ſ&�Lq,V���h�� ����<�L9I�n�.QL?�8 ub}3��G�?�댊@Kk��Z4h( ��|� ������>�t[��O<61�ɹ��<�	��mDj-�/���H����ߩ�<e����T���;_�h
�	
�А�4��Xw����r�'��!)�f��q���Lբ<@�>����qH�

�]l���0�^h�r
�º X DU^t�ω:�l[!KG�S�ڑ������|U�Y���|M���d6!�lQ��l��j>����Q4��ñ(pngJ��$�Eږ7��A�g�/���`�����(Kq� ��� �{�Q.��#4��� �f�lfg\�N��O�B<�S�B��Dn����JbKYf�4��BwF8���ﳇ��l�
{�8i�9��V���cC�� \{]#k. C�
r�LtQF��@�4�o��N�]n#Ǧ�.0���џ�����O�������^�o�U:�38Le��خ��TN���S}�f������2��J��ҏ���S���"�@�@�4���9�Zs��Ow�]���w'�K{�C����@xc�I
M_Ӕ	e��?��R��3}�=��u��D��D[�,����2�l"c���t���i�e6b^۾,P$7��=�]���Z>�P��d$D��Y	;� ��nP߬7��q�BƳ� ��Z���:@C�q;�尚�޽�x
G�,��ڣ�CB�<&���?�W̸�������u�gG�-��y<�U,�����ʦX-ʣ�ĲD9�-��5c�GJ}�����������fU0�{е���iœ�����4��Ô���Jy[�i�Ԗ?�����y1�S�}{�	��e����u��x����[�h�˳[�%�#
�1��眗������!Qr9�ȹYp����%�G:&2W��+itrZ`Qi�B�D��'D�D>2��[����;��3����؎6� +Mf\�T��'���>���>��F�~�;6����C�^�;}5���þ����R��lM�Q�ڭ�� �I�1d�V�%��l˶ &��������j��i�ob]Su�g�Ӵ�E�WG��5 �J�L������m�>T?�7�w>MQ'��9���,A��3i�s��b��n��9&�}��H1���e�:�������%��#��S� ��3�@#�)��،nhXI�ȝ���#?�Ő�Sj{+�A�W��:���Z~��̲G����i8�K��W���t��r�8Z5��4�C��(���@Ͼ	�Ϡ�Q�bv϶ɯ�2�<g|�k�,¢� �I]R���
�#+�C�y���>�(Fh|��B?�gk{��j��j�݅\ٹ���0���]��ݷǱ�U�d)��H|�T�+W�LJ)W,H�N�Y�k�E/�)�)"qU-0�0�@�y�6؂�1܈�������УW�h�aX<`$ Q��(���&��ީt�4?o#���/6t��R"u5��t��F������"�()��1Q�u\���`�/�K��K!?ą�j���g��_�?Ex҃F�}��O���D�K�ģ���iH�*7��c�@w�v�	�?�I4�o��q��iH�]M5�6�QP@�l}�[o?h!�"��}L����q����X�V�����O�����[�|����쬗XS�[�1��~��L������#�e��jՠ�O�����~9��osw;�=�|7*��IN��GU��l��C��u����1����f�����-Z)b�h��(�T1��f��)���t�%�L���!|6���l/�y&����^x�/0d
�`�[���RBBev1D:	���æt�1����E���� �4�#0L�5K����AH�T��"�B�H���OfIͼ�kq�<�p�P��>��*!8�4ۖ�~o�s�{�C ���1��}E��P�\�=��`�hM��0=�q�/`�<�է@����9�)F��O�s��7=?��n�{N������s�/�s.�b�f����s��vӏ�2�^�:�	�>��o�������_���G�j���mWi������!�	��Z�l����D�B'�j!��⋿g�i�x���;e� �Pw p����(�1���сn���%\Gǽ�e����͵�J�T6���=�A`�uq�������sV���z�f�TS8�ƞo�����TH��2Yz_r栯�i�ɬ%fW�B@�n���)t�8��s�:��
�;��$4�-�u�ϨOAع���VCJ�oue��~�V�Zj���/��{�KhXa`��j�,R��]A�x�-�D���2t�!��~�(�����AN�����I�o��W����Wf�IX�}2J+�����'�
��@�o���]:�i|帏*�/ýW4�3(���|�Fɱ��Ő3��`,�\B�O��gYW�k_�����j� �#���5�����/�-��UI{�
4�{O��z^΀���Ղ����zNl�!}S�Ɂ֤����$
V-���SB�e�Q*F���Ï�cn���G,�}{�÷�x�z��b���N��� ���1�BB����g���P�V�;��z��ݕk��:[�	�����L�����e�ѨpF_����=�#mzv6��S�H����ba�j)�����1 ��y�& �w���Қq�`��#;�Y�U�ځ��g����	?�R�ΰ��Ҝ*�����o�J�η%����d_urH�gS8A�4�;e�J��M��~<����׵b��d�.�fkc�=��P��jDj���a2��B�@6^c���K��J|<)�	�S�<Z|Y [���g>V��3�*z�:)O��$���<%�%+��ï�!����R%�pv��W}���+�Y�I���A�&,�s�s��7�3c@Ph�G\C~Y�������}��z�t��M�3��RH|܂S��oo'X��/�ˆ�r8��;Ӏ���z�f
%-���HfC�>hS
}k�� }��BR<�&-��9�|����lY�6A"w���%�y��ou2j/�o1%W�CK��:r��@	c:9��q�������W��B��f���S�Oԓj�]�[@�h?����\�@%�������e�H���Qp�A���A��	��b��Uo끔�8�kɜ��j�0���T����,Xv`�Ao���
UV5U2�R��&{��UB�~�R=��;����9����#�o=]�����g)� ���,[\�S.ivd�$;\u����uz�I�`G�j��؞�l�,�;�SG�Y1�5
�@sS~#�i~{�1�����1���ݤ�����f�n.��k]b�-f�Σ����l�(�|�TG�2.�); Lû������쓔L����'W�ʦ��<���9p��T�-��ؘ�P�v6xu�ظ�H��j��%��,�5��Ϛ�os4�SR-�	��+�h�":�g�c�Bl�0و4w��h��*HO7;IS]ę�¤0Pg���8���l�Y�Ek��s �����e�R���i���A�DH<����lS��E��(����+r�/Q+���@_I=\Q>׆�u�-W�$��,� �g�#c�����!�>�����z�]V[�}B�-ᘬC�5�}�Z_
�ُ@z�+vx���NO���2�^]\l�E���s1��^֪�pP�	�%f(��Y�4��S� A�{f�WԬ�ѐ�����7e��0EoY?8��_�hUՋ"����z��K�$�����ܲ�j'(�*��[h�1-q�����/�򹔓�%>�"��GJN6S�/�!���JCI[�*�K��&��嚔H���B�k�ڌ�N2�L�C_w�����̢H}~��X3����@�ۋi���.��t���\�)��_��X,c��|0������t�Ec��f��KM��͎�(3{���K�K{�wG@�n�1`�X��Zٸ�,��/���؄�y�������Fh.�P��$�M��FM�
R���r˭%���x��b�M��]�b�V߾M�Rud�ր��_`lTE�]�`��8dZ��e�^�LF�N�78�b9��Iq�0������4fp��?9M�(�BT��߿_'u	�A���bx�C_�Qlds}o�>D)F\��l�y%�~�od��<�y����xwwS��Bұ�Y�1��|u��Q$���K���k%z�Ӭ��m�����QpY�������25���<��m$����]��>^[��_�)�$�7�	9�
��S��t���,�ڗF�u��S��(#�d�O
��;��w����t���K4Z����^c~_�R�F�����Ȱ�!A��Q���Q�ȍ48��n�ox	�G��\f,-�[8��L�nh�|m�	��]7�c�}�]��q���L�v���8�-V������}Z�J�Ri���M�D���g0k�bG���D)��V���5z�l����aN�!��a|��;�	��C���^o�)��	k�df�5�?ƝR�E��B��r�i��QZRf�$���8�C�!6l�A��0���N:����`P��*<�fMN�3�p{5͗��NG>8�UlG�1:�T��w�?^g̳t�Y�ߺ��+�"G�X)��X�B��rJ���iD�T�ti�(��像�����^C�s�-�f�4�)9�] ����Һ���_^�'��ď���T�A1u��_C'&b�[f8��1k���eXi'�z�:W1;�։kh������4�,S�²
�̇:��v�5xVI����O������v����x?{��� =���>BB#��8�J.�UF�%b�0SLL������Z�}b�e��\U�Y@���M��:�=��{!��I�١����p.�'��O�u�K�!_p����k��CXHS��jd[�wf%�m�J��њ�/�>�ʚ��jF񍵊ǖk��a1���U�d���3+��BU��(�8YW^���x�8��Ptt���d�уa���-2vv��E�&��lßIC�qsۍ#k��cs�w�&e��B��0�X�9�gd���{j��0<3�+-(��DR�!�R3tc�
�8;[��߭�Gӡ����UP�<w�)8�[@.$�L����
��&/���w���%hv�N��Q�{&h7>�q�rb�.���*p����ј�A�C�@L|=��Ȗ���.l���+7h���m3�Вo2v��X��©Ģ+�o�����+{?�2��r�A�̊'�_�G��DZ	F�b:~�`2R�#@���g�]�0fnx������ZF[4Vi��U���V4�/Ҫ�#!�k���*��|�̨Q�S
���8P8�.w40�m��&�c$4k-ݮ:��!
����%�R�g�_U~B�|�#iyQrՄ�M�g�6�+=X2$ Ǣ��Ĩ���Zn=.\��#h4z����e�Fk)��BB;� �H\c��6m@����3p�I��}Q�G�n�^���Yv� `��?v��Fl t��1���{&t�k[�	�-�vѠ{�a�.,&@ԀT
$�e����\'�:r�P>6��M��E0������>ݯ���DY-P��-�BM�g���b5���?꿒!Kxrل�I݉�0�,td��i���� Y���ʁe۶�/��O��Qˑۉ�X�p�Zw�y�'}�fxy���&vf>_ >4�X����7�E���~�ϤjG���>���O%`�J}M}m��ͩ��5o�|��(���P����=�N��^���@��s������H�g�����)7]j��)"���6V��B�RQ��О��d�NQ�Y�K�pV�ӌ�]jU�/?�]��p`|F����z%,�Yb(D�P�$�VsF7�Pͭ֍���&�������e�3���r������R7��LK:� v
�����}���9�A!jh�'t���yQ��ف�[d�ݦ����$��夭H�#+KĀ.7�bwZcj�����He�m:A��&���3����@L��q�Y�adI('�}�Kg�~o"�]�iU�ʑ
�.o:��܏��z� ����8��&�Zc����ʺ��O��i��-��aR���j6�Z�媊q��x�Um;d�ȉ۹�Q�f?�?��P�YQ�h$,�:Iq�d=�?(
4��Ʒ�:OG�{���p�SxN��UaՊI^Tw=%YE*G��./dl��T�{gҏ�u��v:{��/�+а�߮��ަ$Z�]M�W��^��sYa%j��_����c��HD�l�6�%�ކ\p6�$����j�"�o�lS��6@b%o��横�i)��ޏ�yJjk>f�5�(	"KJ�Im(��##�^����d�4�0z*ȸS;�S>P�ܫ%_�O��j�_��un��#@���sxYN�e�.���$y�b-x����3U$�FO�G�������֙:X�|+ի�E(�D3�Z�Z+bts=������8�<ͯj�~�CC�׉�:������`ko3�g'B[z�q���b�,�d��S�ў�;�?�f��͠,�&4H�D����
��z�oP��<�^�Wɝ���?$|l-D�R�&�qj4�v���2Z�Y���iI�Y���{_�Ϫ ��+'ۼ��������m
LQ����'���1�����ڷf�(�+��Q�}p��o�!���y��WX��dZ-N��V�ˡ[�J`�7 Ʌ7)�C"�S�`g��©��i؃%��E�脥�w��eZPp~�+b���࠷#��V����Ċ�g�o�·�]'u�����G�21�vҤ�:��r��a�ɣ�"�>^"����T	��n�;1vQ�1B��̌`��XG�K{�O>O�b[�@U��e���ha	�8����Ζ���J��ߚ��ٵ;��5C5�B�v���h�_�S��:�繾�Ud���������7�r��������,8_?&c e�W�_Bf[����|�A}(��t'	����S�X�O�>E��|B��B6:"߮����<�\�=Xl)��5�x�0Yw��}��������̆��[\�mj���H�	\����C:)_N�MA(�Iߣ��z7�a���O������>���W��3}��GՀ|3RE�#�5�Q={c|���a3�O�&��3U�.kQј>��C�V��%H��8����¥bt��ooPR|�ŋy'��ܚ]�IV5y�Ѹ��e�<�4r1f7�m���B؜�����.F�(�I'�wT�k�UIf��"�����㿝+�����w1�}R&ZǋXv��"�@Sö�<���6"N���r��/��=��R�� �$�W6�Pŧ�-����F��d:��w�F�Kۭ[�Ё;"���j�5��a#�W���*��Ṿ�
s��IE������5�	տ;a�,��4���ܓ���F8��� � �@@�|�-������6|X����$�e�,`�@j�O�4�A��qVx�4���,�1ə�£DV���KB�h��p+X��XvKW���lC��b9 [�Az��lYTF`��kG]��,��QZ&�I�r��(��_Ou�����Ux����1�t��<���,w�ܤ�A�2oT><�[�m�L0�*'�r���1]�C9=R(-�֙k ��)KJ��k�l��[ D�(M�  BCL�����7�
����Vōd8͊���My!�&�wO҆���cuZ��2��
(�P�>Ы>�Jo���2#g�"���j������c��PTnf3k�{�=<�YL��m�S�2�D� vg�1�<e8���ި<J��q^ܹ�]�\�b����1��.�'�L"\#wat/I�<���{��g��W��U ���)���|k
ܓ����؛�p'�Uk=���KnKe�#;A�����O+B���DW����A8G�*" ��qhͻt.	�RzԈ�ư*��F� g�<W����|O!n-�D>��?�x�w�>c���d��ꕈ8��y��9��{J	�i_���?��� �|/�r�Ě��Q��[X���DE�J ͖�|�����	Ȁ�^W�� � �K���@��r
�?)Kɫ��q9-|�Q���}r|��:�����{Kq�ScJy�i�*�T���}�V�C�G��+;n�[+a%��H4��b��h`��?qP��{�8��u�ؓt�~�UOv�4��#�����`��-Jt�U��|��um�>�O�eE�����ҋ�Ռ�ÑT�=i�r..M��OE~�~�\"�d^�E�x��@|y~�i�Ϙz��o�{e����[#2C�(��z�T�?�)16)��D��+ y�
��d^���p��5�� �=��#�����N��2�-Ϥ3ͽA�.P،�KW��J�A�f)�}��	|��IU뜚Ӷp��0<���/�/��b:B�p1���y�v�'I("�FK�����B�)p<!B�Nf[�Ԝ�Wu�z�QmքZ�" ��+����Y���w�I0wH�}���w�9�Q�z-oT;�^���П��!@�<Yݙ�>�V_!)S��i[+Ү
���l�F�08S>F�(�c��m�;�K���0���@��+ev��,�#�a%t�fd���Y쨄����=���gLKqpQ���c�FL�Њ[:+�N�PbW�9�6��(��G�����{��I����mI% j,�ЈHh,�1�%��\JNl����ԼhX��%D���?Ja+�C��SC�2���R�y��2��`U0�������%�Վ��R���-!�~�GM��W���җ�Xt�~��~����0�7��67�a��AM<k�^k%�	W�\��L��y�z�#d2H�s!�Ϛ�\X���503z򹀲��y4��o��_�0ך�lzFJ��h�����!c����{4A֘�<sT���n7$X��fg�����,v�O0t�x��\�RɎ� iEAhōr(��/z��ϨoAp�rV�
��MJ�?b'��޻�aV��p>�\��*Fx��N����#w�ˠ<�<j[�I��Dy7��9�!w�8�W;�Q��w��O��n� EN�{�G�w��#���+��2��HOQ_�O AZ�O����ɺ�[D���ˉX�߸���o�ܺH	`��*����d0���?���(��_ΡU��� �(!�xJ�k�Ѝ����Ab~�+D,)%��gH��dݯ���]9��PB��	K�I��[�k	ĩ��Q�o��:=��fq>(����Q"�EL�L��*"@\�Ȭ�ވ*��=߃h���|(��c8>�n�x�P#�r{�6]��w�}\��fKv��
������;��fi��	K�h�:"��l� Kwܫi�u���k���7q��C�.troV(I�kvy�?����bD���;���2t�F�o���i2�Uׇ�.[��_�tP<)
����m8=d,E'F
9�2_z3<�T'	��=��i�)�3���c���sDWA�e��Q���gF�^�CN3�+6��:��o�Bμ����;~�}�+ݏ�x�Fn7Sa�k��;�x��/�Z[�}�>��>|ԾNi�d��w]B+�3��Ax�{L1�Ł�2_| ��B��������A�_�3	q�۪5��d�l�J����i�/���}��M1��ݡ����"'����O�yE�k�Ӣ�`����I�@%�й�r�������v�&�n7�>�Y�~���uF� 5��T��>���%m�]cypZ���U�cf�dx�%��KI��(ס�LI��N�<Y��G��jl�Z�m�/�a�F0��*yC�҇����o��)
"M���F��ZH�|x�m5��V�em�C���ol��`Ȯ�YѮq�@�,a�8p����`8D�M:
rߣ�=��������TB"�����M�����9�}����u�ʡ�HCz���~eH��a��>c|2`6~�dp]V0r���h �q_7xc����<��p��[_�Hn�h�vu��p���p�5���N���VS�\����2<P�uiU֢Y_��0��'W�^uN������U��Z$�|�����Tz�)�)S!
g��$
2+pϸ����S'LR/5<ic�����P=@ɮȩp�8?Z.ч�n3k�7 `�S�����"����� �o���"<�!�6�RsFc>�� W\��5i�݌�/b<s����(����]Hy��#��Ј�{�i��=5PS^ ���p�!܌'�C]��d���6�n����U&ߕ�����Z[Z Iޚ�퐵�7��
<��L�i�D�M��t��ɯIz�'�?�;[{��=jO0
.��ݼZ�ߧ1�2BP悜%f�9�&v���Y>}Ew:3����$f2��9�uH�<��`������� ;`��n�(dS�8�r�D8���B������}���,tē$�I���ٴ(���9�������A���.�HtT�VS��Q��T�&.���	�5������~V=��v�.�L`In��'�,3�T�EC�=|�P8._�{�<L��|*gEV�P�=��m��W��gU�*�8�I��4�:�'�t�q�����g;o��R���Ul�Z]�ؤu72�9QCE'c�fi'2G	�����@�JC� �4rD6�Ҟ��{R�V����FJVؤ�Wr�7�=.N��By�X��S8w堳 ���Yz�{$Q�4�u�ꧬ~v��	�cO����{�v,�"9�t��-&%���3LH%ŦGw�? ;}���D�X��F�_!���٢�-N�$���P��,ŀ��&����S�T�wWS��Ъeȭ�x�*+�V�h���*i�KӜ?�ڄ�����G����%���	�3HÂ5��q[7jLb'!'�[�y���Z�$�.	������]�7���O�2NO����ꘂ��RL5z~�ab����XK����Y$���k���w��;��&��W����k��wj�X��������,vo��c�u�'zD�.� ���������������ϫ4+?[���T��L�2!
!�BHqI��IR+7H R%�c�Ԃ���^��z�6�]�̺��l�{��ي^��m����u7Pu��MMu:�q���ʟѷ���N��P�p`�=+N���:
ML��")�&�p]M�������.V�h%�)�#����=s4����J��h�Oh6�]�(�a+���T-��d	Lis{ѷ�Q5B&��	��㋗���)�����o��h�^wg��"&��S��h�I�����b��Ӌ. R�!������Z��;L?�Ee�����m*�)�R��ӱ��1i_����Yc��7��3(��$3�e������c�|֌���bhdl���7���{�����No�B��8�5�di~�� �ebRPq��czwŒϗ ڣj�H�t_Bc(�M����$�C8�
k�aY��2�rɑ��	��9�{�}����
��>���Ƌ���K����X-�k�@;!p�m��}*cRTȴQ�u�Վi�M��/��v���]��|@�=)�.���U�񄚺>-C =�j�5+�}�f��_L�٭#�-�c������O���x~)�lm��#�0y��5�>�#��x�X����ba�Z)hXnA"E���&�� ���;�範�ø�}�w��]�C�{�d����Е��oxl�w��>}��B����>��O�ts�����L��˄/+��tr�|��!��DWX��9*{�Iz�Wf}z~�u�[�D�y�Jt\IP���|�S'(kyߊC�����?���vD�Þ�h%�����_A�V���!�M���^k��o�(�)����}0'�?t� W�� ��[�\�$u-R�o�B��r����>5Z����6��ߝ�>v�U*��N�G��cX>�t�K�߆��<�-@~l	9|���l6o�Z$z��[�!{7@є,�	¥�kw�����\��>�6����H�^��Fڰ5 ����� ����MI2�)���6>�,�c�I2d;`�O���A\R��N�y%n�g*�N+�t��Y�㹯5H�?�-�H�� ��OC$�|T*&�nye�"\y�牀X��85Y3������>��S��V*�2���$�_�����wp��V2��i��<9䱵}X�H0qb��×����8�Fe�����
O4�e��T6=t�!��Q�$����]8��P/i���-O������ˡ�U���b���] �x�����	ޮ��1Ҳ��6����>dSv+lP�Ìj$�Vs� U�ڲyˤ@��,'�����c~��8�sY|@��5N���`�G^�*Q޹�٢9AVk
�!�W�D7����HK�g����f4R�,��HUG��΄��

'����S���]T��.S�G&*��־�{��L���O�=��=H��Q�:/�= C��g=r�eԑ.k��Զ�w�M�����aQ���t��"�gY��¨�s.t� n����{qA���Ḩ�+^��V�ҹT`���P�ץ�gG��9��ź������V�Oŗ��X�A����4���)>���>���1Д�|�m�r��ņ85Q��ҬZm���q1��P?���7��EX��:6��	i=�Mh�<MM/�e4�5�]M�{2�9�!�����)��0�n��d����֋ۿ��}�m~�8��|��{��A�������[L�3��J�[S^F��.13�ݔ�{�t�i.!˛�h�)ğ4�e��_G�)�;zv�%ʮ��$3���O��9�!W]�u��o��A�z���ÒXq�5\�+@�h�E���O�]�}�![��^�`���&���*UB߉�\&ZG[�1�Lp4[R�q�3t��v�%�`����M��#�aa����	�t6ʩx��=l��Π���Cˣ4IѴ�]��L��m:�U�&�NbNp����G�XWTw���e�խH��c>�����<��Z�t~H Ũi>�*4.��ȑ$j���Y�i�YZ�
���G�Lsг]�(Z���~RX��[��g�
�dB8��%�-��t ��lϴf�S���(#���ۀq@��pC�
�����(�JM|`�:=��o�КC�������+X�+�����o�3�_�ď7n��L�?��k����45͚$�ܝ��P0�G���d�EU/Z�W^�4jtM��xW�1���� �-]�Pź�y<O�>nd�xt�R\����w�d�/U�1h3�b�+�@���<3dh�� :���h����[��y�� ~ ޚ��Q��N�����ӌ��˦� G��۱�MF���l�Ms��h�W����k{#A��2�OC���.�U�[Q�`O��uh�S���
YXz�&AGc���1�О�j���l��H�����mNy��[k��B�
��
��g=��f�G�����CX<���|��6���`�C9	+�q3���1�X�>�;%��.|̕1�����c9HW�ǆ�p=�e��p
����B����s���Xfz�>a	f��7o�+P}�M�|�QNj�n*��h�Ey�ϱ2�b��$�f���r������8 �spV��2��z�cv�oc��%ס����?���$��gH�\�^8��03��J ,V8[���k��~D�K�l�>=�{��3^q	r�Y_�;/ c={F$��:*��}�!,MC<'u�	���*�\5�!�l�T�c�5�"F�oe�Pj��/k�o��.g�1��8��X�v�e��Mdi®u4��[��ABeE�t�r���u:���_yQ~}�C`��
;7��{oo�!�5=��o1P�����@BCs�P�U�X��2�?��:}ØŖ�;9 xH[��m_�l
W��UVS��$F8���(���.{ž�}M���&:+m�A�V���S:�-g�����m��e�c��*����1�������R�	����~������Z�����]�P*y�D���]&�3GN���u�����J8�(#���O�.�D�8��jf�\!��+l�d���}(2�l�rՄo��'�
!�S���a �tau(��{Y���e��p]=�]*���!�����_���I�~���&ΛF��$��2DA�d(��,J��f��d�V��֫(��+���W��)���-㦃�5�
,�A7JaKl�����Դ[�GU�&&��k�k|�Q�jw9�
t!�Dq�:��N�Z�ZL^���tH<ɼ�vYS=���A��ѷ͘���gQ[�o�Ղ�LB����X��a�cn��PӍ�a4gh&d/E�^�4�-/����#�@[��:k��y���h&�O�3�7�Q٫�ǉ4$�aNaHX�bA�&�t����	����e+?��v����_>�y+�]�g�&l�^=��T�r"�MbX��0�N�i
������W�y���	��k�S�K��6��y^X� ȵS�<�#h�+����n���1HZ���3v�����%(^��!�@����>9:db|�X������r��S�\0�6��32s�z�S�;gQ����fJ���˫8��C�V�m�,�>�ϛei���JQԓ%'��f�ʲ/�䗦Uee����	4�����YH�(�'Ѡ-?j}���Po˅�s��њ����:�^���nA���zM�*[���?��yꉁ⯦�F�
�j�0~g3������ҿ������!�7�8w����W��-B$ Q��{pfs.Rf�%���:3�ߍ�Htje�v%�V��n�9^c.~�7��<�L�==��JF3z�Ux-�ߟ��cŊ����[�a1�l�t
����e�
x��V������U�^r�@h7ߊ̚H����x��'EG�Bo�(E-y�Æ]� �"�X���ۂz0S�+�0�����s��_ms�d�S�U���ۙ\��k�q�D�g�I�)J�wT]��t�-�G�Z��c����n�S�y�z=��O1��/��� ��ǟJGmўH��ȿaW�o�맘�f�3<�5���[�NTm�r�������	F�������
Q̳�᥊������xK�s����frz�D�p.; $�Ͽ	�$o:U�6g��������NNK�l}����^\�*n���a��5���r��J}#&�CTr��V��"�\ڴ�1n�]t���We'��z�hb-v�_-I&E���`Tt�e�p4��Ғ�͝������p�Cڔ�2���h�f��ҰŘ�f�"��)�ĸіL���<�瑵g�@k�=��uK��R���*���+�K�+j'GyM���5S���RQ`r�������������`:��ߩ���u/�=� �gjj�W�\���� ar��>K��{��Ռ�nmm��A�ׇ'Ƽ��K���#�jS������i���o/��!tb��LE����"�G�i�#���E?9�P����X=,e-���ശ�>1��.�J":Ȑi�	�v>���?��� R��%%y�vz��$�[�G�N��as��y���g/��EކMY|�un�g(��@�414��u�$n\�hT?��#/U4¾J��@k���.��wWiU����wW�18����x�0Z�q@��H�����mt*z$4�ۛ�24��(�$���d�AI*��Q��������q0|��ܕ5�S�1�cF^�r����ģ^��m���LI����U����b�\�a@��t����)���	�rE��F#����U���9�V�/$W��΅
�_�G&�������j&�ث����Ie���#H�Q���N��M`ƥ.��}���J�>�NZ_�|0�2H�;�Ξ��������A��������fO�n�J��P���i�Wvb9���/a}R����y;��i*q��i��J���Ù,��˸��,�nw�mӄ��fǠ#�ʅ��W0e=���>�^�g��+g�m�9�c:��.��Y 9��
(9z�L��fp��_o?
�eK۵+*/�%-�C�~)ǚ�V5_���q����{���5p�r�[�	�g���4��ߗ!&�۠��Dt#�\eP�,J_�F��@Ma�t�����'L�[ p�jU���84�E�\� ���N�I1�?�,Ϻ�H����6Se��[c��o��&D��a���N['�i��@[���b�����֌�FpR��1I�E뾦�_�����n�1HG !�W���/���hjgܵ�E�o�X�6���V�Wq.p��	���,� ^5�me��ٸk�j��d�+�>R�آclKRe���c�$B��N&Ǌ�6U|�/�1��G��`� �E��*j�rEl:Y�m#����z��T�ҙޔ��LS���QR+�v���E7C�wS�WS��)��b��&�� F	���4��8�iȸ�i҅dxը���L��w}H����j��J"��NNr�H����/��h�x�p��m;V�����(W��qsfsI�#�m��:��&��1J%���D>綅�7��^���N�y�ر�thm�����y v���Y����#y�=�?����YH݁#��
ٻc�_^�+�Gp#��#(��Or;��Y�&AǗ�R���|7��,ÌIY�Ɓ��PAu�Ӳi@�Re\׷�7����c0�k�Z^x�9p��E��贎�6�!���b�=P�۝`Pޟ�i�ӡ����g;���Ax$�����&�=�h%����[S�A�%��`E'�K�%O�Sq�8#ff�'�2SMX����'��q��E�N�Z�%�朗o�:�sIQ�����E���Z�������0��'�z!��ꄾ'Q�v� �xgo1߁�0V�v��������r��n�^{��@�$#��|Y&�� ��TU�v� ��"���I���J��7��C�4�D�=dw�b?�8N�~!
��f�id ��� >�.S�7�!,B�j�{vUoK��t��Q��p!��h���8Q+`����/��a�A�u���F}�X>��$�_'c�	�ܼ��,��=�Ue�w[����gvmY$˄��V�P/2B����g�������V=�/W��#>+XL���;N+ca4֏���{-43�]$�3��j�ݞ�=@ߋPQc�lmSH�f3JWD���s!p$z���?�U]��"��k	���R����FܳlJ�g7�k'��E����SB��+R��3�$5�k���s����Kd���[0�N�]��圁M�*�B���A�����Ex^�I��)*J�Z�bZL� �-����3��e\�3#�����#����&��ۜ��'s
�
�ǈ�}#}x�'d��<X�Q!��4?
�
��H�-���}�������}�`0��G�֬�(��Y���i�H�p��|�Y� #�ҍ��wķ�pV���>�h�֍=*⡇�è7�2)�<���t���*�!��չτ�5�.d�SB���FGe@&����� Rm����Έ��~�r�0��r��w���9<d�83"��.����	1�Y=F�д,!q=�.��|�-�X�vJ�)��Z:���k�SyI�&�[#H=s��2�zl��Q��r�-YRxH�B	Ɇ:bV?R��}��t"R]�ءR�T�-)/g�%t�z���N.�"F��%P٢I�޷x�M0�wG�H��-A^9�i��V����e�p���V�ҭ�rviʶMx?�[���/�B��������'�(��pM5R���>E�P�ߡ6�CJ�z�&婊���l?�������
�h�93ƙ�R���M�����X�1H�LP�a����P��G�� J�\������qXdWL4A~<}�la&0D�����m#�f+�ڲ+5��:�0�������w�d�rk�IOq �^�(�7��=MB@Ǆk�/�B-�Ʒ3�b�#��ێ����xK%;�N\4m\bF�`�n2�<�1�.��I W���wĽ�� ��Ci�yS
�Y}W������|g&�ZТ�,h�W���i{���fuk�_��d�в�[��Z6-j$���'},+R�
3_�ʪ�Jt�0Sa����oͩO68�_�<tef>�<��:�g�$�?�s��e���mc@ch��I�����S�/:��t��Di��B7&�:��[��e�,��=��_9HL�.V�O�
y���,���[�0��J�D�P({�-<���T����]w��D�,����O�H2i��?��T�+��P�ߩ���2�!���;�1�7�����nV=��-����o� 8���+Wjι��	�}I���>��n��8)�1.E,q���mbNK�ݣ/��E&�>"[�f��[�!RIꔎ���B]�"WÉ(Y�q'J�˜��CI:�B�b�r_\P���]�p<�6�Yp=�l�(�m]�e��^��[��Ϥ�(B�Ė-�rc��d?�bZ�Ba�XUub0��+r�5��8��<�9��$�h�K���+%��9@V����+k�W�&8�x�0�v�[�����G7��i<�4�����Щ7/ ����&�Yl���PtEЊr�{n��gW�Q?��-�C�ӒFq�w�b��~��n�3y�����<��J������8`7͆ݛ[|�퓺�簨�-�[��֒�ܡ��2�i�]�k#T1~���	 1(�r��#��&Z���ԗ+�l��a� �L$,<|�S�?Ln�Fo,�qh�[��9��lU"BIƀ�5�jdL2�A��َ�{��m�E��>�5M�p�=^u[���!S�L3r�C!)���v�n��k�%���\ ��B%v ���99zzi����0c������R���!0k��̈́�ƹ� ���MS�;���X ���C*l\w�r���m(v�@���S��w\��bk
��l�X̾`^��@�$+�0r���������?��� �5*��y�h�� �ld'�*wm�$6���%A�PE�>LC�5���\E%�u���UW�2Kٴ�<�y�gB%�N&�
���--��+����B*�����C�{L?9�_t���v�{����Y8�([>��@#۹��o-rs�g��C�a;B�у����Ꮼ�C�� ���@f����g�-�#��$ �'��ݥC�h��������t�`(Q�{������^"�I�wi����<�%�NY��/p�gM��Zm�}*c��#��t�t#�\Bƻ\�xMz[$D�{�@+-��~�W��D�D�$�-��4+l�s  ���[��5��ݿ��͏h�{"5��' �,\	�)�Ԁ��4j/���0�p�_mE0�S4n["ѱ~��0�Yʡ�j��S�!	���Ai>>�X5����@�H@�e3�#���=�
0' �L�̚/"���҇2��mN�z��)�iؿ��J�������.M�:�Ŗ�lڣ�Q��ݾH!��:�3mb�G������-���D�1��cɏ���g22v}�H0�<	3ȏ��ѷb����s�!�(m)���Y�����b�ɍ�ԋ�y�d�f2G�k�J��̅EB����
2,~��X�Dp�nOs��	����<�vX�g&��DK�KL��>�WZ��'���=�U��ԑ���ᑨ'x�_�l����c �D���=��~����ޤDFr"YQ�$Y�zv���n���.���F�U��>��;���ce�ҧ���p�W�W����<.���X<���kd�t�d�$�IA�.E҉(w��ڐ���Қ��k�"�{�����R���Z��g^g3 (��>�h��AɏS2*�!�E��[�|��w�͵c�$e��ڷ�!&��i����S2��p�I�b�h����02�0@�N�67�ڧ
�n�Q�C������1��v{���X����@��.k��B�/?��s�2���&��[��]�������*��.E��(���T�S��6�;�)E&q.!q-��TD
 �j���E����;����<��n�F/��?�����J�~�yϪ��c��3]�,��:Zx4�<ŝ���~��84�Ѕ�1��u�m��N���s��4楩-��73�p���%�o%�$�K��}>�hKy��3���>:��QbL�S<6Q#x+B�GL*>z"ږK��k3�`�O��r����G�r�6s��Z����e�k�KH^R �n��
>�j�N�������yF D�y j(m��I��r-�>*j�gs���ٴ�fڠY�AB=T!G�N��]���γI	}n{g"�=9��h���	 n6!��^�ڲseҙ�=tgTv� ��h7�çb�r����4�K��^�Y�}�Xt�e�E�*+-J1g���P�A���T�_O�aG��ʐ���h�b����7K-�${{���S�P��{I�QzTa F��ҙZ��z`˷��M<X ����6�9��ﷅ�
������`i�L%�äp������X�L�`B�����m	n��@�,=su�nc����:Q�Xa>�ڟ}�s�u�q�-L��7��mqYm`�����`�o��k�6��Kz���P�B���Z����}�Y����u��T 0b���@G���l�TD/Uy���Tޗb�9(CZ�)��FߎB��T1�KQ����a��ض3}d���E(���	��j�(4�9�� *����H�_Q0G�y\ɲ#?���΃+�@ߣ݂�?$s̙`~��u
z��Շi�������r2U�/�����^����g����~c��-a��j�&�"4D�a8~^�Kp���]�N��u��ɥx��s�Ikv�^�`l�m�>�����t2�)����M�g�Θ`N�z�~���kH�v'��f �R��|�$^��?�y�#,H��@
	EuB�ӘҀ�{������]���d�wf�A"����� �PSO=�V��"�R�N� �(
�=Ma�t�*��hsh8y:{��P�������o���,]9܁iK����N!�,����).%�Ƃ����A#�ӓK\�j���)_�G���7�6o��l�W�!,=�<�4��?~��<s���K$ֹm:dO��X��r�e����*�_�W�&^�E��.�>d�ֿ(2d_����֭֊e%� 4m��}�y�kv�=����of����zT���/SE�iY����-)Ad��G���>��fU���� E�����8�4��s+?~��(fj�#@T66�u���K�Nt_��t}ˑ�m94?��Z���y�݉-�P^�G��ז�y���;r�΅"��!^�R��8q�G�c�"�q� ����B�{ ����WS�!�L��$ӡN�vJ^Z�ul��x���&G$]i����7}�hOH1�
cɌ����/�1��#�12S�ʈCo��·J�g���)t���.#����聋�"���au)�p�Z�i�U.�N�A���y����'"��}��A��	�W܀`+&&$m�@V{�6�d�,xn���Z�F�B�����$$5w�'�m����21�!�TB����i��"ӲN��}k�Sj�h<�*�x�HȄ���B<j��>RP�5f��7
���2��~�!�E�V�T�P�F|��[����h��G�{
�*�������Y���������=��p���
�+ETQ����tţ=�*�^�!���F�*b��&�+4&b+�̍��T}�M�x��~`PM�E�����f���|��ߞĿ�ǭ&cp��w�/��Mk~ɘ� ���:�żO�:@�A��e�v�½�B!��[W��~x%�e3�-�f?��tm">�1-��&;��2�E͸�g��Lķ��?�1 ���Zd�9�����8<�B�@���ȼ�m�[c�3��F�%��g��<N؜�Hl,�z���!��}!<�:��͕aک�0[����nIY�;��K�R\�����X��h&`��p��̆�&��?p��gx���̿����nш�)�3.AW �����U
���s�ɊH"&y\d]�,M�ƕ����N��-�ׂ����/Ϩ������:����m_�$��cf�aaY8��g��s�S�~#r��X!5���N���_�J���;33ų^��L�B��uZ�nMf�����e�>F��?m�u�2yM��������j����w�]܎5�[��dod�{�������?g��
f !����t��l�Hu��ob�bQ���w���Ҧ�`wa�9 ��L�Ľ��E?�������l���=�@��N���XKR ФH��T7&������:G�:����ާc�l�w6^��7O ��D��y��;5�k�o�6�ߔ]�k �Ap�b���4�^��`�.��DPC���C�xS)bz<{�;�I߼\E_Gnθ��[��"����r5�@���80ƗnA�:I�k�=��˦#�U�¦�< ��3D��K���D*����,|�D����6E�^'�n���յ3���C��%�'�r$�f���m��upX�3c�˝�.��|_��*K��kZ��J�Qo$�QU�����^�Z�����ow�G �>���Q���5��|*|�� 	�ݓ.�+b�Ws�I_�Vl��7�vh�Dj�5IB����P��N�Dq>}i�������um[��&?�����M[M��d���&��8��۰�AX�m��\��ݎCe�Bm�n=�Ee��Cc(Yא�Ɏ�#J��,�Ђ�����վFH9��"�b?�l��c8�����Ű�?sQ�i��h�-h#��M��ja��9���5k�TU�>�o>����Ұ�g�I̾#�%��v�e�Q��6R8���Q�ç_H��|6�J93����М�R�=~H/� � 0!��M)�[�ITq"8�l=rܠ��K�ߓA .ʈۓ��������L:��|Tc&���^������K^�;j�3��򋭂�~�ɡ�{�G���Pi����p3r|�㫉O�Q����磒�Ύ�"�)~��J�oˢ�*��{�r	o�Y?�$	Q+L�wJX����:M�Z�"B����)��`{���z���jL�����?6Ւ�	|��y�]1G�cB��HA>��s!Y�����2+�8��e�f��s0E��]NV,��	���?�,�|'�'yޗ/c�.��a��"�v]�r%�x�ò"�C䯯W��i��V�!29ԅ��b<ɘ/.�)̨5���=<`Vr�����9���NE�ׇ1YrE�
���lKG���cى��fƻr>�G��J�^��c[a=�h84��߆�,!���%��� _�"� �����\#�|�������?ԍ�W%�u��3J��L+F�c���L'���������+s��wͳ�d�xv8�;��=?��@_y�_
����#ʯ�tIz;�fS�	(yu $���ސ���� G��=�~$�"&��`t
�S��H�n�ZP1��2�V��`ԣMx���c�AC��e�&\�R�݅��ט�j<�[�L��;���{L�EgGݙ���e51�%G\m�^E�a�O����vA���o��p��z�ɡ*�h�Br �h�!��5[�8�ŕ^�h��H�!ʴ	�4l�c&��������f��m��	E~Zv���
�G;�O��}�g� ��T��#mI�� �3��c�Bs�����"1�IZSx׵�u��) ��X.�6`��w ��0v|���z)�l���n�_���f
Ǝ���5����2h�	��p��D����`�&��A�mrՋ�Ө�t��'�gаw��8%�g�6�F�S���~w�\#� 2����,?�j-���cPIZJ�^h��zv�+LP'2҆1��;���Y^\;�*"{��0���J,����4�U,�2K	X�|F+����Hv�X�dU��dh���D���.O~Eܽ�)#F�>5���������j<��E�%��L �íq/�&���
\��0������"�����gږ$,�r�i�3a����s�^;8�\`�l�q�����緛I���h�/f�i�v����Z�>F����8n��{�6$�_�E,oO���:�/�K��fr�v�7�-��1]p� o{4�MSWţ�ʃ]�*
pGU0g����b�2+/�"�q��21��ZLg�U�|�_�E�v U�nW����yȥ3�N�ڇ=�=��.��+�?5��O󁈧l�|��>����z�A�$V�����Y ��z� *�� ���~��k�s�|�Iim�1�O +�E�y�׿��������l u߶?�i^ߟhlvW��ng9ܖ�̽�y����t����$ۿ��SE 8�������|�Vr0��>�	Ku\x�~�1�t�k̐^MA|V�矎��v�$�d�;�z�qk������]�V'�l����F�a*'�us��w��+_�(����wD�[�Q��qᶀ�F\�,���ט���*�N`�|����oӱXa2��:�$�oqem��e�+��|kl�U>ݤ������ra{���X�k΢n?[��5'M�X���y�ݸ��ȃ�������凱qۍ(�P
�R��L�cX�V�J�׸:�_����[-��\;�3?[�HC?��'U�x�<XO�����12|�U�����������p��ie9�-�m�r�E�j�a+b�x;)]���5Ҁ�k����
��R,K ݫZ�YT�EB�ĳm�4.�߼1�����#
匔���}é�A�Hz}�<���2�9B"%��3Wz]&U�������)8�`�ߏ'H�{*{d@!�����P��VR3dv�7&O��Ͼ��F�J��z60 v�����E\6��*�jM8�P����(���'��W�y���-�	S����_��Ȥr��WK����0n�풅�u끆��d��@���������S|�~���a�C������F�,-z=�'��XU+�@	d���)a�H��iX\i25$]T��W�*1�|�`�蛕�rи�堬2�61چ��껕��X��� ��RG���Q1��A���!���
0Ƕp-ܧ��*5҄?q,��!�����Jk��D��s���U��uD���RR�ͧ��>ƦU7]
sc(����pVU�%��#��&��pL�w����f(m6"�d��{Ӏ���h�\3�2sT]����PU��s�Q�o"Psl}��c8��?��{�}��
$��������[��M������#T^*(C�e	�>h��%��p�����ji'�/�1�\���/"8��d���a��ŏ(r�}w!�a�ևؔ�R�U;ʾ���A���
�T���})�����Lq���o뱤���ض�)����K��]ۺ����돚���e����B%_7��.`u.�ks��D�rГ�#�?�ϻ#&��3�%�H��$7Z^��ˁ8���@g9n�����S�Tt�/;N�'��bݯ\j�<�X�.�?(�.���=+_��|rr�"��9��6Ww�g׵����Xý���~��@@.��]��q�m���~Yg�]�z'�r�`��K2b��9���7��u�1�]W���o1�t˔�0�-�8I���0S�^�� ��B_�u���F�^v�����860-GHlQ�bO�o*	��`��}�HM��ҦČ#�im�Z���
� ����C1.�9j|�z��C:Ӳ���k������Ӻ\A��i��a���r�b����n	�19���πs�遙Cb�>5W~۞���pq2#��g�)���d�!�}����Ŧ!(�
V#�w#A*�x���(�LJ��!���j$�
�p�����[�9�2��wWM��꺁1{��D�jA�=J!@�V�rU]I�3p�|�V��k��R�-�&�~�ph4�H�pd��e�.͞%��0��w��8,;�Jf�,�sR��כ��y�Ԁ�>�^u4�%���u���+T�MԼj����f�8��<O��ln��!
��k�ߴ��,iQ8w�}��ÂX��V�8VV�A�!Y�&���z�}����v�OG�����Uv�Z�%�n:V�K�{�����fF@х���4/u3Y��9s���|�N��<������E��?�1��`@(5NH����+׿�Y���uk_�12���~��,��$��� �!���S�f�ӯ��fû�$�����h�[f�%�L-���Z���4�,�cf)��|��@�$����a�&��5kHsh��z���zGrgl,��j�}	@�<��{�(5H1��8i׆��k�jÎї�z9��h�e+��u�5#7�0���\���11:K?$�Vlb����3�İ������Tq��8���\9n�@���3u��b&�I�\�C�Zc!)3Z�R��Ui�욁��d)���κ�o����?Dt���U�w�z�bbBk��B״�`%@E�0x���4�w�����W��j�2
;�	?\/�
Q�b��B=}�s�P8�mwITu`:�䥘}F�}+�g���
�7)#}N�����x5�v_�v�!�K�޿�Ɣ��3�Bʒ-��'ڶ�k�y��~��I3���2��Z������!@�5u[1�Z-���iR�{�ŮG�
xa=�ИR�q}W;��}�n�Ab֒�f`� ��Ql��Z{�K
�y�������M�����&�\�W��¹�}{� ;�)����d�4O���=�yLB���őײb���@�y�E#B�.�����}�<�uw`��srmo����A�m�
�`;Xc�j�<}t��{M�H��Y���N�B�x������@�7�f}(4�7�O/�xy.�\���u{%�:��dZ�����ܨ5%���U;����)�
u�1����M;&m�K�dF�����||%�#lu�j7|PJ��_�M�T��0}�*�P}������XŸ��r��#��T�Tb��{C��-��X�	��n=��<5�̰��nq��������fd�3'a�=	H�$�����|^]�n���E��+t���.zk�����)�V���5p�{�c�����!��_c��u�nצñ��!#v�&�B�X��~��c�_�>B��N�G7re�u��h�=�6����җX��dd�m����C��B�u�"Ks�Mʰԅ��5�`݊GMs+���k�;!��%t�������)��	�L�"�R�u��/��~��Z��/Y��I���dl݌s���~c��܎}�މ%P5C�B
���]�	���q7
ʄ2�U�u��"��U��,�t����W㇡�C��� ���F���b�W!�u�J1J|�b�ʪo�/O.�'7H6)|�c+�n����e�p��a����a(�r|?(��Y x�ofV�8���']����!��f���Qr�'+��
n~��s")AalJ���y��¼�S$��Xq�ψ3��[�BF�ZzQ���:C0���>�,/���~3o`��O��
�DM#F^XsU���3�Z@�l��Df�n��I�Q��!�kP/\/��\���\·CE���<d���+S�U��&v+1UW��$��|�K��Od�/�.ˆH�0��4�9������w�2���.����(xD��1;�����(����%�s�y���@�Rw��#z�K�0g�;E��⍌�V԰S~�k̏q�"J��S��m�������KHy����;��޻�"���Uin��i�XkyY����1���'y�N.�ȑy�`�]h�X�lM]_�29�}�ô�𓎒;ӹ���QH�D�xP��ʐ��m󶣅B����p��]?H�m�M:+��}a\����SNaJ覐ر��لxu�U'~�'������B��:'џL�/, Q!��/�E���-s(���v����3L�aA�G�37���V��@_�Ԫ��p�i���sĕZ^���ltP{.�!C�m�?b��:��)���>�;�����Z�m��A��>�j������)Xujs6�+��=�b�-�Nx5�w�W\.6�H����/��f)�+X(%���Iq�OI㉐��a=�<�[���,
�����M`�4$�1��&�VW���#���~S�Za�V��)��e�lON�������`E/�L�d�%� �g`e�&�Uiib�R��#Tv(�dFy*K�ܫ�l��?m=�NM�6Gy�#�k�����C��!r��~���=��B?϶�4��6��<xvsve(7E�t��v�?��_�U$'S���c,A���~¦�8�� Ôu�mM_�@���$	��@����n�~U�[��s���&c�V���9s�� �z+�U����
!��jPa��!J�e͋'Zu�EZH�7��ZC���t�F���|��$�
�XA�[8�~���.,�/l�K���6_�<o��o2mr�8}mr�MpMk`V�H�*�iV(�m=%���G�p�|\��aɛ��B�ö���D���Y��:�BC��[��md�e��+n�:���$�U^/�}=Έ���D6m�x��D-�~���f��Up����>(�fs-[����ߠ�z..�-�@;�9��t= ⯮�COт��"�2�2�*k�Y`�V�����ړG�qtPB��	'L��'��!��!w�P��;e�� {�7׫��LLJ�"�c���"�X%1˂�qa�zAI��IȰm)&󱐖�b�CXs�(��>��u�&�}<B5az�(Ĥ1����i�'�	�<Ї(R^��_���nr<�W��o�H�9�;
_H;�b�ʰ��Q�7��XV���#̏�f���E���}Mcs�kU��3{)��#��F�^�Iq3���=b���L{�3�",�|C)��K�n���lÚ��DW��J'�&t��qF��i⩳6	(��߻��<@���q�.�e�"��cX����Ζݻ�s���2<������d���i�������+|�aN��Z���3��O�,쮭�	�O�U��9�z0�3M�s�7�2�Hx��H��>-�/���#>g|*�#|��i6���rk*Dzq����̮��1��	XQv�*�E?��q�B1J�P�{�u�Q�����O�)�������N���m�*�3�z�8ݐrE`�
�ه�\�l5�s*WL�i�g�����{u>��+��P�D�g���5�%��5E�ŧ��T����>�0eθ�g�䫻U��u��ƀ��e���E���P�%���e*��N�L�jgݨ�@�w2Qӂ~�?����(�!@Υ�?���ԡI~�5�E(_�@�0QdI��K<���|���;�5�U^{},�~��&�Wb�77"%�K2md���0��`v������ˌ���*w�<i���T��owZ�i(ί��bL��W�{J662R�l)f��l>��zH�e�1��lW���5㽃0�q)�P�D�c�})l������n�ӰCs/�_D�pYE�7�������ė2ui1]n	�9l����������A���qؐ��k[4ʾ쳛p�'�� "2A`J�:�X�_����4b�!P���,�1h&�?z����К;��6��AH��IM/�i��aߍ��D�N�[Y��j^�����ߍ�HhzX(��l,Y��kXO���Q�p�ޓ��a�}���aQ�i��_��9N�MTɬ�H�kl���L���9�����#����E��p4��*�)n��t�9��� և����z��w0;�Cjr�Ǒμ��wg�T��$B�A�Fku�Q�O�u9��Q�[�bX�v��Ď��s��F$yl���s��f����i���r�5��.I�SE�V�Zkw���8l<Q�q�Jr��y,T�a�*~`���b��/<�h�D�$��Wϯ��6��	�c���6��O�OTы���}�0�c���ا]Õn���L���¾�>�n\%�r���on�FtÚ:�8wɿݵ��Kl�O���0��*�8z�E+�2M�x�b��Þ��Sp��qu���+ϟ��G\H0R����1�D�!C��7�C�]n`&��YK�;wp����#7q�v`�����g0�3&��&���e�b�o�T��I����"3�@P6�[�:�X}y���R�lyÂ(�B��`�Z������3�6�4�<�A'�� *�/<B��L��� �U5��Ae������3'׹U�����x|bp�I�^y��v[mX�_�p��Tӎ�5{^7$���n��R@��q �
4ϑh�+�9�j��\��sǄD�����|JKl�x�c%I���\�\����ǲ�|zAˌf(m�?��r��平Lۈ��ԎN�h]kpCub�K"�OӖ`{m�L<A�ݔ
�/�9��<�)�q�R���E����h�D���[�Y�q���̭?�%!*�z8�4�Gx-29k<ѧ�%�.
�rB�9X/C���[Nī�~<
�eo�|T������`�l_��ʺ����>�g�[�挗���4��&�!���Os��qc��D��)��]jY��_1)���ٌ��)�����wXz�r�&���BC(�y�K7{{�n)�1��O�R��_�5J�)�X ��eU�>�S�;�h^I]\�"T�*�`.��YM��7pW(ࠔ\�=sX�7:Ԗm�B�C��̍8ܥ��X5����ե�з�=��}�7>�w���}hS�u�k�Nl9��Eo�QM#��/��6b�8��)zO�5���.}���t/<q�yRow%����	��O�7�O&����M:Q����<��N
�\l������b0����o�����x�x�62"f��j2�9�hQ����%��[�<!�/��q��Zy���l��i#�C�f�(}۶��]F�\���J��73"�fg�,���k5g8�X����0��<ql�w<g�ʌz~,�OD};y�9��i2e鶹��
�Yg�SSߥ`/��
��|g�oPz%&IȖũ���K�U?.�.�f���T�+�:̞z��w�5V?��"�	:�CD0K�6z8�.�tH���6�<���S��W�Rf�o��v���"��ש�y�C����\�Z��ʚ���>��u�ɐ�?�t�9�d��+�jM��
U��K��h��'*RI��QeQ�& �D{��o�����5�2x=/������#�ԙO͟xC�z�rO���g�Z=������w�gju�S㠧H?ϰ�ॴ��ݣ(}����}���X>]`�,O���y+���p��ޅДM����r�|!Z�{�:���!
Q��xc?���QV4�Ư>�y�2��\��D�ā�Wγ��/t�@V�M����3qX�/�0��o�"-�.��9K�[ �F �W��5��S67�:��v���	��{<Q���Wy����mrL�1�D��@��9V|Ib��:H��� Ic����t{�ajR�l��*�@�) �oq�M���~�{�F�(++:���
t�7I�>	j̙dU�_�-h�I�[d���P�1Jz��6�#L���9+�@�]� 61�
3�D���Y�[��� %Z9�s�"�i?V�@��J?Q[�\�Qy�����؄a�]ݶ��;�n6`ߌ3��6�8���� ��a�ۣ��s��(��R$[!�ڔ
�O�[�����"�@򒫟H{q��>�Y�E���C��Q�J���j�-�S�c6O���5X9����+ҍӑ$���}1��2����鮘�V8K�Ga�UM�u�0j����r�>�A�N
�M`$	MT�G�&�ߵ�F���CٰW��_@rv�h"�k�10�g`a�X,�q��8m��I�;�������U�BJ�h��J�VhtnYܢ'�Rۦo櫓M!�yq����lO����0��riQI��	c8EX7��"P�vC]�D�ə9	b��)K�mz��1Oӈ�ʬ�-����,sKvx�%ۢ;�.��x��}�?$�Z��44�R��#��X�G<٣���J��c|"_ '���z=���IM��� s$�hh�u��(�&�0��!tK��+���$�ֿ�q���1�nl)�Ã��S4~�kgR樹rzR�����3o��4���ː.8ou�ܮ�����nq֑FQ�r�y�d�gO6\L_��9g�H���?D��b��=����@��@DD/���U���"���*�=��~>�d�g��|b����|�6��;+4)�hJ��/6L�U��'�l���~n% վϝV���H�,RK�-x���l��O����m�J�sg�+	�"�����s�?��S+ Ǐ�IQS��P��Gtg%�.,�4�%�_N��g�l�����,�Ե�XŰV�TГ#���lG�4��V_Dz�K��z��l�Ww�I�Iݮ�ڒ+eV6����&^���[M|$Fy����áxSԍ<L?!�)r�iȔ��������T�<�knMcsHY�#j_��w��]j.wea��5�􈮷��V+�KN<��bŎN�MhT��5�,��T�:^��O$�&'��� m��ҥX�v�����^{6�4OֆtQ�ar����e5|���P��ZKf�R~��ُU��d���a�8:����R>�"��.�(��l��S;~Ѽ�afU����� ����x���O�,��Nb����LY�92q�2)�=��UC�M�\'�*�YS�?`��x��:+���KKc�Z�ƻ�ZP?_�h�P��1�8��/L�ӮeʉԹ��_?�2@7E6��J�]_;��l��B���*m��#�oА����2�����NYL�%A����;�V#��
���PŹ�Hn�5~�d>l���Á�u����g��|��@��#n˼����v .I���*6���9�7��&3��� ��;}Dڕ2%�&U/ ��h�4H��!��9h�ۊ���Z����3��z��踛��,m�1�mes4^@��%�XR�->�"-�<����y��^��'h��a��4���$�>�T/e�)ɔQrk}���~p����(���i�
�o=��H6���� �:@�?-w��YU�(����>||��\i�PG�l�C�*��`���p��@mY����ˠ;)�R
	.$��#��?������&������+�u�� ��~�\��*��y��>=�]*��]���w��F��X��k��`ڞ�s�������Yv�@x%.�W����2)�J�vd觉��؉�Z���w�_�F���=��Йy�d����O-����,0w����*X�!�MA5��H;��8���(5M�ڽi�{7=Q|z�hn	���	���3�E$���ۙO�֔Q��L�:�7��=���M���Z�I�r�9Q䂫��sq�wc�5Ő܊I��cRrHz�ʹp�N:��N-�-m�y���Y%-<��@a?9���F�%v�<�=o��N��
?����,p�r�$�w���#��)�}d�E�M��A��B�M�Q9(ּ��_�jV���
U+�nH�i�Uì�?�=��]�1O�c�@X��e��r����Z⣙��y��"�f�P7���_��j��9K�@�� �6t�ϙ �C��d������V��ʹ��t��������<� z�����	 Q1�f��iy�P�~�5D?�ХOǢ3�w��-6��#k�I�0|�&}�G��9��E�D��*��G��r��](���,F��g&^����Q����Ή��$�8�g�4�Z+¶Q?"�J��`�"��,x;sԩ|�c�^Ӯ�@ D�d���� �߳�%ڱK����9�5� ��W����ϲ� �� c�;��]���$��"٫؊r�)���ɇ��F)zi�`T�CDuܥ��pX�i�yHCæ��U���%��>����!�*4�InR�N�8��B�qC�^�S��fT�B �B`s(��x�a�z	�R@�oA��� Hg@*6��7���MCfd��6���!|�Nv�9aE���?P���Y�gf<o��]�ޞ=��$Y%2�uLM�V���Y���C�,t�`0����f@�޺GR�(������n�/����Gğ���U.SQ3$�ڞi�p������޼#�@9��>��L�Lq��YgE�)���2w�y�7�}\�K5����e�E�sŊ�9��y��8��[��M�!hpw.?f�������3�����P�Vͧ��E�zE�^k�� Z�P|v%�8��q㓯��r���i��h�Q��#?E�4�Xb�-���X;'�ex�d`=:x|PNk"i���?+�k[�ʤ��.��%���,�y�	kY��'ϖ<u˘Y��A�('e��):%�(V��.�	�z0 ���T�	@��-�A���{����q��x&�[W6z�/�:h�Il�̹��0/��D���_�:f��y��[) ��
�X	�g� �<b��Ô���,�����'���s��P��-J4�¹P�П�8�_�:	�}���~3j�1�O�wtD8���N{��W�3�J������:1W��㙠h�����uS��J���"˧�?�>/�����~���x�� (�.��ҝ�܎o��Mr$���P��J �8��|$�ˣ����u��_��V�W�*��nmF�8����:Nدe7�b�O�6J�����.	�"NCI�\$^�P�
��GEl�Ѳ3Ԉݚ����ɪ8������eć�\t�o�5���@5"�h�كUc-1"�9i{�Ih���o��*nRt�
�$�ߙ�U����v�f��l�e�\�;(p��gӞ�
�����z�ڧPl�����/�&y{���k>g|�i�R�mC�Y�>�b%`W����@r���DLy��ij3�����|�3e��)���*��8�<����L�D����.q�}`u2�_���.���,�0�(���8��\إI�?�!�r  ��j�y�����߲D$ۥ!����z��oI<Nv>c"('
��3�>�0��Q%��Q� ]��oz�>�$d��������_1������?��or9j��R�t�梉�:#%�L�M���4"�Q@$*R�ک�"�٤y�5�Y�eo��T�����P�j��"Fq�ߠ
ݐ�$�Y��ؙ��y�Ɨ�F&���X�?P?��괲x��S�������;��v>��=�1'<S�2�fT������w�&��@�]�*߭!ے���5D�;i��`(�q���+�~���?����� �r�����gϷ�rJ�+��� g���Y;�Y�ٙ"���>�ʤ¡���mo(�sk�oj��%.��<)k&qcݗP��O��;���>xx|���E�T�#��!=�86�[�缯��M֊��ѷ�OD;QA�!LKl[�=��r��4��_�O\�c�r�o�j;��7�ӺJc�T{��U�)��/v�N��a�ߣ^YB�=%q�&�bd�H��DA��/�e�an娽��G���R]H�޹�T��z��>K�u\�VA��gúG=��؂z�:�y<��R>g<i��J�Ϥ��,�)�s�������ix2�Zw�\��E�C�h�?/V��}��n{��py�2ȍ"���O���ة��L����mϣ2�:�k2�������}LHm���D��x�����]+~j7r��l�gXF>I�e�쥦�XR���h���.-=5vʇ� p�4�\^V�~��>�w1��f�����0��L�	�O��@5�`��m�$�� �n)'ԙ؋o�u�Q��|婕�j�_��t����Ξ0h�{@9����h5Fh�J8��Ӈ@�R����M�?��_�^N����O�K�/��X���PR4�Kz=]1�����	읋�FG(��	��Y�o�~���/<L�@a� v���^Ѿ��٢ހT��\��&`�~���&���^�����p�9D���<��4Y�kD�*�n(��h���	����Be��N���������?k=�s��{��x��ҫ�j`�;�??�烁M�����~���e.��pR�_����fO�]b�V���:�ǌ�C�0��c�����j�f�C^�^����3: ev�xOx&,����
�3�6$u)R�J^ oZz���T��\��g֟�x������vp/�����?tI�\����91ȸ#zJ����[k0�'��Y���2UX�-F@�Ε/^�*|i���(Q�+ja��T�ԃ��J��	?�ZZ:��GJe }��L"|�q�6ım������Wqɒr��jH�o�гv���v�mA��Y���SG�ʕH�n�"Jn��>���~;h9h�+v�5	T?k �E��wG��0�-ukPIJ� ��G�n���_��:!�5:���4j�'|�ƅ�]�����v�@n;`%AeI9|JbhS)����}[����N��+��a�T�u�W�S�ې�L~Z�~c#'=4��l��2�i?'UDU~E��(�t!I�c��^S�����74N)zoo
k�����I���k�^#Vס�g7 c��Z�Nx
�s��a�lZ5��-��hb������
���g?��S�Ob��l��ڑ� �ƉSr�̠4�L�p�U����Ĉ\�͉!Α�'\�:٨�$@oԦ�,`�j��&#!Z�����2���<��97��k�V^>�z!���������q��9R{XV�(�賤o�H$ g*(B)R��W��@}���X;2m���(��j��E��߹��` �`N[�~0�vY�=�\K��C���C*51�;c�g}Edܮ~�,VY^`@-����n�Zb7�'w|�-qόŋ�p�'?wO�}1A�z/�JGh�� ��_!@�i��M7��	��Ɲ��ڝ�J�Ŋ����y��m{X#$���/�[f8O��o�
a 61��yR���
�[���f��F ���Nz��\��l�P�{�FZL2~�v,Q��-�=����c!	��������đ��WO6�����U�^��)��G2�&�z����/l���B��Zj���v����N���F��Ѱ��	�[}���Yz�aP�t��
�2L�K����g��S�r��u�P{�JIy�X		�O��8��uT\ߏ7�;&�>�[T��@��A q| �ѹN��+��-6-���������a3�V^ ����zW�3l��=�ʚ)19�N���A���h��`� ζ`'�Y@��<h�~���Ȳ��u.N��R��U��1�� ��x�l^[.F���wb'��r�5���W���`&{�����8��.:{����^A��@,
fw/�s�X;_��GL��h%F�ܙ����f�N��<�]�z�(I4�꯿k��16x�96�6ʱ�V�����dz���s�o�Ih(��c���g(e�Vf�Y�b=.]�>4댋��"��d� n�N�?c�d�/�AJ^����XV	f� �i ǮOH�	�9�:���)�~��&�4T���)�ĊV��;��Ҷ��91���&n��0E	�E����[x�"�O���bD��` h�96(��/}�X��Vv�%Ck��f��X�f�3ʃ��X�D�ܥ�D�Ŕr���XXb���q%�Y�݆�Kd��J��Vָ��?�ޠ�wA���G�w�8�<�j�c|4�F�m�'�}%�A����m���%�L�J�W3�HZ�d�@Eq��ѧ0�mD|���ָ)���)d�mn���f!�tZ$́jγ�h����N:զ�a�*����g�e�_��k�D4p���_��9���E�E����n#x�GtG�e���6)���^ڑ�|>9yẐ��>����q�R�e2�w��Gx@��L��K�-�'�a�l5��|O�
2H�3\C5��?6�D
 �����L��Д��n��6�ee���Ӄ�)C�%<�k�E��T<�(� .��Q��3�H_aؑ�G�;+���3hA
u ���ƀ���n�8�8��b|�2`�vb#�������r�o�۩ݹ%���ѕYm��/(ߦ�:�k��֖��z��~y���Xx�_ke��C����,�>*�"{'�v���/� ��l�����
I�q�˫*��s��fJ���V�����ki�Jo��'�B/���E{K��!q��@�y��2!H�ZʦV�݌���q�@e��Q^���j�����c��z3��n�4X�qm�N:�TQr�1Á�B:�q�d�.#¿��N6V�b[j���Up�K���r�����J�,�V��8�Xcf�����Or��0.4*`�#������ٯ�Oz��*{_Z��t��i�X����F��`}7�'r}�dw�������I�����������^uZr/CU��%����R:�DOf�Ąo��;}�j�M���\�؂MN�eK7/䧴��5Z�D<wi�VOd��tM�~��J�V���m�mE琉Z)����]-��{-��ͧH"R� y@�����\���׋[m����~n(览�$<�ÖM����ua����Db�q&1������ֲ��*�^�(琂+ǚ�/<E��o��0�Љ(]k+`D�m��&1O2���q���#P�X�@kx?�ͬ���!��7���#�9�V����D!���[����`�s��J���+Y&�;�^��HKi��>%<"�g>_�*K�*6�rP�/��![���]���s�� �,����?��;���+��'G����C>0
J�ɮ��� ��O.;z��ED��e�Q^Nj�6��v=
V���δ���>2�� Y��E��R�5!J<�Z����9;,��R--����8���|P� ����׽�3�I2s T� �����s3����V	)�����_k(P+�u٘�IK�k��0G�K� R�RM���V5��l�\�.�z|�LG�L��%A���7��ĳ��-��چ�)�D�c:?v1!7�7�p����s1Dx�;\z�T�l��}:�+�s�Yq{0T��f���0��?��LT)�3͏������{ĻEI8Պ�ܻ���b�za���q�)��|\C^�nN��|me�3w&��'ot�?�=���3��Ӫ[�K���%��^�c�[N�Z�<��]"��� :�Z��~�5a��}NO�?Tv�_�hd��m`(`�fe���0u;H!o�p�s���~�TI��i8]V\�@}ƒ��k�i�R�ҟ�������9�|��~d#��BfE�yɩzr����ևiplh�8^�qo�ƍe"��`�1/���V�/������R�?~�x�C�K�k�{+��V0���%�bw+|�p>�������fD�5]�K�����\�+� ���9�v�:��M�"�P*���s�/Щ~������lP��gY�J�-��%N	RG��O�X�7�3�3F����>r��~�%M��J*Kp�+���/�uP��uI)��0lr�a��Gܚ�f�Ƀ4���@��$��n^�<"��z-]���ق
j��&~���i���xOD�_f93}��;q����-����Vi�b�5Vz��:ȵ�SsX�B��~��0X[I_���p�^{�PE#Ť�����]V�E�iu� W6����]@��6��R�Dq֗��̟���f���m�Љ���c�zq�B귢W�^��ػ%��Rs0@h�m}�X^ݻϳ�V-�B^��6$q$�'%~���)�Ѫr��~�aʶ��uK������¼�3��H�B�&����Fo�i��:c�ͬ������V�a[v��^9��ay:F�r�R��q����Yl�it�J�1��ٳ�8EL0��A>�����$gj���*�E5k�xC���|aA���if�_��ٛW���L��F��fKa6�Y-�r!9;; 7E꼐 a������V5l�[�8��uxм%EX��|G$����*�H�����;��O^��u�E*Q�E��%.h���t��e����iu`�����%�)@g�@�Uɲ��@,�E9|��"B���Ž~(�ϴZo9	����u~��v�AL_�ɜi��{���Ƶ���O H>�S������Z��Ue75������9�pzs����Π�op�F�+2m'\��a����2�d-�T14])
?\]�ePo`��y��E�J��8���p�IV�c'#��?��W��� �k�����@���i�j;��~lΞI�Y�m Bq��I!�:�|&v�Ο�"��V�?���&��K����z�U��HB!tZ��X~fv~2=M[5��G*�"�LӮ0��̹�8��s�j�#�
�oW������S���j5Γ��bӸ�QI�ڊ�?��#\�3s$����&��M��'~�~؛�f5�t)�%X6�A�����k��h� ��DÌ��yӓu�T�l��*�������~�"��3��-S�⨣�ۓ�<��qo<���>Y�7-}ߍ�� ����ә�(�P���S�$'�$@V5O5�QV��=>4e`OH�9���hi_�p��.r+R|�x�u�KrE���*������В��-@؆��c,:��V���p.�Wޖ./��^�0�
|����E��1�{�k�7|b�(Pc�\���Zf�0������Z��^���f�!+CH�!}��]�����Yq�0n��N���(�CUֹ��3)�
?n#g!�?�H7-���8��i�Q� )l�#���z����[ڈNb��p~S&�t��M9^(7r�#㱁�/�`�����fz���D�#�����(���#x7�����Ƭ��4����l�N��8ۼ�[�8�ݓ����#rK��^n8��t�r~�#��f|A�G�HϫV4���44�c�
	p��8=�0���e��	Diۏ�(� qt��/��+H�Œ�$��dVpk7;dɦ?���̶�qra����\�'KԟF����Փ;�A2�~���  �R6�<�F�֒I&<���~�Rܤ?�m�3
$�_��`���Y��H�7_�2=�yz2�s��p��?�K��%Pb;!��߿�nIB��1��.�!㖢]c[�����U��C��������n9�Ex�� �j����b
!ޜ+�!�3L�4�b��0V�Ӥ�^36F�{"�/zT�����6�:UB��R��:Dʿ8f,M!���̩�.zz&�V��xxl�م�a �e�����yW�D�?.&F <����ٷ<�Q3�)�E��9X���=vy�ި������,�l�#��J�nr�h�[8u$�^�%�NŎ�M���Eg�^�Z����G�`��י��J����:�{�JA���KX�������'\�>P#�'��x�x�m��i�b\����Ŏ4�w�̖*Mv�?Z��A�YL=~;uDj��s��2�#�9n�V�j�d(���!���K��+�L���D��#��0c��Hr��y�)vǷ��sT�W�:
16ڄ�Ym`D��Zj��E��{P�Y�կ��I����=o_�藁 ��yb��P痌��W�z��>��P����R|�_<; 	C��F���+ DK� Ր-�a���e':���ܔ���U��x�c*��J�Tx(]7���E�I6܍o��ho�7��X9�XU��iQ_�X�ci4�G��A�9�I�4�H��9x4��ĩ��fI��V���x��=?�SM��0;��$��_�Y����߀Y����U�x�ՏQ�B�v�\1��jJ��'\!c�b��d��p��*���>&E>\�ktU��{t�~��VN�$)��2�?Ne*Z�צ�ˬ:�L�bdq�x�Q�$�A��7��К�A%u [������������N��eH�5T��i2B��a��_����qp~��ҳ�՞�	���H����vx@�(������V�X�[�$����$R^��V[�=v Z s��NZ�ag5������~?���l�/�Hm-�����i)A?Sq4���O+�R4!V���n2����~�z���fꃥq��U3R|d��;�^��s=�B�ނ�D�yb��>��i�$�'Ԕ~���qL���JJ�b_�g|DӺQ�"Wׅ�'ɚ����7sJ(S��뛉;��K��5�H�lԀ�3�2�� F~�gd�iV��؃�9�ީ�N��ŸA� �B@#������m':)�wΰ��#�fNG��?�*E���*Y,��̕U�x�%٬��?�}���=zc� k/O��?J�ר�qđ�F��=L/�n����]�.hn�)�J:Z^�\vo��7'����Q���]}��V����M1�����1��yl�Š�a3�B�=K�>l���>I��'�g�<
3R�%�&��]IԄU�=��׎�h�� �\k��+�x(�,�Ućly�{G�M�.�,��
L[�ڈ>�s�7N�i�h�q�Ep�RX����쿺���_@������Q�[|����F���HГ5@W��F�*�`	��z��M��?�z�Ix��TU��uBڿ�@�ҋ}�������_ A;�05#�~E��F��N�ӝ�-2���﹢ID��Ó���+Qr���Gu�q�T��"y��[�:�8����7_� |�FS��G쓹G�'�����Ю� ��ҏ���j2�4˳& ���;*��[���-r5��ހ�������6"s��_Q��(NΜE��:*#�m��J�����溸>d$&����\@��,+�� ���i��g�۠�.x4�=*���CU$��rx���3m�c����T.��Q��H����I�f�)�u����G�d�+�,5���[���XV/~,a�����6�|�������!FX%��88�(��v�pA��st �{<ld�ʳꩦ����tKJ$��]`PQ;#{���y�*��$h:��T�]~q�[30���:`v\�D\/�o�]-G˗+f�{;3|R�Cn"R�ɧ�~M�@���G����Ip6�;'/S��h	�7/dU֧DGF٪.+�k��'�Ω�!�a����y\� �	�)�/ ����uXDoU�����~��&l�+θ�se�e�=��s䤄��@��I���-��:�Y�|�x8�ah����+�����[���K"�Q��Ǭ�?�H�"y���3�����z��=�;@U2u��mB�ǐ,!-:�-\�hP��ݖ62'��C�d��@���S�}>�[Yvm�4AM8�g+�"�h>�����GZ�m�m��T�k��uaQ]_�d}�M���`��u�|h�����ܢv�%���������w��>:/���("g��+5�&�ˮu�fh����`T�<�%��)���d@P�1HS�,��Y[�I���DL��NX*O��d�Hxz$�d�n�G+ǘ�>�)"�,��;�*���7�����m 	���pq��TQT���7�PP���Ƌ\4�� ����]�Q���[�����3�dJ0��G�n� �2����C(	��ݐ�+}7��c]S�hW� �Z�6���n/Y�pt�?tR�>@���u��E��8��Ӏ .�p��TA�n��l��M"����a��\�����݁��-Z�2�a#���q���	�7��E�Y��d����`j4 ���mC�7o��Mc;*(����a����Z�$��fw	ϸ[�Eb2��F�+�|ӑHU�s�'y��2�<6cQ�uz���F�<ײq4�eN-8�.�ɂ�;t�0E���	�wH���*��fQ�M!^s�S�cU�~�O6�7�LXS�I��y�]߁`�ٜ�/v��//���\"#��R��1G�qo7g�Jȶ�$���lrU
Y�C��o���
�1rv�U%��G��T��T�O�0��?
�~i|0$I�W�>�x�K7([Em�/���O��z��<<Gm��2Q�̶���M�����id�@֦1�*�T�K�<a,~���s��ʔB��=���,�=~�W�_�����Le����;���v�^�R*}�:�$�� �R��;�9����vK���R�p��L��c�+@���Cko�����5��Wb쿛�7�e�����A)n��R+S[/�,�=�b(T|��t�A� /T��ilqN&|�O�]�@6A���턶�ܬy�еpX٩�u�.եO�yo��s��b�G������1w#�0m�̈.�-�P�/����`J]B��\�E�ư�B�]A�},���	g`��\ؿ�zui"b����l�5�R�i�=��cH/� �?+����S�G+YG��|}k��r�5��n��t#3�YA��a�|�;X׋��L�_q��&��N���ѭ�D�Ӑ��}���v�(�?"��E�80�%���H}��?Q�h�cu����U�p���	@6+�-�D`��nO�6�T�:hҫn�u�QY�C�J޿{��B�K�q�u*��ة�Š���D9����V�$h�g���4+P�-d����$0����`ѣ�ԑ��9F�O��2�]���u�SXR����^�ʧ��򽒛���I��Hwl0yŀ�[�W��O_xV�K�gL�dНP�ڨ�/G�^�b��R,���N0:r�`��E[ѧ�%�_o�߻�^�p�+�]� �iU� ���|C��v2C�/k� Ng �A�$�ؚg�|������,%y��_`����x�(ڧ�6��A�G;�� �߲X�.��;�j��R
o�S�ģ�zZ�5��0��Н��>�/P'6fV\r���?�>=�|A�z������L+����A7�Kl<��\b�׍6
��Օ=����'��9W�<>A�L=]Bv��ٺ���g���������dI#�7�!�<t�T��Z����@���ʗ���k��b�R����b��خ.}5+�r�#z��H��|�B��Zqh�f��/�s X(�=C�����:{��.r�4�e��ea4I�ٗd��M�t�HP��@�
��?���%�����ꂈS�-��x�/����n�\wH���uz����f��AFs�s��[�d�ԉa	
-l������P�<z&4N�;�a�᱇��i4����w�M�}qy ����a�.� M��f��3�=��pT ���޹B�&xzY_�kL�'���蒊Y��C�gj � I9�����<���M�~�:���b�;���.Iz���~��m�\�8�˥
�'�H�Aa��x=ho7F�+�1�I��hgG��瘆Ey�cG�u�e����[�S���f��y�M{����Ǖј�	��HI�}eKܕ쇈����;3m!Z3|��(O��ґT�t
t�gb�liǉ���.
ShP����Ͳ�)lc0D�m�FR��*?� �Z��)��?��DK��<�vX�R��l��� ������3W��:։|����e�X�Α}1�r������o�N�y�7ke�ȣ��\FA%�`�ǫB�U>��M����&.u�kD��'k7�	�-d�i�W�'d
�v?���M!�`��� Ix���\Ka[KI7��װZV*q������b�2��)����s�PWz�9�:XV�A`_a]F�'��������.%
"�����Ӿn�pμweh��o�DA��`�CR�`v�H����i����&�':5� "#s�V��̜y��D�FS;j�Djs����J�q�}��`.���i���C��nϦ�o��%Mׇ���&j��mر�-�:�A�2���hF�*��	��i�r���e~� r�?\����
!2�62�H+��kz1v��dvf�J5�Xt2��L��1X'�~N�(k�Yn��>p�l���D���&�i����+G��L���.�;�9%���쥺���@/���B��0�%O�jh���fa/���B��� .��\b�>�rf{�o��h��qD����hg� ��F8ɑK�T�0֬÷���6��d {j[@�{� �N�U�8�)1ɆU����SBp�V���2���z�A"��������M�-�L��"r��C�.�9`�nT��I!l�]=(rɳN�q&�<b&�✵5��
�T�E�(�4�d��Vp�k ��x�/*z�Ѡwc|�l��cw-�AŎF�ۃ��M��t�&s�!y*�4�gkVsql���Հ�K�z��ۡ �j���;��UO�����0$"t��.��!˗sV�J�Vlo��ˠ����%�߬�v�,-���T�F���Y8I
J�U�Lvu��liB�� ���n)�����w�hgc�?����]�� �'��Ĩ��c��-9�!;��"����3_�ߊ���IwhϓVS����&$CL���F��ϭ��u>�&[B�`�wA��_��4�˜fB����6x,��-4[V�6�e�� ���ј�u�͊�J�P���-.�������>�u�7�� 7[���y��S��>^.$�<#��k)�J`�hY�j��A�ٱ�?d�����m�趱Y!�C��So'(�1h���>��|��nu�1-qں�=A��C�tڨ��ځ�+��wG�˥��ޓp }��PZ�s��切v8�2qɭkU�v`lE?G�l�5Q8���vd�\��ڂ�?�W�AW��uEJ�%�LM9Z�ӃS��~)ѝ�������0>��l����M�R,�E�l�_^��|O�r��᭧�:�H>���־�]�d��x	�?�$�u ]q��~����RuQn���,]��8�qx�����U�gS~�?��,�:�8�;���]�H])�P74\�{��ؔ����G����f�C<�1�rslڗ��WÝ%�����ӓO�m����-8'n��F(�=��a��Ɉ�Ε�:���=�&!V�j��� ����h��!p��qQ���=�7�KO?M%�����40ǏI1=�	���-�S��	���|u��LsO���,f����D�����{|��|���ne�N�~s�7�|M٨��y��f�(��!�R�1�I�M�!3���{^�Ez�����EGP�a`VJ��4�x���m~+TNRw����\L��L1�?�߄$-�HI�	,�}$��r)�8l&�ԋǻd�E��R�=��@�ET����ߩD�qxp�[,���ڼ��̋�)��)ѿ�9�gc�]�����S�^�x�	�PV�=�0�c�ެ�E�!��]:V��8�B�C"�v� �0`fsE�Q���p�p�C?����%=
���*�PK���+2���&����H���K\s���|.���}���.$QA��m�wbqF�ix�nKI_j*s��-��%J�ͨ�h�A>���:C)J=TfWD"�T�%��x��	��8U�7�D@��,�����g���J��
m�:��km�`���QjLj��s9Z�=$�kA6� \����f�����!;�0�W�"�|��u��?p�35�t�[���2�nQM4�dTz�><|D|�G����6��q��a��~�X������m2�&����ܸ�h����vڜ]���܃ͼ��Vʮ��#�%�
HZ��>�5(0�����He��#��8W�V��Rh�w�6���*��޽.�0���^z�]��M�bX)�7�3 �{�׏͢M˘�6q̆����|�Y�'3���"9WlZ� _6�������Ó,���M�߾�H��`�v��@���t!����*��c�`a�F)�n��|j+�`cN��� �R��G?�,*J��T��Ѹ�ڹraB��eS�ttR�ˆa����l���
�0�����ֺT�"�+���ƭ	�A�47�iAĜ�v��I��ͱ���QN���m��������T(u!�ǿB�{���c�J��xB��|xj�R_�����~��Uߜ���̗u���v�w��]�[�Rh:N
-f������$�s&��h����I�gE���A�jF�oQŌ�Eյ���y�^$�X9�rlc�Pl߰���R��C�K* ��W�A������{�Fyg��v��_�+X���7:f�˻�e��7D�n���]�eb��m�w��:�ϳT_�O��43f�������`H��󕑰��"m2Y�]�.&@,#���D4�Ah�w�j��LY=�����ҵ�V*$Ӊ:��d�g�)��VxD����6���?H�J�����3��_8���u�k��?�.��՝�e�mn����=l��V����T�����b�N�5�B���q����ȫ��"�V^έ��B�0g�m��Dؤ�/ ��<X�γ���+��p>}3H����ͽiJ�r	��D��A#}3J���o���<戃uЉ��}Z�<{��!$qS�$AVP,$oZh��L�9����%MGS��K�v����BԸ�f\���f5��:yV�`f,_&�+�r|�X�$�'�'�ޢ�������#qu�Գ#�6C5נS&��i-���z���:���u'�V�+�!��/|hzs&�5>�ygw3���@�@c�Qg>��yτ�����"nJ�o��Z ��BAb��A��іr��>�����	�A/:��z�a7e�9�%����
���Z��S{�@{�pp���a�\КZ�B�!��d�O�c�	\J4qk�fSWx����(5łt�2y�F�����%���/r��@�L�@}`�=Co�ri�d�Z���!{B�� 7?l�]��C���.�aa�%��95d7��H��臟��?H����o�:�˦�����s*����Hi��*۲�ߦT��>�E�~_�� �����u�ZD�N��ip����
��e{tb�``�Z�kP��V��O��+�<�p�8Ԝ�6_�΃���[q�#�)�������2 ��˸h��"���u_��x��K)�`l�V��Ik'{
F+F쿥��rR$�<�1�%%�~C����H͡
�ŷ+�A�i�`6�u��Z弉lJ�V�I~�N��Uoe~ ��\�� 	��E�4P������ ���`�kČ(���G�Λ=���[0�3!k����h7b�p��A,���ǀ�7K�D�nE��՟rl�p�A�[�'�6��"��/,,�N��b:�^�<���\]��Y�����)i��-&�=��G��#a������9�C�|0��' �Y����~6Dx��/ ['����+;q��K����vDi�RVv��W�
w�u��^	I�`Q3`��mz���gy/��bK�	�;+��'�m�]�5��"��fQCs�޳�M۲�J<��F���7�Q�|j�Iɒ�G�r�,��&&�%˟����cks���:���d�Y S'����~���*��j��\$�RIUeu*H����u^ߛ,}`�V (F�SB=!#A���0�	�&ZF`�:%��`=��gq�$ j���n�U�O������{��)$�^�o?Ы��@?ƶ��?�a�x�U�$mb#������J4|y�\q�9B���᳻x��EU�{<�]#LN��1�
"��a�-������w��2���C�%k!C�&g�ٌ@��OR^��z�,P�q?����L���=0=GE�z`�"|i�~n�@�$܂�����g�]��)5�Z�Q��lԦqfc�n�@�ϟ��;&BY �ɲ����LH�Wa�,g���ۤ�4[�O/�d|QV�=�U��^dЏ7lЂ��jԸ��bId79C��5_�𐷿?s�~1JM%C_$I�%PhV�&k�P3���4�+�G�:ie Bw�%U�F݅���Y�"]b�O�/=�-|� ˄������D'�`~�.Q �Ox1m�3�A�.cm�� �H|�}��jr�-G�
�@�L���r[*��=t��	���j�uW�%S�ξنh��̩�,H��u"���?a�^*�X��6����O�hU}|gN��I��y������&�E7�h"��[��=�~�j�(�d_�4 _Ğ�L�>�k1�A��R�Ԣͣ{x����������j�-���"����gab��^6S)�,�$���>���?	�����_l�qfj�����J{�f<���|l��s���O`6�F��
@!T�x[��JQ��&�<���.'�YFk<A�v#���������~U��Q�4+]�����c)j�.�ܼ���-VA_R������$0&D� <������%\ @�p�bi�����x�
�o*<�C��Jw����ZQa���Q��
Ǳ���ʡN�&p���ڰ�09=�\������U�Ah�ˀU�?�`�6��\�c���h��qw��Z}O\���'�ۍZ����@r��|�|d~��iq�uh3���*�����j��=�+��n9~�TS"�i Q)�b^k9^}In�����Iw�?��ue��b�`֘F�wˊD�o6����������K��0�L1&�zRQ^N$�ɺVڼ�I\C�����w���TYԍɋ�K��aZ�N%sd�\�
��L��e��Z�������~�+��'�"�!}8Z�Y����R���Y���[ݽ��l�h��*a�&��	|�}F�G�g�M��y�LR�G"}р�6�a	����)��<R�6�Ӂ1|L�3Wx"�@_���g�a��4\�0��(,��0�oɇ��sZؘ�������R�@N��xK�Kзf�~��!��l�w&Ҏ��iN�)�$m�8�����k*wˎ����YA�a�*�b3�ݗ��b��T��ԋ�m6��L��h���9�Fco�%�����4s��X�2��ڿ�����o�I��M��z��˕sQ���OT�]ύ�{k���ek��߾��n��և��E�	�Y�>س��?�d�o|z��,���ae��v���%Yjz.�tT�
�_C�����D
-�"�4b���]A��Br6:'5��}���+#�����˯���dH���p��3)2���~��L�]o���r�ˆY���-kJ�}iŒ7�;h���a��p�y}�K��Ԕ��q���l�C�a5�Ʋ�U)�j(B_�IU{\���J�E��q�:�����#���v���G��p�����b<a7H?��3����e�ԥ�~�H�F��Y�xN�Y� p�e86��~��Jb~�o�2�k@�Ϻ2���ړ����j21��SV�n�s._��g��D�IM�����y>^�qL0��wP�U*�HWI���GC��J�&�lB"�U:a@[R�Yq1��l;�b�'b�b�}O�����mA�y�l�+ <j�t�z�H��ϕb�ua�)��y�!�h8�;O[ ��A�ԥ��+��/�� o'��zLY�J��hZ�Re#�/��o���c��Y4Ɋk%���p���������R�>�ߒ�HӢ`<w�����@���
�El���uN�.�z�r���/���7۲J8���hPXwVm�U�+-��^n.oq���<1=��6I��	K,�Vt?�͏)3�[a�x�͐�z�U._r�7dQ�@��R�{dW�겷�f�E����@����Y�6
�_-�X?Zl9��]�N�x��2��j�lR�N<�F����}��'�5Is��D� l��Ұ������kT@�I�ìl�kH4Yq=���jFӳd�fw�c��?�	�(�곶�r��oˁ��9��U�򚀭C��+o����e0t�|�����4�Y`�&b�q1tcW{	�{ �n����Ai��"�L�A��ofP��l��5���RC.N�c��:���D��e�I���� r-�fi����a���27mʣ���WCȩ'-���p9��j�|ƳCz��=F�i���*,�@�ֹ��f�Fy���" c�JZU+J�،|��2��X�ejI�r�����\C�V�+���Op��lnZ���8��Z�>�Y\}I��AI�2+��|5�.��T�"���1��3K���/S���� \��'��� _b��,�^Oq�����7�ˆ2�1�^��j�y��>f}���2���2r�3��gbJ�S�����$���-z��4��`����Cc�9Ѐ^��ʙi�hb��yv��m���h�*(,(�T��N}2�ZI��Wͷb�I(���ٌI�@0�$)�9�����"H#�L�y=OHil��}��'MP_�z�z�T�ẋ&�d�c(~h���'/df�R~U�/ SK��&�x��ŀ�`�`����7G�9�Po� ���R�$����l%�7}���H`u����=���%T��2�Fs��O%�	|0^[�s��\�5�m�Y<DBo1Y��$(]J] %�\���b�$9���	&c���̇�]Tù�uȊ��i$���Mb���oV߈Pi�Ë�u[�qy&J �i�y�8�UP���I�����T'%N��Q��*�!�ʑ�;�PvˮvMݚ�_��ĥh�-Z��,FD�W����K�+�' ����ZhB�?�{M>�����.��ޯH��ך�Qᯥ���4�:A�o\f mw,�0��j��4�#��WU�T��R^bЀ��QiԌ�� ~R9ӏ�2��mkc����~[�w��C��.�V���[CY���B9ys����<�ڄm"����-�q�GN�I!�k�<6�����i�Ֆp��#����H;ο"���a,�I�8x�������i_NT��R�ߍ�3�bo`�m	0��N�
DtLǟ�^X�O.��١��\���L��8�&����z����_��O���k�?ş�.x���L5�&x&��}4亼�=7�%�SvK�]]P�w��ܝV�Zz�er$���K\�E�(;OSp�>~%;7��?�S'x�c�s��o�˃��w0t��z%31�+�yiY��T��/Y�~�>�੦M�8L5ݜX4�5�I�6}�ΰ��]��`6*������MœO�F�kڝ9��ykD�p�.}g�{�q���^j%pX�XA1V�WN���� @`
���O��)MP;�\�3eI+�v����Xd�̬W���x����Gm�,���>'���k	���J�^�+1p?��X^��@Mp��iIJ�;s
2`�IM�/F�Q���Ïi��[ vN1*P������Mѣ�6z�EO�Ļp�������Ҧ%�zp�$���5�5���ū{�|�R(L�+Oh�*�\!?U�Y��/o=��D
�P�sX���|x��iak��w���>��#�)c$8�>�w���ލ�	�!���ؑS���r(�
Q�'lQ����nQڬ@G`6�8dj�>�B���6�-P�;`%�:������h����'�d�+z���"����S��+[)����0���7"P&�z��Q�c���F9���g%G0��pd<�[���_퐥KZmW�T�%���9Ny��ִ�:��=)���M���#dX$2/'x���z�=�1v�_T#Y��S
��孰�㇈ό?���R�`���W�V�q�r[G�JF����3��Ua9�1��;��ETx%��0��]D�+r�8�y��R3K����m�/�:����Ŧ���x�KUT��0Ι8�x:x��^�|$��CW����zoyN @Z�y���L�����h���)%�%{�)פK	ų(�/Ѽ�ƥI9�N��}�q�)aEBGw�)�S����y��'Z���	�\kڝ���T���R_y�2��i���a�h� �6�����ŭ��m���gs ����{ECc�cV�i���k#�����^�|�#�)?Ph�)n�=cR>�l�\���ӏ_+�<�&����8g����I��&+|:[9,|k�֛j�Q�rԿ��t��r��=�sp[
�y}�#���ܐem,��3J6�b`2cBݓ �ΞUBڳ���T0Ԍ|��zJ0����	�L{���M��˼����gz<`mOd=h�F�M�
e����@�f�<-D��&jN�>hi����Ru��@�(2��4�V�T�:<n����=�r���3Km�cS$%U'����td�ʬO���D3q��D�]x�-��8�߀O��Aw��=`�k�s��5�J�s��׾߳$%��-�&Վ:������'��5%<q�reCw�g����ꢸ�e|�թ����iDV�\��Wmo�0�<��ڧdA�ݑf^�!73"9���<����!�&��5RDO3>�����]�#�.����fX�zj��o�8b��
c�����.��Ƅ�|j�Sm5����Vn&`H"�Y�O�n��B�8����%�ygfg��+>�.��	 ����̃<l�
Ϋi����5 �L���qASϽ�_�����<�Uj�4�Ǥ1������_��<q%��'!�q��W@���4
o"=�u��
�ț�G�[�����-���7�v����^D�R��;y�h���
G4�����xY��RW���D��R�㑦�Tշ_<iOo��Aʀw�B���	�SY�Y�8ǲ>�����~����P��������p~���C��ńN�6� ��7�(@�>����[.q��XY1�
�̪E1�U�Y/7�K�2��+��e�-�m�G��o��X��G営�:8J$ �i�Q�k�{� g��O��:w�#K��?�OO�������Mr�Y��?{�;�t�����/��A����d�Ǟ�fW�N���\���_9\�����[��vI�&�כ���)��NG2�Ⲉ�:�-�u�*�v�i2����R����5�&�����3�y�(v��8���`����e���u�A$�b�7��<�~/��j&��wv�!�	�3�v�&�^�m�LMx(mm�\S�.E���g�y�v9��?�c)�^F(r�{)ĥ��$�������=kQH�pR�֘{f�f�빜�0D�(ϓ���'aO���/F���q�w��cU�X��\
�R���(v�9��%r����Zw_Y������w�������J9�{���:A�b*U�{��t��m���uE��ϝ/+���b��
T���+�:�7H��j�)�8�9|_+��d����4�C�	Z��[�A���	�`���|N���@����	�0��̔}җ�� >J�:Vkm�Ų%�Lg
B~�i�%.m�&����K�kǆ�5P&��m���(4�'%�s�U�E��//�Yy27!���d���F���{����'i%�-7:�m�N²/[iz�v��z��Z
}�M,�f���$������4D�vq�M�J�7��{qf�r�	��@��6N�����262V���"+�X�j�Q�{3N&m�^��lC3��K���A|T!�A�/���s�m�D�U]���Տ�R�C�ئ!qҒ����sw��3 ����������@����&s���R�z}U��t��n8h��,;��%�0�cN���>G�l�>?&��=�GUiR��1�`�}�"�uk�t�f4ձZ�m0���B6�V�t�
�NS�0��@�
�����I;`W�|��ԓ�`{�*���O��Ht#��Oc�}/P(�mg�5ǆ�Vl�e�|�&�����`��W�5 &�H_v�ЫBc���[���+��U���hL�Ǎ=~Rܾ�t��M/EX���
�x�0�-�v��z��4�kؕq�~X�#�:�ƶ��ET[�,G�_~i/��J�,�jx�6���i����N��|���΂�3��(wi�6�������h�A	�+>ձ w�m�u�@�"�}��Q+�k7E?��x�)�d7��u��h�_K[��Gx����̤rĭ�v��J�Ȓɤ�~����-�H �����Ʋ�䆈�<e&Ct��������� �Q����#���=��7"��)�'_N!7���~�[� ��k��}Uw#���T2QK��w��%���-K1G��9l�\����\ht�A����Rf��Dr��2���%�iY|��(���n�]��4��%�̷҇W39��Գ `G,�Yp�4]�%�� ,r���t�-����;�	�,����渪�(�㶭���Z���F,�ϐ��&���I�R"������CV�S��qY$��+kׁ�7��ϐ�1~�|� �,?�qb]���Ş�7Hb�D�4�?���V����'���|KfoG��ί�m�������?���=���r�B(t�n/��*������)6�~y��Y1�+�14�7�W-��iZC�9�K�x��~�v�&�
�3xA��6?�>~ ���@�F�����f"m�LA�g�"a7c�vQ��k���y��^b�d�/"^1?�7~w�9���0�ʺ�4�q�pJ��.��L��#�#�UR�8���̉#X�"�	�a=2_7n�*�xO��������t\��_!�tQ
����W��X˭�SH�p�X��V:,���2)=���Z����)��9;,�>�-���]	Ⱦ�?�]>_"��; m���-���x0:+�O���P���'�|�@�s��E�/H����n�?��ݟ%�{w�ѳ_1�S��Ϗ;��KpDM���NǟL@i��s\ny �0`J�d�ڏ�P�Yb<����JGr	={��Ul��[kU'�z�9��*3Ф�ʌ;������w�T�����c^N����b�X�`cS��S�)
1!�;����G��Mnʊ����g�� ,�6�9�u^H�W��Q t��Q�[.|@
��k흫�H(�*�L�ٖ!E�r:?�{���O3�KJ�R�>�
�0�qD,c���y�D�� �ږ�VzWӓ��u�=	Q��=k7껞Ȩ���W���t޸)x��R��8�b�xi3[O��D�bx"���	/���9߾dC����:4�~h[���5u��`��[�kv�t��w	x�Ny�[��$y�aì#�����/�_
�k"OE-�Viͬl�C�V9�N�"�7�I��,�dk�:�? �Ds�+YQ��QU�z"����T��^��|;�EH����0!^\�HG�*�(v\���7�Úf>��V��yq������*t,(W��NU�b>����֗\��OF"���r�M�0V�^z1�8D����Y85w�g=���ڔ�g�b�|v�2?o�($A�,s�G'�lH���/���;i!.t�K^��D2n@��p��
��= ^�X�y90n(��4����J-E+j� �wj/$����},�ǣ2���H�9/�	[b��?����f�V=B�h�E:�E�U���U��]̪����A��
�D٤�"�EfBa���+)�_����^F* �3�}��~��c�R�"���5��.��7p�� ioI#����-�	�<�� |���q��W�l~m$�i=Ր�	Q� �Q�TS�r5=� �v��98��b���������s'���2�d��ۂ��웵��B6~:L�6��=ӟ6m?���#���JP5�����'��{`��>tl�}��jD/`:�,�E�:1���;��g]���7�^���h�eI�"��i~3d�xA��M�X+E%�bP����u��&<>c,8�7�-U��>zz���g�9r.�5��yx{��f����w�oOf�QF���M_��Y������}��Sa�~����v0�q[�ޔ������`�_���U�B�n�E�ϻ˽�����0���є���3��M��L*i��2J���Q����Z>�z8Vv!g�h���+�����W�ѩ���|�$�U��v�tSi�L1/aYV7=���r.Ӡөq���~A ���y�p[N�N�A�b+�OE����V�����ٗ�M�P�w�:�A��M��r��,ڵ�e�B�Y�\ǘ�r��7���q�F���j�|��6�ll�M�pR�`�e3|\�������_>�5���h�&z�q�W�A͛Tg������ M�}�C�^��S�j*Q�D�+�T19���N�Ro��U���P�|�Z�n+��$ƾY)C��� \#eEN7�����XK����Zx<_ipV�qX���J>^c2Ee�N�r�����&Xx~F�w:���
W�G���.�r\��t��/̠�n�IO4�DO�=��MY�b��gdsA<9�jڀ�ߘ���k�W;/u��_��� #�c\��S{�);S�7�T��/���#W��j}�ߛ]��N3�ד�;���	���^}Nφ��r}}�˳��!�dz��LȪ	�W�k�\n�tп9]����9zc��n��#��u�VxX��t�Pբt���؅£!64Q*Mۘ[�nq�¢77�0(�n����s���p�(�ۼ���$_}3��ti��Do�$���ȫ=g�|��bv4�~����Ӷ��O���kF�X@�|Ҷ
6ceX޶bN����uǀ:4�e�vSw�(v��%�^'u�E`���PB�M����]^�'s�f�.�|�qJ��p��EȤ[*b�q����~���B��?��+K�+��g��5q�n}�Ţ�;� �}
�Vc��,?� �q����<v.f��Q�FXU��F�w|D]��l�DD¶I93��j[��GFh�3ž����/
I��KB�'�⍪����R:*�a�3}:ӱ����2�<�wn�n8�R���=��
=tԣ���8d>3���H��}e�By�\c��Cex�DH����FbR23GG��^E����ucq�@���1.P�l1��3�bb*06�2_s���������E4C��*i��hQ��B�/���*�x0��RE�����u_n�qIR:�.mΓ.Ԏ�7�nt�ه�.�Z(9��uA�Ts}-�g�O��.�i7Nf$��Vx�Ɖ�;���8�+�+����I�c��q�<��i6�^�r�NGkp�A.@��U���6ϐ޺�މ��K��&��z��|X`�܅�N���u,����������y@�!x�"���q��������tK-4�� �HHwi7���!w�s͘�V�QE�:r�s�q��kN�5��&�6�<D�*�[��0�r�|uP���<@��6aC�e��R]��}��;�t���&;K���� �:H�Xط��X!4r�V��ݕ&)PPM5���1����gʂ��e6�nCx���Y:K��ɗ�f�W]7l.�P3�D���|U2���b��
+���ݖ�b`Fw��Hw"k@��_<���l��C]�.2tI���Z���6)8����O�s?)�$a������t�is����$�<yu=|?5�5�:�w�oI��}guI� ߕ�����tF���m>9_���X�=gJ��^����΃	X���Y�P�2�bP����\�s8R�d@�15���}YH���n��,g���.E��>d�>�4�d��Q�/\�x>B�\5���'����~��S=���	pD��<1�A�Q�F.�wB���:1h�x`��pJ&Q��16�>�"�bu� aS�s��������u��1����b��d�M���	�-U���9P@e�<U�����~A3����n�Ct/I�#�� �+��%�r�4R3K���[;��2un4�a;܄�+�˶���b2P�r�u�#2!#Ð�
�b������T5O��g�'��������>&ss�>E�x�4�Č`��20��GDV(�xYp��XŪ���94��.�#N�/��	= �:�#�Է�M���!9Su!ւ�Qk�/�5�V��A밌;�~���Ah������&�ޖ4�4�����]�W,~D0�X�N �����E�����=HEz�F�t�,�<r����FqQ�@�����7���g1u�=[dE>�q1��6���$�5�������|?�׫k�G�L0��X�]�]\�)��X�t"�X8�ۦ���:#�+O8U�}��G��d�Ua�i7����%/5�!Q�����Y�0�.)gr\g�,�S���,���Z.�{��xX���TY�����r�����!�(��%����-9�y���.=�&f�)�-�.�q�dOߧX�P��O��ҡ���B����������Hl@r���_܋V���IO�ٵ'a����@�A#c���U�d��ωI,П��Ͽ��K{�<��:p*N�\��	��HHÍ�0Q�P�� ���÷)^�9lj^@.T�ge�C��?�7��ԛ��Z�"#�\,h7�?��^�(��ի�k:^�l�%-��y�!A��;�7+�*z��¬"[�E::��dJ��t�-8jN�c|�/��?YǒL��͖9����R���gՔd�ϟ�� }�y��+�Ü���v�u 2F��q�s�:Yc�a�aNwz��Dr����0��ɒu�h�Nɇ�zq�f䩃L�wǧ����kw�`��,��^��.�	�.��q���etKv��Sʾ��˴|�B{兘6�+�Wl�y����� �ܦ�T�<s�k����+h�aT�rv�v�S׳��܎����A�Q�:�����6��\B�>��.���1�wH�i�a(�>sg
�]�/��;��DՏP�_������CXAH>%���2���x=YB�޳$7���gU`�f���) x���������07��� Bq�;)���!���F0�?����#9_��T�`�\6�P-��ϵ�/�'��'�H�cn"��Nx�� ����'~L��M���G��ʹ�5���"?�Ӟ)�5M�dJn��h?p#����ཱ�G%r�W{A��H� �7tN�Bxb���=��k���{�o��ܲ��{���6����]�������d�E�筲�n��u�Tß�z�𨧅ػ�)��K�/�evV��H�L�ɽM9��_$�b-�r�*W4����Yyg�U{�cC!*�G������u�7P<J�^��eA�M!��iw�('��cR}L�r�$F�연���m�+�r��5������/�$���Z2r&U`���b��B*Rs��x�(�_g3�J��of�TB2�}�"���S��nG���?� ��3w�M�u�LC��1<�D��]��� �=���bt�	�n�>Ɛ�&�a@C�ã�ʔ*U?�N���g��s�K�A3@Ψ�3-7Hλ�ŸH�r�����ئx�0�u&y7󟍥e�ò�&G, ��^u���w�8�e��}�i�K�����-����*�T�y�A�ǎ
���fs�X��� ��#��yK�>w����j�-��_x}�������^�:��+�01�>Y�6M(D9��+W��?�<����9�4^N�+�K����ޚ�mj�h��˓8��TN����uG^(N�㬌$Ytu�9|<�wOI�N	}��$Ű<�Z�Zu��2䲌JC.��+�F�b�|r��վ	��[1*G��Gk�`�-����N_�����4�O5��g]�?�ce�HI髊	��:�C2|Ǭ�l���O	�ٶ������r���לGge�Fi�T�|BgXZ���#�������:b&Q���eN�H�]P�;.���4���=K<"Q��I�nU�ȸ1��@$�8��3[d��ig�1
�E��Es�:�O���-T�0�%�@���RǵN��|R*�:��t˜ �,ִ�	�1�D*�����x�cmh��K����,�m�=���Ш�!��S<��G�&���j��RL����a� n��S0�Uc���%�7fZ��9���2b�.�b�u�/A�u)�
���D�My����(�N���a�V���fq�5&�����hf�9^�@�x��/���A!��	���=�����i�/�TM�=�,9�4?�J����rնGVA��))B����7&.��z��/��)�+kXrjo���c��'�,��(�8M?������n
���d!����4��/O\�B�F�亄���k������t���0�4 Ͳđ,7�چ@��t�v@?-�:��@<N�= V�c�F��vN�|��qr���;�2�&}�ӳP�<s��M���dfo{x�e�̧T�#=-�>mEZ7"D[��|�d�[�Ż濐�w���M��[��q�,����_�VL�t	���w��V�*��������{���L���^�Δ��vp�PAbz��=>:ER��"g;�_# Ȇ����G:`��%���02>B01@.c�J)��c���/�T`���:����K��ٹ�]V�ˤ5K��\�y��k��� ��C���I&�(�Lg]�I��>���[ބ�yUy.�=�Y��%K�[8�֚������	(�E�)�o�Ӟq>��a��N �@�}p�8Y�"zL�����[�&">�����22�HƨZ�g��SVz��;�d7����˧��TuCa�;ad����Q�x8�l�Fz����RE�_���-]wHe��]%��>�F�޷k�0o�J�2��6X���s{�Q6fy��SkRG�6�㬋K٣��E1di���E|�����r����0k��!r+�;r������r�mY���K��Ö(����=�;�e7�V��$��eA��ζS
&�+A��Y<M�9��G���C�铐?��_�%�����`f��K������q\Ub��*<boVxH0���e��{�����)�P����d=�����Й�J�N�]׆���X�}ミ�I��_Y�w���1���kM�������!�o��\��A6�lD��p�"	�T��V�ߛ���o޿�X�e�/��#{&�$$�W�v���16`2��q�B��BU �s�'mD��Yh��	���k�f�Du%�=#� YM`����n��WiP�}���]���6d֬믈��T�ye�ye�����Z��l�LH��A@d/����8��%p��糺��
pR&��d���o��<1,wh'Rf���]�Cz!�'-+�}��d��s�=�s待�l��i��*���f9g�zV�L���|M��N��YPQ�S�ެ���|r�Z��Y��e������Jo��&���M��!!�v�I�<������<��S����M���#�7�K��~����;*o�T�eZr�Pb�|qv��l,�>��%�����eK��ڻ�⮴.� o�̝f�5��e^�ܒ���F��^<�T73���{v�%ԏ��p��)<@�$6= ��V���THt���'%�mər~ gQ�z�x=�g] x��5g9sw��.|AjĈ�2}&��BA��gWg�C /k��ōRa^��;QEq9��]o�@7��I��i�D�Z:���O�T�C��0�DX��m/C&���/�s5���C��MD(����r�Clf���Իd?ÒӴ��cg��#p�n�� �H���X�|�CaH������Lx:�LD�@&�p����ѝ��VT$�?��p�i�`s�:�;*����/�c��<x4���ҭ�^�_��k�k��(�"&�t�R
C�����|D�
�J�@�i
߳��bO��6���H���
s�/}t{����R����G�ב�%u?�g[�ԛ1ч˖�YޱwF������oU��4[S�9��@��U�����0�������i�-<�/=u���]���W���=7�!����66_�G��g�i8oz�h*�#�Ε}�xT�N��[P�M2<�L���c�m��`=�����Tj[w���g!z&������¤#�LCOvc�m?J��v��Bms�'��WF���N���� j	�X�k��2�XB��Vy�Օ���*��\f+T��#P#�&�u�C�5�m��nĤ,i�.]v� )�-	ߎ�F��j� 8
�k�9�U�畖B�������3;L�%Q3���`=.��̋ŧ`�MtpZ��td�xj���v� 4�׿�l�;��^�u�d`����Ī����?��L�rb�~�'�s��(;��"�mq�nř�"Oq���	dw!�й�KŸy�]~�%�+/z���gv
�{&�;Pj�gE�,3�,x�"ۏ/���@�0u	��󖐟WA��?���Di��t��V�-�R���k�!{+�+y��q�S��D��p� � bK�T�(�\@�Az�����>g��n��J�?_�ShQ��:��d��K�u�tw��rT��\2��V�� ��\h�+I�쵾P�%	�΢�EdII#=qJ=H����>�Vf�9��[�:Ya0���w%G�r�M룒O2$F�gz�+�
iTI': t�@�#9H��qe�Z�F��l�cP��5��3L i'�؉�
耄,Xg�#��;����K����k;Î*j^y�! �v�.������W���S����_ޒgJ]�Q�/r��R��H(+�i��������#�eDV��JctO	-׋i�������- �����D	��W+��Em�jP�(xҭ�NlA��C�� �~�rgu:�絥1�2ī�sB���>D�#���Sִ&{:�p��̕����I���8�?�ݑ�j3���_Ҽ?�� ���Z��Ŷ����sa�:��H.�Du��ٻ8>pm!����!�9.�[�0�}K�̿=�� 4��W��mC�����^�M���}3[lX07�"�@h4�V���6���Ň��x-�f�;�)����*O�1cP��N��;4{Tb�e�@�5��h�� �9��Ԡ)t�+Ub�:�C��F�t	�k��d�l�77�]�IDEB�|��� S`�D��ʲᣡ\��~-�e>���Dr-2���[%��>�4�ݏ$L9(r�+�� M�^4`��д�Xg�|2���9]�$qQӜ���O�-0�������Aߦ��x׮�븲N���W�e�%)D[�q2}߆@K1\�?J ��ͬ�K�X�>.3xh_q<�&�������uA��K��vיK�����j�A��@�?rQ��&z��>d0���}��Z��῾�.:L�̧I˴mj)I����M�z�Ԏ�X�b@)��ᬸ���~�`a�����n�>��qj����i��	̪S1/�:���xZ]P�V8������S�Z�?Tm��u��C����i5L�Z��;��'^DuzWO��~��R3W��l�����2�YU2��1Ts��j.d�G�{�a`��q�f�f��0�Q�����q�u!3י���'��GnL�z�L�aڞ>Q���G�U�鍬�G��-���d�	ld��=��Du-ӧa�p��4p��Epj��w���[
?;:SN*�" �/^F�UK�/2��`+��I�"Ϣ���v��r�{��|DBv$!5J��l0�v6�O�Ӝ�x@N��r�{� ��Sb��� mx(,�ܼ��:(f~�VJ�&o&U���2C�nقl��7sy&}����׭kn��6����0�1�X�M�����F04-L���)�$���%���a�7WἫ�-R^ )�O�3u��9a�t��#��/��(v�b�j/��\F\[Z��J?eÏAfQѠ�,=��_tLA!��� �ѧ��,I�sɭ</ ��j�|�6��2�^�� 	�5�ՋI�8�uE2HNO:\�~W����W�w:�}��S*X����^hd�8�l��p�9�#	�=U������v����iR�����@�+'$��3��"��k�F��MD��X��x�:�
�X�f<�<�����IU���C�CE���Ӈ���@
��_�"�C�t�>��%!�;�N�<@ѫ��z��*�����R���N���?��P8Y\�d��Q��F��a��s]�E"b�������P3^͛::ඓ(~�ڍoF.�M�����8_K�U�y�˛q������BJ�0�Aw*xQ�o��cr��)"щ����fm�U���`Y�R<��䫘t�P:O"���1�֦>���q�>���1�5HZ�̢O�}�2�=�>+��Wbuӵ��&^��Vp0���#��6L�ͭ#&�	t6&��I�����r[�����AA�)�dH	�j��S������J�z�S��?I<MŔ���H�
E��|�q�q����i�v7Y ��V��7l��bu�� �P�w�F �����ͤ�e�� 	��7IBճ硠$]��Cݑ{�D�I�NB��� ����$XF�k��L ��Ii���>�
��[}@~g��Հr��`�[}��?�(����I;��eq*X6�H��.!�����ѳ��A��u�e�+�#�mw��_k��9gQ�����6Bu��?�P���ƌ�HW�i�W�"�r��ʀ�O��!��e���!������*FP��!!1��U����CUj��'�d���������E��E��C�����"O���#�j�G�n��Nꁵ����2���Wc3��X�g�۷��+�K�57���K)o�	#*� �`�!��������<{��V+�����'��=�~�A(9�y�&!�y��ǞLKk�h��������dfm(��.|��j|5�C�kӼ�D��Z�+q��Q��$ik���������o�42�1�x�J38(����V%r`��d���V��W=M��.�Ry�21=Z�1ȳ+�	�ς`�!����}�0H/�,r������;��Qf�8G�?�����`0�g��)`KN0J�ݢ�p{?�d������ʷ��D�ɇ���M
���`V�9�*�lG1N�jd)�{������������w)��ޠ�0�Q��Z+�â��IV_���1z�W��S���2�J�z,{�$-��"��q�Sd���Z��W�ci8�S^��k�d� �{a֮�&����kL"�y�T�d��O��T������ @ԃAr/p�S�A{�Q�[	���)������n�i]��$�4{�@�˸��n�n'�
�{�n��b�����	F5�9��a�ͻ�������<M^J�����˰��<^��R7��u<�U]���<�%i2hB_�}��i�c�l����^OMS�J���wY8	%�*hn�gy%$�4��žUq*��p�µ3���6B�b��l����QʣCٟ߿n�;�7� h_�S�f�]�}�G�d�T������Ω�3�h �����,��X�؜��&�{J���X�5���a����W`�2�&~"	0Ck8)� ��ugs���iGҌ�n���@�9[`5˯ڄ��cU�)��O_���c	���"-��W�7��zt������	H��������N���YI�)�����N�<����+W����C��w!��
���u��"�u� �kk�+�nC��xF��I���0'�����F���[�Q��@"��U:n3T6���DA��]Hʐ�ʧ�H4W̒0���~ &�?��������4�9v.�(�fԜ���"��kz;fp����{e���֐�1�nI����[e�|�$�ߔ��%����ٗ��������v�3�E�!�=zc`]H�W��yr�.�*7��hU��h�������u��M�Ċ�ƹԪp��/�>�7�F��s�b�����5@�� c�q�R����}k���,��k����s�����n��YyɴU�s�.����Y8�f������>�)L:�vbƄ�r�>�*r�=��
zv�A�n~����A�4�|�P6=f@��T)��ƨZ@���/�������~�|Z��Z2�X�JOf��IF� C����͎�|���C��� ߭��M��(]EoX`$�~gs%���dX��3D��%6�2��ـP7ur?|P�D�Qg�u�_����jE�I�]��P4h8̪8Uo��e0P�js�B?��XV"\N�%��.��ߗs�3{Wiyz(���}R]vϜk囸��/�a��T���amR$��3R�]�8"̻ϰ�m�e��P�Ӂ��J����9�t2�������Ŭ՜c����aW���i,�G�n��gSl%�MEa-�2�����ɠ�G����s+2�*�7��=/so(u�8	ū �x��ͮi�~�Ӄߘ`}�j�Y�'��:�m�(�DH7p{�&� �,�T %r8{'x�Nh�3(��>�%���9vX�Lcj0g)D�{���U��d���E,�D_��:�l���u^L�q�B��_͛D{�����FS�7_�7�J�E�w�V\v~H�
�P�W"�O��x@�&��ft�'Z�s(��zJZ�m~�"��1�/[�|�cF�+;������"X�������Hҧ0�oˊү���n���6��c(�҉U�_��9N��F�ڊH���d���}�v#J��O?��*v�Ν�#DF��e�5�C�F$����W�,#�W'�<)!�p�Ҁ�W�����~�p��L��τ!�W�^�R���e�,Gx��e)SƮ�Γ�{ڭ��#U�nn�l�Y'ͭ���\�V͖Q1�4;3@��p&{�9��c�m�������Bp��ۙ���H�<�z���"i�%*�yD?D��qnme�zZw)��	5W��'��Eeh��P껹�uԣ$I��G�u���6w2�d@	�?��C��{f�jL!JQ�����}����l������_Fi��FNHA� ��1LW�d[� 
8j�����y�3�u�T����ȳkڈ���+�p��b��kmz/@��c4<�!�er�(g�ڻ̄�b�Ԃ���̥�em�X#؜������Є*����	����rqjr�\�2�!.�`:ͮ�V˭�/8�\4�N���@��;��|T}Ҵ�hfI�E�\E��9�?�YG-�/=�"�r���)�XM�ί�$�&�)�������-wy�y?O��)�#�A��R�b�y�,ʩ�˒�b�(�8�Ƹ�h/)x�V������~���\+������.�܊M�6�I��R�	�7�D����p�L����	��|��A<S`���w�D�� ��zЂe��/����Dƣ�r��/�)���k:F�/��/������*a<�n�?�}gA��U7�SVgt�M��0��HVO�D�$�7,=�����N�v��u"Iظ�J�t��}��	�� X�S�}'�2|.�\���L��G�WVGCw,�ͥ,$o1I2��I�7����~)�$���\�_��JϑQ���L����<x$��.Yf���AtQ�Gx�4\k�.�
��F�)Vʆ9�p�H�[]�����Y7N��#��p�Iv|�6�"n��u!S�Ǝ#���^{2�.濎���-c�����w1YQ�oe-O����^ђ�X+����7������h;��9�9�=:�@��tċp���
~Jk��?��h���s���#l��Y��9�=a�IK�X����B*��p;]�޻[�6�~R��a��3�t�a{��Fql:\�<g�a�$��T�Bj�� �W�-�E��3ð���'�p2O��3�Y�a�=��Yj�i���B3?�Q����,����rX�56VT<�C��,Q�JՔ����ީ�T�3D��~W���s�n� GSzj�A"3�]Q>=�O�@a?e�nV���2����a�������eNi����O4�H[���j��(=�I��v���Wl�/�/K3��G�[8U�t�Il.0J�_Q�8`i�3�|�Hv#1�B�v\�ěk�P�Ɨ���Z�l�']��%4����h&;���j#�B6a]\#h4ϼ�B�O��uk|�0�aD&�az;.j�<A�2>z0�%G�B�xǍӦ��2(��9��ՏqĴ<8^���Č$�JXB~�m�ɫIq�|$�k�j�h����E��T�?2ɣ�G8��z<��%���m6�g/���GSe�Y��,Q{f��zY��;wB����W�6�K'e��7��ζ�)f`G�	}��!��<(�{*��Q��N���xK��a��������Xـ�g��<����M�5���c�b(��5�"T�E�<�����"�d^���� F�ې�n#Y��.�ֈ���� +2�wG�u�,��L.r)cH_����EӜ7�DX�l#�����F롗Hc�7O�Y\��N���w��j���Ў�t(K�����	o��?B�c[��	��{c���@h	����L�fM i�/j���W+G��Y����_4�ʐ��h�ƾ�[�k2>��m~��l IQ���<�COo�dkOmW��6I'<�-z�  �d�.azp(�RUW��p��
ԣJ���VI�k�:ٸ���7n�L'��<�V-03�t�T������VR�a�����6T�tʀ3�������*�I�ӄ��cN�!��#+ g�q?���(	�� B�vEO��bǜ� {�𮵯~� ����S��P�G��^�$���YJ��~�*��۞�򬜊ˀ8�!�.D'�"����5Xv�ʟn�f�W�\���B���f���t���i��Ca
��0��p	M3O��ʵ���
 ��!{�����m'�a's$��{mvuC�>�R���#V�,o��# 
���n]Pgh_F�,#���w;���n�o �Oҽ��A�\D0އ	7�:��o�#���+.�X:mJ�d:��vRfp��zx�'t}��ImĘ�W^�3*C� �'F�6��k˽�"�	�D[�e5����\��R85~Q��$!w��j������9����6Ž0Rs���ZH�qY�0H�J��&A~�!�!&*���CRW�g�C� |��<�U���j�Z�pW��(hw�>��V��rH�`�*T$%���5��F���dh�=,'i�f��Í��8�~?Z;ɮ�F�'�i�07����j�α�&}0�W��!�?�S�r,�YA|�k�G�Lܴ ͇�u;��?ڰ�*��&ӚS�Q�l;�
<��Xh�ҁ�9���.�7Z��;]�a:aN��@��@M�\~zya�Q��Ig{�7+���!�[Si�o��9LZ}��Z��N�tc��(����T�٦8!�Y�ɉьDe�+�� �����J�mKRF̳N�W��h6���!�y�d�7���Nf$���G/@TH�x�y�<�A�R���őv���ލI$ϒ��/��,n+D�h��nb&����&����=�������2X���Y�mq��nǐJPAc�6vj]����N0��ymL�+y���j Z��i$s��G���t�C��#v�&5d���:W�d'ګmG�Z��?���u�d�o��4>��v�r�V˘��:�N���)?V�o|�-4�Pg3�C����W�Ob�����(]��N<�$��@���}�T�pIg���1�{|��m��$3g�'���(a�Z'X#%h�b��c�g�+P`#O.e(X�4�|l���N��:��s~u�V�h�܎q�A�{�ꍵ)��v-�p��~]��/����ac�=���7����/�8(���!h��BV�,)��./��E��}�7={����7Dک��m�2�u��ym�&��uZ5���h�^�b�Z�AU_-�[e��4 �\c��~�C�.�W�ƍn�D�sT<�`���n��`S~����)���$���b��&>�Yc�R�L�b��*tۺ�2s�����dYBkץs-"�g�i�V�\�l�O[�.�s� �V���c{]��j waI�F~,o[���h6������`�8�K�
7�6�j7���N�2Rm��f���}�i%h�܁��ɼDU� ^Џ��N��aWŧ�n�,�ǽ���5
����._�xa�B@��Fk�^�#�	�w�j�i|������KL!�t�ÎuI�H����,��BN ��Uzstm�A��(�w�������A�:�\�4Nd�YD�D��N��y�/�c��j����E�g���ndt��ۚƬ�C77�J���Ae�M��,?*)��eY��t�#�Z�=w���&I�z٭C��`�ɡ# �ݵ�&���E�x�
�r�qӟ�➖<�k:w��mnۇ��JYB-�g��O�����l��B���m>��
��bt�O��i>BU/�?-�s/�W�����D�+����*�I�M#T"���,:�)��%�b�Fύ��ן "Ve:j�;%��bM Q_e)�A�G$�,� U�8��_	��R�h���+ ��5�E�d��5[\�ٖ����x��)L�Jw�)o��_I�J��Q��m(Fa��e ��ڒ�xF4���q�:��OK���>��1ff�uT]h�۬��Z���߯V^�M�3F!��պɱj��_H��&Fe`R����J�׼���5m���ƀ�S�A_ν�'L��)�oW*^���vd4���Z�� &Þ)v�G���T��F�W�?�k�;Y�d�n�@�[j������0���3���P���lq���ȸ��љH�������C*K26)�`G��e�J��e�.h��T0���e',t�+�ղ�U�}���$�����=�, 0�S|o�H������FNX*	
���A�K�V�(��1��!�$���ZN�7����б�	�UX�Y��_�\�%����y���{�:|�v���9�xC�ֺQu+b�(u0@#�O/���Ke(|�C&�O��:3�y�j.ݫ*g?`�>��ۑf��ɓPq�O����_��#���Yx�|I���̥Z�+��J	@zj{��5�ȗ���ī��z�Q�0�B��"5��*���ݿxt�Zi���b\/|y_��"%�p��L�~T�[�P�.��z��R����͑eS�OU�N���ۄ(x��=�{ׅf�ݧ�.�P4R�M�0�q7Y|&V)/��k�Ǟ�'�\��͐R�z�q���xH��7x��d0��Bu�:=�嫋&u�*V���Q֢��,b�ܶ�+.y��G�>f/!}�ŵ�ʇ� �������#Y^�Oտ���яz׭����o"��Ģ8�]��U"���,�����!f|�]v�Jt<��� J�Q���v�)1��ZH�&�J��v�p��`��	�q<O�̰��>]8�-Z�-�_��~^)����2��J�AS�H�ĭ¹4n�>�:���!�Ĩ���f I����ր�Ӱm�'���1s��,a��K!�?�B&��SsA�֮���tqz�x�s��Z^����Jr ��Akg=$~ˆ&
b�`X`����cDUm�}w���e�4��Bг�_Ӹ���F��o�B�b�p���m
���::_`|��/(�Z�S��hnQ��Ș�W���y+*ĔsW���V����H	r �4����(��}B�k1��j�f�v6��У�a%�ЈK�U#���~�(�@�	�����B��G&�(݆�R�Ӧ� �V�'l�0{<SJ�}��W��,�K��v�����L�^�$��Z��
��tND�}�=�^ވфN��%�UO��7��[ �P	�]}|��q����%�A�{�@�6e�8�z��Tf���Dt�ꛡU'�`�F�'�ps�ũ��)�Q?ƌ��F^7����r���(��a�8qYD"���u��Y��?��4U4u5T�|�Q�6r�!��w��U �ňy���߽7��E ��\s��X9S�H�\:��{��|���]�'8�V8����o����#恖�reVm�=����VQS?��p�Hi�?;.(�S�����2��2�L֓���1$�r����p��\��!��9����׌��l�R�#q?J|&�C���)��6�R���7-�v�k�υ�@1�H�c��eX�o��\���T4�58�������k�t&��4��#��P���k�p�Z���a�S��
ۺ`�f����6�!�}����+��y5��VZ� wJ (���Ƕeƛ�(��a]Q>>�.����`��[k<�G�+��aS�M�]�Z��_ж���e=���hG�I��3f�]*>;���v��6__���/���9�WX:1���B�z��f� ��O����|Ǿ\%f�Y�R�~;�� г#�sː�x2)��֗>�*d�j6�#���l�Jm������I-��/��0β��f����W�������'U�2�wAx(ԝ`���o�#���4� ��MM�X��`#h���+ �Xf�c�%K�ރTx�2��ੱ���c��@�t9̍�SW�֣͌eJ-;�Q��=>HF�p���B�&�0芥�X1���%�2���A��q<}�?���}J�k�cSSh-���)�~��e$��U#��.��OTxq�ƟF'�sZ�ٞq�����
R�Q�ǀ��ϗ�}Dס�e��Ɍ�>ˋ�\�<g.���ч0K�=�O�D�n�Eu���a)W"��y܇�����
�R��q-5kMB�#Jq�&��zv��;P�������I&�-�;��[�g*A�QXo����j�Ǎo�K�<,R�u�8{����Q�;�]c�'�Sp��`�^4�џ-i�����VK��b�eĺ�W���h١��{�X\�ϔ�Ⅻ�57��C��	2����&`��ګ�b<ʿ  �
��U[����U%���Q��L�P~J%��`đ-���9�}P�	��R�����t�	�O/�X�,!i6|ħu�c���G����|Ϭ�0�c]��=����>t��^�L��,^�w}
��%� N������'��w W�TqEbk����lR���2�!��.#��6�`$���Ks���'`�a���� ��� ���Ҧ�.n����+�a�lDg�>MjgS<���<hn��-l��5�˚�f	�yE����	�[՞�v�w6��TE5nRRnx��bOG���(u�R��n`O�*7\S>"�kln���N��T7��7���C���Tu\z���'/BY�x����6[�\��H�x�?÷"��<���K��S�ҵ� t?�`�H;��[:Ipwڭ��Ų��+˨Z�]rǦ�q���D�0�"��+QI#�~˓N�b'�Di��%����-|�#�����C0
�(M��е�ތ_�%�1�5�|�r�q\���+x�msd�o���A�T�D��a��%�k5w(�Ǔտ�JJ��h�J��5�[��c�PtJ�"#���Q_�)��	�{G0�=F�8Nu�u�ݰ�f��zЛlB95$������"�J14��� ;/]mk-uAW�W�J�u׺T��ZҢ�����$���gȡZ�i��r�y�A��]t�.��G��/lm�=1\���0wd�U��;��)���	E�� ��(�����ylN��\6Z�����؈ݺ
���ivl�C��s�6#��?�Ȍ�x�2^l��_$�[̈́t�;��
-#UD�ϡ4�,8�M�����X4
GǑǲ��&$l�|��r���v�2����U\�|�UY�%���^�R4�'����K1��a�DYW�)����?K�gQ KHȃɖ0r��g��'�9����	�Ƴ0NT@vO�A )�!^��kV�0�T���$!�Y�P.ĳ�^������#�eHdS�V۔YL�XN��P��`e �\+���@�"�t"�@!��R9ca�>}�$���%�DZ�؀��
�JP�L�?�i������+���+~�!��Ƽ5"{Kf6�ʲq5�BڴM/v��+nI�	�4D�'�(sc�L^vx3@y�I��2� ��l���(�����P�:m�<�����@�0�0a4(C��	aB:�T^�-�!�BGW�\��Lh;�`��w|o�s�IE������k�IA%v@%�S�/挵h\_|}<����'Q����HkI�Y>�u�����ّ�0���������!=���������l�D�O�Ʒ3>%���I��!.B$�trs�뚉���f�ś�Ƭ/��W�l䯤3���J��V6��<í�K+ěOL8�&��{z]�]�?p�d7�l���RG�O��k�0�-�yLaU�K�׶�J���(+�a@� ���)t�<��
W��m�%��q�P���h9�8EL޽2ެ��O�Tx��R�:�Pe�G�H�H�;2쓕.����m�ć3�;�Y��io��a��������ҽgn�2���)!Uቋ�W�X��[~���p����h��,g)lJ�hnw�o�d�-������/|��f�7t$�@n�Q�)5T�G�Ͳ�v�{4
|hx�T����..ȢXnB�}%����!�k�պ�N�1	��C	���b��U�;-���	�d�D�'�ɗ�5��Ę�^9�� .o��Z���2�-��k�"~�8/��,ΰ��`�〢[ᬎ�G���������O�o�$��L^72�%�G��0�3�yC<_�L��Q��7�J����86���O���[�S�|\Hk�i���g��X~�]�AN�#:c��S0�p6ԡ��E2s�s��Z�ȃx�;�yaH�+bں�k�����t�y�\z�S������ߵa��b/F�Q@2��w�����U�o�[(��b��>x8��M/=.����+�M�G����w�ΐV��_�6)#�W��8�[;�7�3S/���'�2M��;� ��N�XKj�i�(л��Z�-����ܪ��7�yQ��֦�%�TCX!���:��Ql7�_��	oj��s��|��}k7's�`K͜,�aҞN|���q�)w9�I�_eh0&ju�6?�����I�~�;�﯏mt�ω�b�%�JQ��#���f4���b�rg����+�N�I���/���_�H�� �%;���7P���?_�����X�tA.k �Qk��:D��- y�6��Cz4:�B����F��"g-=���}���a������[C�x'C�;(Z����ԅ2u��D�����g3��LS��� ��ܮ�� @/p�����0�v��4��D$���><��?4���F�Ux1
�V�%s�`0��I���$��A��t�?>t��Zz�e�Dء����k{I��;~9�س�^�+�еO2�f֨���z��!�Õ��h�G)xC�L��h�Խ������Y��=D6?V�S!���ӿb�x�V;߃���r>T	&���2 T���6	r�"�	hW]�m!˵����-Ο8��:N�ō:b�Vb�+����U,�k\s��X��4h��K��gא�y6�v�2�u�it�~���»L?'��g���L��&�]�S Y�w�.�q�I�Ɣ�V�U��,m�i�=y�]��F�E7�N��3v�U,�D��;� ��:f[^RۿJZ���DZ��&���U�������{�� �%�_]���&��*�Zh.�(�Yy	���9oG9oV�KYFC�Ҋ�`7��mA�'�7R��vӑ�c��^+S�'P��@ͮz_i�M�c~ɥq��?������Hϲ��d��f;���3Y�x��S�i�f�;�ӱ ��*����:��_�@�nvE�L��̥�iYb8`�ʳ��or�AI9�3Q��-ʰ��A��V��M��A� nE�:O%ҀQ)��5"����� �O�Y�M��xÉS��QpJ�XT7'�$��ܰHO��3*2vs���3�+��1(��¯YP�>����C��$M������QCzB��})��ے���	�I�h���a;=�c�Y�G�Q��q��c �eΊ���3��j��ހ��Sb�o��7&�@���Q��=�_Z&��P�B����9�v �/`^�/�����_؄J����2��.�=�'(���U�d6tS�Qh���x�|���a�#����>��̚�?3}lԶc ҝ*a�<���Ӿd����
M�kP��,TQE�E�o�p���R`|,��O�"��f�Y�wc,݊PP5�3(��}o��������$-t~��ڇ�>R�		�^�ҝ�������[�&,f&�n� lX�?2��Q`�ނ�XrW!=�nK��U"��3��|��LQr[�A��E�AA"�R4�EFj�Q�����ӑָ���+Ə� �$�׌y������	�Ê�]3JwO'L��q0"Жs�g'��GZi�O���$C���t�F�r�w��q&���et��5x����i���F�����q��P_R�D�曄�{?$���7O�$��X/�;D}!F�+��x̡{M���#��RE��9J�)���2@-A.����4�C�����=�g;3|��7�"y$���M7�:���_O���>O�K�)MP���:��u� _,�l���.m�G�[���.x�.N~���M�T\ׅiz����J��^��	��YJ�
�~��8u�ݳ�GuumU��Aٸ�Pv��X2d���C˺��\d������یs�I5F��ٜ;���L�:c����'HĬ���%���$¶3���T&�s�j���aB�(^7Iѣ60I��(�I5��1|</�$����U����]���C��L�w%ށ�|E��
�Ʉ��î��k�YL/�d�C��)��ǐ�6�k��$�5QRC9�ܸ� cڂ�����vy�*ǯ����8�m�~��Ѫ�y��9=��}h~�V�V��M�䗯餈:뎕 ^A= F��w�E�Q�*_<YR�Ю�7p%��*Ă�_C��5Hv'�~q�ۡ=aS������H�r;1;_�-G*U�LL���ߒ]�v��~l�6��@s�Q�;O?���n�Y�	���,Ǵ0I�q�W�Fn�HD�s2�L���唱K(zy=X����G=� p�A����(]2��S������Y_ʝz�#s�� �~0Ð�[d�N(Ԫ0���x�1���1��T`s#q���,�M�C_a�JM�����Z�5/����cN�mH�u#��F�\v��O(v�8�z��9�.��S\�]Y���j&�頝(_�a�GH�
�w�?R�TE�x>0v
�kގ�ޛ�ƃ�k�D�����( ��
�{(���ڂ�<�+d*?�
lNx�\;�.8�e)/$>�_�l����{`�k \*��N�VB�B}�rӳj?���oT٬.���,�+ǌ��Ru���u�ǫ)�vج%�i���I���CiȌ��ȎW����+[�K>+}<��p2���]3�����wrĮ�I��O�������$� ���7J�x�~#)Xa#���CVIh֩~Խ���tf�<++JK�¥�OnL���M�6,ꢅ^`�Ǩ7z�g�-^0�3�	���0ᱥ��R��#�J�!d��v"��#���q>,��V��2����4�۶��/�i�,�0�Ŝa�'�}��ߛ�00�5\&���gލ�W<�~U�2�:�ʛY�x��B��;k?�q/�FE�ę���[T�`�>CB݂I���q�\���L��~�)�p-k/����b�Kgv1 �g�E�
�y����u)��[Uns�@a�60W.+��s�z��\�c�������Dq�%�L�]�%dsz9>1Ϝ���fT���6�Aq͍`G⢄�s1�"��kg���a�1�K_p����3��&�5�_~Wʥ��Ւ����o2�G�2i$��D@k�s���?3W�3�-�.��p��?N�e�����~����5|�\�8d�����,Br�3+'W/�ՈL�EE}�ޒ}Eg�b#,�f��E2ߦD����a��Q0�;y��{4TL�w��� )�d�9�-����[��}�(�����-�k����-�^X�qG��/����'CV��'"d>4�������ǻ؍ch�Q	�n�ƣ
��~�Xq�<�ų�cŨiO�4¯�}�5Q�X��0N}�1�/l8F
Z��̼���RO�C
��)耛�(:Iz6��9�Wߑ��S���)�+g5bBh�fE*�b����U��/TF�|"����F��izi �W��f%Sq�c���8�tDl�cm˪�Ы&ĵm��-=���Uy^61��ǁ�@��Z�V�^O��h��ƥ��	�l^>b�b� ����f�'nfu���sF���*�2�*II�p5��;��?��Ȕ�Z��Kv��n���e+H���F�ݥc�N���l����!�A�>�?�_�|�]S��y�������vaGE��)������qhGdE����-�Ny|�[����
K�p��hW#�Ć5���K�ym񴆵t�Tde����!�՛�.W�Ll����8v=� ��<c㇟
5���D4�ܝ=�߃6�ߜz���J��Yg�QA?����TWɣ+�Û5t|09a�5>���t BD nG����9(�^	C"�X��9���j��fJ�c�I(Z�,?���������W?��;�>i&����hY ���!|�ĈtK��Q]���%A�,m{$�FIڷ$�:Ǒ��CA�]Z�H��s�U� #�X��&�	8Uv�u,��S)�����"����Ǥ*q/��i��Ĭ�V�/�L�;�NV���Q7��ܗ��$Z!
8�m�1���V��{ܦ%}�$����
���`-/ ��c9=�^~�}{��Y��N6LAv��~��y�8��3�a��;y�E��o���4�I^�Gk�+��a��+���	6E ���i5˞��w)C�.�
�\�q��@AxbX"g�'��^�2�f7��}�{!��=���Y�\m�c%�2-�@���r=q�=-¿?]�q��e[/?��;�Ĥ��9B
Zu�}>l{x��c�p4@G�aj�=��IG�m�s��vH�e�� A E��"�D�G���$:��zg�����tD1c�-8� ã1�ѱ|9��cg����}�?H���s/��}|�V]�$ � ��:?�î!Y�:F�.�Ԣƅ�:�]��&2s�f7zM�`��R�V:�B(Nժ�qR�{��$:D�d�M�K��ۦ���yMQ+�f��"bl�gfᣝ;HO�@;R,��@Ps��i�����_|��%y27zƿl>�|Uv����@����Zd����1��.�r��3G
��N�Z�����z�����jK�	sX,�$��>����jQЬe/d.��Y����+ޝU��Bu{� ���8ѼD�﫩>����=�#��>q�(��b�����W����c�N�
��
��B�����F�Y]M�����#5�/���XEO��
���*�H^`X��Z/���$��	���vg�vV�Cz�����
Z���y$�v0�f��]:����[�����r�%�E��������� T�o_�K j�^U	Q [��V��Ne�}0e�:�|h& �9��нfz�r�8��s,�#��I����;bG�W��ܩ�6�`�]�PǧWM�H�aM���+��l��b���qs��8ψq����\þ�A��s���B�&t�Y'q�h<q\$���+�tu/#�(�a���'^�4��^���z�>�� 4��-�� $ܔ�ko��k��u;�@��i�蜏���}��"䕴��Z��d����h ykt��N�T8�"mY����N	�ֆڛ��:pz�!������B!�w}��R?9��O����fI��U����R��^��3�#�šǪ�]Z���,"��BPZ�uA��>Z�D��坢1?l���8[�����Z���fR��G ���-&fڀ4�%:R����������-��6�O(�Z�܊d�&�a1Ѳ��(��L�G���R�Vq��2q��s�܎(�˜%����pW:�}q��z�q���mο�$�P��\Yl?���ؙ�_�?e��z��C}� �.Ƶ��>�^�F5��,t�pr�x����
z�r��,D�
p��Ƹ]ky�d��8�6<@��b��^�Z�7�S��P�����ӷ�) ��&��%�K��b�DG��Z��#@NJ���Zc�`����.��y�9\��'9ɶt�]�������U@兮ΰ"�9'��!*kT��R�0%ն���<=���n���QG�?K�s�f�{�rk�5���2\Ȃ��E�N�Cs/�'%��nk�X1�:�ZZlg6�4L$"f�=�pDÏ���9���ՠg	����A��!�י��`Z�qʕ�iO�{���%�C�WGA�����j���s��Х�R�};���TVB�Q�dk�����P�}R��0*PE@��E1>��p��[�����y �WGm"��,sZ���06-�x���c��_��aJ�uY��i����23��F���Hj�jvZ4��8��{6��s�[�s+5�NؚG�*C?�O�O����m��m�]H+�_�D�R�����k�\�����������]�;�� �ay��'���ˍ[�f+&���%Q��A�'�y)ZLC�̚���'�rU�����\z�V A�dv������n�.�2�>b�B�l��--���GǮ���d�M��l�q�"�	�Y�2z 6�xŉ��5���!:�b�mZ�"B��_��H��6�Ӷ�W��{�O6�C7��1�B�G�{�2���:1�J�4O�G*I���8�$oɡU�z�s� k���m^�YLKQ�	u�:�v��#и]*䎟Ɂd�v�5�l��[��/1b^�q��"z��~E�wd��-�Į�|6\�4�m�_�H�T�4GHDD>�pl2(;�V9qߍ=�鯋��M�;IQ���r��]�̷w/;��_�L��$�G6ZJ�l^���뛛'����!����=.�(Jc��˗���A��[&|"�Y�織ݑ��3
�և2g<(e�Ճ�ZM�ps�5�v˯����o�ڦ=�v`�!i�T������1uw���̍�I	�@p%�pj�^'9���R�bo�����})&%|񇏵ѐT9�e����n�+�;��z-f=_g�%j���9C滆�4�?��
	|���76�D�Z¾��(gyQs����qB"nїx�Ê���o�a�bk#��V\��o�϶�pw�91Is���'m=�.�Q�������RF���ˍ��y�[¿e�-N9Yp8n�7���O�͉��5&�&N��#�Ꮾ��i#� 9N�}5?���Y??/���~E�d��������΍����ބ����g�$����B�[�#�K��,�`r �:�YZos��	L��=,R�^x�Pc�6(��/���"Ajev\O�k5�e��:7H̟j=ō����>����*�z��j�(�z2��ꭰ�B@O�C�>�354��Bщ��k���R����~�oӍ�4V�ȣ�N��d s�Ѕ}�q�{};v�*��g���&���Ƅ��'�a�{�˗�j�5?-���ء��\���01?�;>��U��Oք�'���Qu�Οy��z��go�G��G%0�����WF�R�?�o��Y��{�r���E�2�$��_�w��{	�aY�6;�����V�_r_xd�R����-ub�G�(���Y����s���	Y��Uߧ�I�6���ai��:�^:ㅄ��į�YBP?
-�����Jut����RN��xa��Nb��Wd��o1��`�����s��~��;���S$x0Z����'sEd� ɏ�]���P�:���n�����@�|?cJ�.mc���2j�b]��UA�l�-�[ZS6�G(�$|}��q��Mt�ˊ�V�e�q6�)o5;k��%��2t�k=ߴmU>�e�$DK)a�{R�:��=�ALŮ�g�v�¡-8��:)����҉M�S>�̊ě��J��|�FώVt������B��'�=����9<[]T,PE���&�5����*�]ז �C�1�k����'<А:.����2�J��-����\����C�À̇�Q�2�VK~�����DCK%(�A�֝8׮,�G��5ԔE�}�0�&���V7�!�K���.�b��՛W,�8j>���U|:����2��q��?��2�y����܍�3ϵ|ò��l"����5.�͏"�lsi;<��I�X�O��M��{P�Q?S��ʶ��φ� �W�iJ���ۥ2�feJ��k�s��� A�%��1�5X0?���o�[�s=#��>Ȏ4a�4e�n������k�1�~Ok���u�0���T����D�ž]S��p�z�� a���YY�����������M؝ʓ�Ø�64x���J�j�x��wFHa2���aK��~���
��@�ם-�ȣu�j�9(_�'��U�un�{� 6N�l�Vv�*�&�bQT��	"~�T��l�~���=N��[�vI�̆p|._Dcg��ܮ��TуnYF��1"��s�f5�aj��k�Kt.�@`� CP���j���C1�ګR��v܆2��*s9.-R�(�E'
�q���VT�H�22�x��IYM��F*<`<da=�HQ(���]�Gs5eJ+Ә$}_E��~�l[<��H@aa$���Z��N��t�JU�}�N�?B�J�j��e2�Nص38,���ف&�pI�KD�m�=�`E�w�#Es�v���k{v�#W��ɳ�ʠ]EɁh'4���ɰ�z�G�]إ��V�"L�sa��Ø�]M:ﾂ{�%.�0��RNi n�ҿ;f��9���&	�ᗲ2���nU�G�����{ �p�N^��P��pD���T3��� TzJ��Z�AKWU`S}MM�����J���&�0�Mh3T�H�Z�6���*�b:���x�M#�, �6
ypѨ��H�8�%��	��w,�i5�n��W+?6dC�5�Ģ( e)^'2�2-�ַ)Ȼ��y���J�'�co���]���5S��@�����	lׁ.*V�t�]H;������i��P�w
a5�\ �S����F���P��Y�
��I��b��vl�&�/�ٳ/�{Y�(��ۙ�O�(��u�R6�Z4n\FzѦtaz����m�t_5G�j@jҧҩ�����d�,`GK��[�}�R�R; �Ac@5�����/�7 D#TžH��H�'��A/���Q&��,�m��C��{v�����(�h�{h�q��a��T����ހs#�3�,�ak�$7q���QKZ)a;�L ��� Y�������jK��v|��9�:�3f�=V���#�P%�,���M�G��є7����	�DZKAmugOu�Yvms�|��2�\�Ђ>&*�����qP��l�*��_�����\rd��7�@��d]!��Q�U�D
'/, �`��3�e��FUy�&��aq[��P���!����Y&yk�w�u�
(��_a���a��(S�����ݒ����4������#�h��gkeʬ1�Ƨd�����@��U�L��'��H�2�U�{ih�֕�%�ȁ����CL =�.�O�zC]���⬄0P�W8r՟�VB��:��ʝ�c��n����'���{i4�˄����Ɵk�"�E ��,�v��!E�s�Ȥ:RR�:/jِ^\�B��P��IV���O���B"�QPD����i�S�%�j:�w�a�G+���P<�w �U�B�4l
(j���	$f�,7o6]�"��V��yW����K�#�%������8�P�NI���R�oЈ�k�X��9�������ѿ7�Vm V���D�;��l��O�຀>b&�<�gCd����S�����'�ڍ��+��PF`Cg���	�P0�>�^CP���Hِ�C�9�������H*Ř�S��VU���i�>`ui%NA=�����aKN�����ne�Km�W��LK֎ROJ
&�5-��0�GX��`p�5HQ]�hp�	󙡡d�"�
#�l�BA��"��	�d/��s����H���u�պ�׬n����!�����M �=)!2/��3%^�%�OF�+�0�,���4%�Kv� �b�n9��>l��hL~�=$ީ@��{�^7�յ4e�=O�|����]J/Z��x��&���;��Ť��c\�hv����,ޮF������k���Ψ�%�7�T�#�ȋ��s�6�����o�Ϫ;1�.�n����n`e�1�ߥ[��|�q�4�-Ļ���6Bw�C%����=ϙ�0-�����@[*��O
Y�z�.5���%[��8SC"��c"���O�b}~S��V�w;�ʫ����?�eK|�v����Ҁ1Ŭm�&�[]�OG?B�g�t��+��|Me�����#R�G���1����__�1k?�E��L��'yxφ*E<?�
d���4�;���G�ҋ�qM%���x�P�e�e$GjC�ײ�<�+�sߐP	E�i�<���1�5���_e��78�A���aa�q��;�M1[ee��4�WC<��h�h�qD���qE��(�
ȧ���<��3L�"�\F�o<�i�i�s���C oܗ��,��	�j.���O�����d�h�=����G��J}�����X����h��1$���o�=kϢ�Ёcjm�Q
�{ҿ>�A�6V�o��ԮOTj��u��Q���~c�^#˻>�	�꼠�Dk���oڱ�X� ���2g	yk.l8�6�wi�g� �=d�&�,�1 �ߍR��*r�8B|G��K�
�l�
�L`��J�pɂ�#��Mo���%"R�W���5f������;��U`\Qb�yY����(Δ�$��#
..����nCZO�.���1������8�+���!"���M�p
�b`%�Da���Mۗ���v6�Jojtp?|��j��B.�J� �j�CwS�.�g0tv?d9s�q��\M��ؒx�NWR��ՙ�=e9����%���6�8���0�Q�H�$���pj�������l�a�f��_�Ihô�Y�'Ʃ�:�LW�����[+��<�0�*Wz�	�	��,l&N�Kxd��ƍ�*<��j����e�����+v����	p���>�;�>��,C��g��"�1�Fʎ���x�S� �c����0�ٺ�f.1��11+C{M��Ŏ�3y+=8�0��������
�yҗi��ɷ�7/G���z�_c�P[�$��'2ܽ��j�Gl��{�NB�$w��o�E�%�w�c]�!��� ��3���p���ٮ݉�T��B+ܔ��z(��*2�!��E��<Cw��V��6"I>�#�_� ���\�đ��09��k�G8�̠>7�	��#V�#�:&sl��
�3���Ӝ��CK6!\��LZ���}�2p���(���2F�9yEs�Q_1�K��mv�)�͖ϧx�}��zA�q��5�����d	������`E1*���E�S'4�[8_(�L�?�zP�"R�����p�[�����"E(�\^t�
���X�m���K��xs<<c�Ą��m�NF�2(���UU��l�H`9�]��ښ*��O�B��_�`�������f-)lk�2��UPB!�K��|�b�)�8_���zT��.��Iѭ��p���=�Zp�b�;�2�A�3/\�@��������0�]�����=����f��Z
�!�f�JɎa
f�����܎#�x
L���w�Co"KG�guU�,��}�ؕX��A��c���3�<��ѐ,���5��Hj��ѱ0�����}��h!�W�j2��LӞk:����WI�t:���<nS^5$�*�~�-��}lg]���O0���u�fi�#,;�J���36��5S�#^�{�;��f($�+c�1��LlL�"�.�}�H�ӾW'�;3�B�h/�]6-y~�{��>�VK�y<�!�K�d{AE��u8,���`,�C�s��E��hq��,�U�a4���q�������+�a�X�,ʩ�PLccӮmگ�Q��y�Y�?���������o�iU ��}o��B	t��@I�t����s'����%�J��!Cݏ�f���2���l�����R�%6��Ʌ~1� *�H�'�q��ٰs��ȩ�(�����:2�}�m�(�f�ꪲ��7@���h�B$���HX��w��X[�|2O9ȗ}�یd?y/��������H�����^�brl/ibD)�/������3�9�bB�O$\��)��YA�� �1�!�p%t�'V�"f�<*�^.δ�ꁛ�m��Y$Y��yE��?�w�ή� ������ɿ����yi��S+l���� ���8T��/��D�QbL�5�����x�&|��[q��҇�S�.C��w~T��}E�쬟7�@�D�����zh̕�Y����D�%�]���Q��4��]z�D�ݥe
m	�fi��аφes�g	L�N��#x��L��-���G9hOQ��̳l�;��k��FWr��fU}�ʴ9'f��j�hɈ"�K'"�G)1­��I}�E>��(p�Qw�=s:�g��dV^�\�	˙�=��%����ӕKx��B���Dp;z���̳4�[3Yΰ=N,�Y��,�)WCQ��l葚0�HT�������c�����J�8;����7��t��?�m��Wp_~|�aH�U$��^W���+�V����Vfw@�֓P�2}��M�˽��N���ِkba�~��m����5��v�F[6:�_}�vT����%�>�?���2�#��
�i��!Q�p�{ʷ�.�y�����Vn��H)/�z�ӵm(�Z�rb'a%k���Qբ|$6��b���QTf�r������w��䶴� �rt&1M�j��Sv��ͽth���W��l�:\�mll�����/�auԜ-�D���B˛�Ni��u�N�_��	�v�ݹ|r�@J�V1��z~������gu�AA�EM�R)`��7Jw���)*˚���lP�l��6���E�u�}íH��z��5r���r����m[�Fy`�������l������7dC;����{�W����Ն�M�&����� �D6<�4����a�����_#`�$�����Ȍ ��	Q���)}���zW[6k/Y��!4v,������������D�T��3���U���?a�I����=Z>�s�����~�:HRblr��;(e<d3�|?r�(-{{�+Ȧh������>�ft��s�½��j9�+BwAФ��K 6�G�;@;���U�߄�95P�k�G�/�hN��e݇t2�Xyg�����k^Y�N�G	A����Rq?Gбg�������X"�K99�U�L��vi�C���ê<m��"� W�I���ۆ� ��w���W!z	�UR�j��B�h���%�2�
��Q��?�:�*_	#J'+�YV�_�Ed�Q�xQ����h�"����W"��Xzt��ł�pD�x����cǆ�3��Ke�1I��> *Ëcb���$�r���d%�@|���s�G��������Ӓ�~n�\I/N�����D�~n'�ȳmB]Ő�Uv0�&�l6��2�ܽy����&I�	.�3���&~3��ZO)wJ���>Ϫ�+AW���ہB'<l��%��]�,�触�?�[%�f��mEt�.�aU����Ŝ�U� ����O��0��}�f��H�1�+J]���D$s/*-��/�"r7@���rr��Gɚ,�"1:}1
�)������r���������Y{(��.\���.�:�ܗ�[�����T;�ʰ���ش�X{M�Lβ�A�:U�Ͱ}[&����Dcr��V+ylR�2S�X���(���L���闂r4��� L��������yD��w㦅�I��pA��!�ȼ�	�!���4��R��4�le�z4gh4�L��BGW�^�u�;�"���q��'�!K�X�4��Ja�Y���t�!4���2�U���?��!��DM
폯�����:A����(�I>Ϳv�&+K����z|N�����Wޜ�C5�÷q�.�9f�[ܾs�Y�~
ET��"��WGyh�2=z�E�r䰜�9�d�x����lȉ�!B�<W���:�#'�}��oXo���>d�5qVʳg�`*��)�E��,9���iT_\�i����q�/�axhS���e�cp��P1k�_�#,]�W�`��� ����D��N��o܈��ϒ	�;�s��P�`��-�,1P���%%�E�mk%g}���)Z���#�MVbY=��;�^6��3q$��:U]��X�ع�u����[O�Q�$&����Pe��ق�	B�LW�0'�s)�x���
e}	v�bWЋ[t�K�v���Y�Dr٧tgM8�?Kd��+�b�P^�ax0Bρ�-�@ͥ����ߨ���02#67g�j���'�G��H� �C-�(�u��6O����U�Y�A䊙D�O@ݔy�������ؑ%o��x%p��,*��� b(�$ƙ��i�F� ��	ڪ&�`%˔8*�|C��7�����0/:��p�?�}4����j"{��T	x����S�P�Ш����̾t8^�����	!c.��O��Ծ���U-���_�49tsZ������3��x�%&n��Hf�<����:r��J����^R�x���ևШ�Ky"F-O�$Y}a��� ����E�r�D���E�W7�ғ����;e���
�=�a/� s$��l�5|� *'��W<'����#!��lga��~~$M�'�1�y@�kRyL�B�Z����ۅ�t	��7U���c��7���(\,��p�b��__ .���@n�Z���~�%���o{ϥ��@�3��\aaO���VƦ�"�o���1�B�V��W��@���9_3G�j���{I���%�k��uX,�'�����F����VZ^+��{��i��?�ԩ�ȫ�;�|�+'dZ�р5#�l�d��8�FfR�:�0�m����$at�m��W5�_���7єJ��߂"�<:�D9�Zr��gu���#]�Ӎ�kd�,�� ��ɵr��00�r�4�>Y�+�e^-:ۼh�爰R	�~͇\(a}<�W㴲�.Va��P�[[��IV�¨LA���S<H׼_���Aﲢ�Rz�"{ݖ��%ųX�@z���M(�#a��%�����b�׎s�5^��b����y X)!i`��bФ��u+��}�?��09}����)�T��R1w������i��sw/���]J\R4:�Q�dd����pd$� /Z�U�N�D��$���-.��}ﺢ7�&A��W�G��]]���}xh9�f��:���U�c�7o5d���Sd�jjz�f���<%I�6xsIĬ�9���$�t��[�|퓚Z�C ���(sԵ�m$|�'(Xs�麸&��8 f��WT����+��>�Cb��ڮ��h�I�?�͑�)��=���)��O�m��G�a�j����$�� n��D�H\�LPN�w�'Gٽ<`p��W�����'k���e]��VE{#�Վ��R;�+A���X!���6N[c�״X�"���߰���}t�N���Y+ֹ\Lv�^�?��nn�fA�}?z���5�6 �}�3���zl��[�8�R�Fj@����%i���g��K��a�[ ��rG�#��`>�û~
,�2��gi�m�^���Íe�<��,ڨ�{.h�b*,au��d��Dg�l޲���VJ��9�İ� ����_�?i&��JF@�a��=�D�tp��:M�����9���"d��+h�>}����3�]�~lc��(9F��l�?՗��Z7ʛ�������S�e!|�M�N�zK�V�dۙ�6�.�ŭS�K���5_Dg��C�T�m��3�8�!R������H�g��6���C��2� ,a��Hð���7*w��l�#l��=B��Q� �~���t<h�z'9.o�� �(`i�i��MK~�
t#����"�B㥓�y�����xF�4�
��7$���%�3-ɀ�M*����9;Nr���� �dLP���P_/y�x;�V�V3*�ˇ\RA�-7!��t�=��g�FG~Y��M��Zt�����ي1�`L��bl��9t��Tb*�����������n�B%@Ÿ(�Բ���K�KQ�'�
��<;	\��	��'֘�:)��w�,��#��{7�m���'�4��r������Q�Ң
�c����W��o�Jn¨_cJT���|��?�o~���)����Pu���H�}��LV^%Z�{����#�)`4@�68^�2������-�4?O�g~�[��j��}�;�E��~*�h����!
���6M��B�4|K�M-��8��C�3�k�4ne�Ռ&S��r O��Z��Li��'����HL �B�!�f�^� i�ۢ{���k�J}��,����^�Px�"�R�>�!"����&���?X����ճ�<�<���R��0d����*�s\��dIB,����j���"v�A�x=��I?�o�v�q�t�ȳ�C������n��͡ڶFM!���Iގk�T�E�`x��(�5!3*Yں���4�{�p� ��Zz�+V�j��3�I2���v�S�Uީ�G�%:R��%��_��5��K͊ٳV*��bC0�ۢf��0@�g���[��R�:WS寋_ʮ�������
���N��6����Jp{-0b?�i��� 	LA 	���#b�aة�1����p��.�5&'#}tё�	18�,�4>0�8Jh�G�+������> ��G~1�Y�P��f?~.m����D��k3I�,�
�_W�ƸN��$z3�l�`:�/g|Z��6�4�m������\��:�­`��4�%۟�H�� 
'���)��m��說�\
��b]�v����i�w�^��:ϼ�U�9��2���	�e,՘^��7!�I��0���W٣%|����k�IX��%$i�ʥ��{R57��E
� ��br�ĕT����>���!eJJP3m^;�r�2�]GaA�O��Xk�]�q��`�n�M@��z�눍���Ë�J��UV��C	�[�Ѹs@|�(���,�H���m����B�̓���y�\�(��TMs� ΅+���N�F�q���3�c�v
+��� �Ʒ��,���ZH;k���s��c�n�*c9�ǰº�:n�@<����D�VՐ���X	d�̇b����72q2�i�+p�"M��D�!9���E�]�.E�R1����L���z�\}<�V���I�MGY$DA�h�7ic�@9���[�z�R�_��Y/L�R�թ#�m�y}�T��}�����ZA�����M�F+��Y������&�Sn���=�K������C�X������D�U-u�r�C����� �:y1?�H��{z�m1���Ŀ 3�,~Z�_�^�2�槂^�:�lXs �WeOl�a'��8��r�����*@��r����'b����*#�a�%����ސ�!�iCG�6��k5�g�Ǟ&ij�sĈ+�+`\׹����#�C�Ad}����k$���ϊE��X���#�ښA����U�>	a���Tb�O�|w�}ow��ŵm�?�5&���¯��ϯ�p4Ȥf����Vu��=��t�l�͉��7_����!�o)�u[�LO��=/!|��H���*��sJ �!�5��Y��7���{c
�'�:���@���;��h��f^ݟ��U�+K��3O�tS�W�9fQ��9d����!���S�~���������f�ҏ��@��!8�~Ί�uY�b��?����bAĚؗ�'<K1.%G0�HA-[��M-ܯ=(�Z�ғ��9$�PX%��*��f~�36@��^Or4�6���f��EC����K�t=J���~�����e�DB`Tԋ�a��D�}nR�y�]\�%�O����8�D�yV���"�����藎Ҙ��@C�ժ� ��I���� 2l��� ���s�؞��~m�W�@��h���@M)��LF#�Bv�Y�	��߁��#���⺐k������id
)̸����~�N�'襍H����|�%�9�3*���t�1HU+X�!�����c_{,� ��=�v:��]��%��u�7�=`Jj/h(��B0�K|7K>�GS�9ɑ�S�ڷ�λ�����ʉ�Xʷۧ�Q`s��3+d��۫'�R���O��pv�G�PE-�,ߴ��Kf�%5h���踂�-�/�#E�>���f�=����]vq�}�&:Ȫ[;�q��B�c�[4�(+Ӥ�3��r��U��}��W��MG(�}�������8�Z}O��F�N*l(g��̵d��4�-��j��lw8��٠G�����֤�q�)p�ʳPJsD�E=���^HV��;�	�M~���]y7����f���l�B���������|����wN�FD�NF8y��r�IQ��b���@N�w����L���n�.#ޯԽ���{cm��2�į�HjU`�g�V��>G��6>��I��j1�h�  F�yoN�a�b���-�ז�X
jc;�k��SFe��-��v)�!����2W��&:f4��cy��;C�E��ko�x��S�)� �<������a琛�k=�!~��0�)��d%��<�x+%?[[��Sw�����[�{�Cq�@<x�%tB�ZXV��w3�������`�\�W�2��CB���7����A�v�B��u@/0,��sz���qm5��#��������d8�E�����e�w�ە���&�J�7欳P�wH'()@��T�e���Sn��v	\t���'��0Ma&��4=f��>�|�M80�(�S���Se���Xzx~g9ܼ�6��u��؛|"ic}�
�6�)�/_�Y�3ECYٲ�� (��#2�}qKxp��Օ3��u��۶�#�"��!��A�NU`��H1MY�͝$������ې��o�KӤ'���BY��|����j����a)K+�s/�'>���ET��s(6";��5=�Ø �5
�Jin�`,T�kMÏ��?;0�3�寉*Y���~��w�9�
�7��(���>�}�?Mp������֎I��k��1�3e_b3q�I�U��T�i��/��#��#Ynڲ<)vK	��zd�6���$"���Z�����?�O`nݞ�1�b3�u�X��
V��a��0��f�����e��<	�S��}BM���ZE�☘<�c����5 �BכW񲻧��NP{��8����I��}����e��R���Y�����JF�u\��o��u��)����+|�l�Q��Vr{ϐ/�����B�x�Px�R��iI�q'j�2j��0�[��ك9g�e��à��|�8��ߴZP�s���D�k�DҲ���-Z�3���n�(�C�H
мc���-mDq!/3X+ �Ȫ���GF�v��VY��
z�&����v����3j�`V��/�� D�q�1��Ï��~ ��Yy�l^<nϭ}��D����_��%�F��`٩���aI^�r��Ж	��X�����3M��)N��9d$o������7�c?[�#���7	$���\�#p�`�/rq��V�wϲ�I6��[�?]��ո0�|����a!3��ι��>P�W�Z.Ц&�4��Ft`% vvĆ�50�������V*���8Ӄ_���6�ҿy� ��Faۑ�)Md�ς����+��}���ƌAIL�-e�N�U�̌ʪ���>�n,v狑������#Fj�<W�0)�hq��"�����
���r�xģ�T�	nɢ��ޓ߹�[����Ƈ	J	Ź�F> �﨑[���儹>ה&s/��ћB�L]�?������Q��@���Y�j��V�e;6(lޠ��N�L�/�������P8��ʧ@Z�oI���EC{(?:�Ǚʗ{��Bu]QHp\t�� :ھd�	ep��i�yd�����F�s(sT�^����C����E���N����#d������m���ճ�lvN�;7���߰�*�^J*޶Ύ�ܳ�ɂ�e>�
�q�t�It��9��+o��E3SF�]x�5S���.{:��JC��E��_�@��z~���%j�V��g)�����C��	��(��7ln1q�|�8{a8���Ւ��rS�;OtM_
��5�N�<(�&��nDҎ��jⶴ�ܙ3�ڲ�焒��vn����ъ��"���3��*;��H�F ��l?�ѼP̟(��w2Iژ���%�]�������}�	�J�I�L/w�tM���Z?�$
���=��)=�%0��5.'R@���C�����p�J�$�1�_}�* �`���e�!v�� �������Y���Q4>�Ya0v��C �Ր/%-�����&.7�tF-pE���زp��'u�Y�6�߬T�&�KgT����
���^o
�oůCf��Sʨ��-�@zw0�*��u�9�egʲi2-҉��b��gOu"�}�������;|��>@��Ӟ1��h�	�I�_�<�x��:�c +	B�s�+� �[�:�-4�*R�"1ގ/o~�ĕ���u���\��V�v�$�=��g���n�Hy�F`Ye����gw����u��g�ɭ��Hy��b���z�,�Q�{P�$��š���F�$ς~j�$����~�y ��~�@�`�R���>�)U�4c`�`(��-���*�K�~��D�l�E��P���	J��	�W�|(����࿎�El�\r�/�|%��ߙ���3�1�m�����C��z�g�؟\�����a��;���b���ЖXD]쐻=�w$����2��cR�D����40'i�{\B¡8l*s$h�������$��(�p�?��6F�o�Ih0?�����"A���P����b����m�W�C��l��253-bqd�m"�b�$�X���,��ڤ׼��O��h����3���%�a�Exi]�*�֠���G�I:6����-�w�����#7���w��u~��K*�x�}�
����q$FFf����FVfJ%8V�@����9�0�l�|���
jz�V�DĜ[��+bl_$0�c�%��� �,�|9d.[���l��7�ơ��y2Nl$�����]�<�ҁ���"/���,�+7	�.*��Cc�Yx�?�9m��}�6ǐ*�\��}cĎ�A�[�Y��~��K�Ý��:/�f|/1�"�U;�,y#�̓*�)Y
 �hm!7���(C�5�(+�O�����P.�X��g%B��+U~懪�����ܲfD$ ���_W�M��N�7uG����8+���_a�g^�����tE5�s�=5�����p� 9_���)��ps���>I�jn��Uχ���B�f�߬�����;�*T��c�3�R�r1�A�@&l�+A�N-��Ki�Nc��S�7�G��=��{�������D'��n��V�R��(=��m�dՏ) K�&�H9lz�(2��m({3���%pP����Xo~d\�Ѿ���i�L�RE0ُ��8#B��s Ng
3[�mkwwqdn�1������,�����l��1<�.g;�}��mrr�.5v���|X�b���yn-Ӷ��,��3_��_��p��s|ޗ��WT��(��N���s�
��r�s<��C�k< �8���h�lE���`r6�xן? |�^'�����#S�T�@��ZE����"�!!2<M��i<!�[:������0e�XkLg�j��K~	��i�,���7($m�{A�%3�f�x���6���'o���7����U>��Q'k���xx��F�0�20��}f�3��T �W/��'7�It����w�x�N���I�l�]O��'�,	`��Q�Ap{ڎ	٤V��*��xʱ�4t��R���.�^`>���P��32OlN�Y�h�\נ�����b���)t�z��Z5��A�,qiIʵ}1��h{	$u����3�vS�{����a�M:o���J�� Df��0��㶅�[(!���}@����)#+9��g@���,�,�9��G{1�۹�.����:�ɤs��xh`d�"(�,�����+FD��4��b`�1�r|�)ӓ���dV5X���3�a�`d�� FG7ׁ�:�jw�J�8�/B������L�� �#h\i(ѧ�)�&����`�CGNp���\j^�O��߀WG`:ڝ|�6��p�8?=h��4�����q��c�
}o�T��J�jT�!��(缸��stCT�=x͠���D��,���up7^�?|:��g�6e1N�t�G��٦~��6�2��P�5��M�#�:�m39q�~����s���gFV�����U��%C߭���оm��T#���Gw�=ӻ����^���Վ��q���1?F�.�Ƨ�_m�u�%V�1gW�����f�p,������l�]�鱗nd`���
x��di��iK{P��!�ӽ��}���������H�׵�o"�L͑L9FV���+Eq�{����}��p,x�yc�W@"�%���qJo�����(	�+h#��yS:�b�֙���p�r��.pdS�J�B���	�\��Y���YhE����`V���AJ���&%I=l�������
�;�^56��e����}r��gM\���(�T~e,#2�n�4'!�S�I�R�����n/`��_p'�{��ܷ�C�?X#�E���[��V���^�+e��\M��)��9���Ң�>&���$c�(�Y�	lF�Q5!���(i�&������9�
�����dnd�s����tE�FΒTޙ�!���~S��?���M�0�3p	!��RޓUX�{���&uxx�S����z:�x!�^���-�rżY#)�O.����{Z�a]����7r�5�B�z�,����*j�-@'�[�� ��e�S9,(8!�/e8���؃γ�#YE)�?6���~"B���/,uC���}[N	�up
���%���|�e�d�p�c`8�3."_����K�L؛��j>��l/?��9�����jROQ�b~����,�2��U�ډ ���v��4�4kd6�Iti7}�a)_e,�im�]�a�	.�dFϴO�ڟ��z��.Z��c�.g�����
T��/��H��/� �uÁ��X���ڂ�]Z�?p�����o?��5��Lr���4����\l(<�r�~1%�.�\�W戕�����G�>��.+9Nc,K���D7l p�)��M��ɮ}2h3��5��QLՔm��;��p��v�E�7Al��'�eY����]��_�A�
�$�؄��gg�m1!�RY*F>C�Ϥmٕ���P��ܠ�
�>1��/'���F�,'5�n�(C ��Ұ�+��/��׳M��/��	k�{�k7�����_ġ���R����(z��|CY��	{����(������<܅J B�Xd&d�q;:#1�.φ��Ͽ�A����张Qj�d$�W$�~�ґ�w�n���s�:�,�.�2s�H$0��M�Y�G�_����F��p�k���x�/o[pw���\'}qup߲t�!
>U��S��~�	���~�t��y�/���-�a-䖊�آ����Z�3A\-tW*�#X�ÍM�=����q���=��w�T~�ra�H�r��������"�V��%�P�F���Xzc���G��fKɛ�.53��H�_fX;� �f�Q�|�N{ ���mt�v���^����ūKvzuߞf������r�
I��ƪwb�G���&���� a�N����)�.h��nO�~�Y�n���z3�y^y��7�~V��1��W�C�$/�1�I�دr}qyS��ϲS?��CŞ�r#����Ѝ��l������A ]~%��! [�;��uUj����Q��׀�����M�/�r$�ŉ4=h�������9�{�r[�o�b�I�gy(0Xy�)t4�:e6�Ei�_˱T�Pk�`I�AZ$�e�P���|�-����æ) �z��]}���v!�	��V���=�}*"�`�<�0�����=ԯ���OD.�d3�� ����*Xph Υ�5�YW|-70D�`��'�!�G1�Ӧdea�,���H/N�XA�����':�繖~2�.�G�I³���P9%vT�hsm&+ (�A1<�B��a}@���I}�$p�4��&k��2-�,��:E�h�ٶC�g�x�T���w
���F]Q���3<�նN]i	��|��h��	�o����:E���榃���q�J��{�P�,�q,�nz���5Xt`Q���2
�gB��������|R@cSC�x%�ag2�����t�U<�!�eߣ�6��ch.f�}���MK �U���X��%}��}�����_���)ɴ��
��� <�b�3�C�x��N%r����>��,Ǽ�X�� <�O����!{ ��R=�-n��'9\���:]Jy.��<�~���0�q'�4�qz?
��֍�j��$�B-r��<�Ci�����M�䊡�E�S̨#��6�CVuQ���DUҥD\���Ng��:�ok<�݌}�?S"�72�Əa�(��4O�Miטv|������b�Qq��L�xkv��.����y�bד����3.�?�*�����,�}t=�DO�E��'qY���(�WI�)��~Q�ymO��g�^5��3.{�$?�%��J���i,�p@&����_2��AiH�ap� j�?1k]�4�(]Csgd�?�&1����ЫH��"-�����0���{�5v���u�(�
D��M�B!CiCj���0c8k��:�J��%L��|)>
������f6��X��1Nb@��&�k�Ԛih�~�ⓕ1�� H2���C}�şj���l�a�E�� ;$I��됢�6l%��d@�mbD%��B�<3g��;;�WP�փ��s(~(���f!���T��T����#�����T�p�����HP��S��-��ţ�l/�/aESsz;���o<CJm�_�|�]�1(�������"#��׸������C�٤I�t��YZ̠G�"l����Z��bA�n��@Ȳv'���"(w�%&�rp����`d��8�|���5�qw!6	�o򬖔ξ�_�dݿ�IR{
4�Jg9�`�A�Ts���V4G�NUg����:��x�)_靁.�E-dj����TUYѸF=k3�[���ڀ����K�.g���@y���;��E���M�s �ǥ=`n���1��)x9�X��ե	������3���#+���epҵ���b�>V�5���p�����Uٙ�	����"��DV�A�������0Q��¥����i����4�s��[�LaY�?1Ǯ���f�c,���J0=�e{gy"�,lRP��oG�@LEsɡ���c�ׄy��0�O�>B��$qK{�]Gd�"A�̗����7R��,��ZpAp��ĥghw@��mr����\���yI�O��i)ۮ��O�����(jQv�v�8Kܑv�Ϸaq�~�(�Ņ����	d�d|D��y��5�Ce ��X�>8߀��l���\�G�k�l��o���<��������o1����i�j��<��p(LS'#��Z��7 *�����7�<<�֍S���5ϴ)��Oޤ��_��p��_3���e�=����K���􆆭<�%s�ǀ<g��H��.�O��e�G�jC+?��+M}NGb
ǭ@�L�p���%+Y�sto�0�)�许� �4`�T��#XH���v�ރL��c�``�ޘ��Qƭ���9S2���G� �*z�+[a��Ȩ������o�Z���+��V\�N3�����6Vp�֙��U	��尀9�U7�-a���W��7f��zR/^"�rWU�͂M���ԯ�d�Z�Z��[��N�@}�4�J&��9{G�D�+>�-�����O9b�/�X5G>�~��k�L�U���7�q�&���E���b��_d�Td���%�cp6����&q�;[(�f(��M�&� �g�8)dBK��h6�pq'��-od���g�S%��!:������������U��ќ���`��I���Tڥ��y����r�-&mf��՘T����Ъ�	�c��C�ٶrӭ��kh���o����`S�L`������E��x��[�b�i�\=�� �\&��BX�	���%���l�c�Lޒ�L�㔸��GQIN��B��yC� 6�����l��F�Х���'IVM�E� �j�Ӓ��z\��u�u �=�x%hn�Uj�NHMx�|�i�rIМ���(��ic=�`!�?�իq<�mB^\ten$#9���fa����|_	JH�(���"��Y5	ϱ��W��;H7|���iX��m<SQ�R�HL�����c0���S�[�/a��k��ذ���������زK�.^�.�3c���73Č�(�M ��Bn0 Ή��T��,���\��X��\BM=\
��m��0��C�NA2:Y�F���������a{����()��7pɣҸ![�t�]d����R�zb�l{e����P0bvi����RB#��²Ո��A6F'וAr?�ɒ�\j�2.�/��{�H��PG�3�ƍ
7޹G�jJ���CI��^5��ռc�"C��p��2�譛�U���K��,wT=��d�/��"(\g$�Ճ3������ �iެ��:,N���f�~����:鸧sR� �vK1�3�0���$�C�Z-�ߩ�w'Z9G���yiR�M[���j���|�����#��DR���y���E�I�ƚ�D�0�&�k�4�������bH(����i��i������b0�Ot�T�k�l�Q�٤ �#��\��
1Ӂ�#$G�t(V-��Y���`�ہ�X�DP���K
V�ˋ��&��a?��;o�b�z���d���w��dV�@)�8���T���Ƨ�%�M픔���.����b(�<N��p9TgR˿�5�Y�cez���,qB��kě�����,F�Y!}'�[Y�� I�����v� �c�%a�йi�GW�2��ڦɰ�'��͘�F�%�r�c��|!sr�Z)/(}��(�J��Q/�ǎ@�Q�>:J}UcK�[�
^�i�}ؒ��	�,��	�0uM�3�rbK��mܢJdPs�̯Pd{�)D\r]	�L���ޯ����;�	�%�g�g�`�OBEuEk���9]T�cdX�G��C�� �+��6{=$�����Ŝl���Y}�5\��u�"�W_ooW��uJ���Г���/�+�X+&⓫� ��?vft�B�=-p��ɺ��"��3��P
���u4���u�Z���&�xl�����x�٭ �s/"A��#>�r�xلՀB�^hr>!�Čp��j�Y�Af�8,.��;��>D�`�~'��Z7�^�Z��h�����m�����c�H��5X�@�7��F
ʨ�qj�*�#�;��RcȠ�s�� j םV�ו��C�̋S�Ya<���Վ�n��#i�R�dƞ�F.hu)�Rl��?i�X��ռ~��1�:�;��t� #׽����,�p%���v/��g"Q\�i�I����Z�����ǁ�Oqi�pv_ |fʩ���.��#j����1����!IZ#��1|�Պx�h�(�L:	;�R�"3�W��S�쵴jm��sa.?nW�����1�@7\:����>���~kO/�-��Lb*GD��Ťt!SzM��|�Lj�m��h�}��P,ʤ�oD��������"�Q�1X�wp`}i �&��$4$�Q��:Jۧ�]~P���=��3�X��H������`٬�z�}�ٸ�Q����C���%�~w�*�͡�Tb��~�J�S�	v����h����+X��x�Z�K*��_Y�$�9��-��!�,�Zbl��m�T��z(�����ژP��j��6�+�(�]^?b��Z0Z����A-���,���p�����U�2��A�Vog������U�~�2z@��&���4p�Ȝ�I���c��f�؅^����C�i����>�l>�ڮ�z�~V�(-����I�6��$���O6{������Xc|(�KXN�z`�Q��<�Md�|�Tm�52�+H+�W���p��������R��A���U����Y{��,!ă���}ž�
3l� ��D�e�2o�Y�R�>�+P�2�F��~N�,���]ExR�'�V�ǁ{XQ�38��w�3�H1�ԩ�l"�0W�bф�y�����.ņnU�\ǔ�@ЇG����E��7�f�+�q��`FSt¼�������cK"�Q7��X��.?m��(~:o�G2�"��?�vs��M�M~f;^�	��s������A��qRh*N�&*R��}���zA��6��\�ڧ���AӘ�`؉]A�3
	og�Կ[}�w�mZ;�pz�]�cdc�)�<��|��ْ_GC�{�N���xEP$���3 �l{&�%P?Х���p� X�� �o��B���,<B�j�>�Y���h&<*g'k�
T�g���-qtޕ0����y���:�L�-�A�AѤ�=��tx5߰���UT&w�Ũj�i�K�X��4�0xs1L�H�g���/Mmv�G$i��������v"��?�阨9��۸�۪X(BF1m@�v*o!S|=
U���5܏q+rGP`_DA�0Gl8�$y���u�c��
}-P�t�TP���m������d�u�"-���ْ�2,Y�� ]��2�m٠�/���ƿ�΄����?��@K
�\����&�[u��ˁ����f/u7�c�������D-�~C�z�D	֤��1˴h�$K�6d�go�N0��b;�l<f\�[Iʳ!��_鸰�[�2؍��ˁ��ءO�'k�7�Έ��í�$�]e*���%���:Y4�܇5-�:�:���kQ�R��o���h�|ʞ^t'�	�zgZ{�&Q����S��(\Ӱ	\��nXhE�_�8�<zby�Z���?�w��S]���&�͜��׵���??"�9���2��$�F��dc�tj�1z�ʧ�c
9��0�Bz��1,�gA�ŹvAb3C�ᫎ�Q���☭
֥��d��ڭ��|$_<�&6���1��$����t+��;H1�����/�5I��3y>�����L��D'������T�%6��B�n�J���O^2���٥'���/v�^C6P�?���Ԣ�q�ᗦ����Z�>���tl#�Is���d��>~���ث�r�Zr+��ﵽry�\B�Bq�����3q _Ol�xZ��^�8?;�S��-�����u������Hy�d�?`� �PkM긴K�]D���u!\K+P�Ͷ���)�*�/�l([w��T�@�횤�]�����&ԩUZA�8S��6��z�塃�zxa��v����__�5.��	�d6������B��Lj�t���:��k�;�O�B�:	ڃ�=ԕ�G�'�l5m�O�����k��]؝N52�&+�Ee�X��fz�{�G�<����4Y0��#���}NU
u�8���[����֚��С8	�Vߚ�CQ=�5e�ǀ�	�1���2,��iX���ͺuX�jQ� ᦂ���n���|e�Bٞ�t̃��Gj3����5Gf�ݝ_3�8��Wn�D�O�w�հ�w��1o�u���DS;D3���d�1X�όY��W����:�v�M�F�/	#B �l9ik�-�ZG���3���C���M��AG�x� ��0U��ɭK�������Eg\���s�(�4�
��g_T3�2��b	z��#����qV1m��f�㳆�?y�GTn��v����N��& ��b����	���7/��Ӓ3�)�����36�a`���F'/�ͬV\����J,5�7�#��l�ָ���R/�t!������\]�m<"��w����\�l��sv�E�K�r����>�zi�-�m���f�.�$�N�[�k���5�_n����=1�?�6�BXT¨O�v�-H�h�|����Z�ܘ�<~[���V�/�7�}u&�c?s�/Rv�k�K�/_�`�i�A�\��P,�����@ݱprux.I��=iF��r�FTQ~L���Q�p&c2ʈ�|�+Ϳv�:80스@y�{�cH��L�����k�����E|��ƯO�K��2�g���Ra6�|�9�Q� �կ�n#B���j�vY�)�������Y0~��͌T�9�=Zб �ѷ�;�3`{�2xJjA3e��孝����a��JC��a�v�+�ڢ�����߷�����u3;�8QS�Q�`�D�sWI��HXj�8�X����{��~m;�W8AO��9Y�F����[7��~~��K��`�4������]1}6�^���W��dY,�Fd|�g=6��1���F�PZ� !��׎�6$@K�\{"��5����bz�?c�ډj��uN��5rJ�f�uv?�Չ��w��MR&	���ƙ�t�0C	����w�lT{�
�e~/n%�/��mU�O���5lW�ק`&�N�ʆV�w��#�:{�n�5�}0|)y;�>S7��~
DlzM���(&:��ȩ���3��L���5O\�Y���(�Z��w䁛��4��~�~���gD�4b9�L��Ǯq��\gn��39�uĒ��<����'R�)�Z��\d��6�J�@dl������P��X"�U�| ���TQkk����HYJ4ă_0��"5N��-#`���������
*�Ř�}G��rF��Гf8�����չ�<y��e�",$�>b���d����B)�7�4&]���&Fї�)z��5u���a�B��s��0��	��x�/n�e�RPﶕE,�gU��(랎���{r9�M6�	7�l���q֣��uL���eP1��?AŴ�'�
s�N �Kژ\-��5���'V*�T��޶��9��4`g�JB��n��E�"[(5-É��?8(8��)H�3�f�fT�9�Y����RL9l?6����s-��g�I����Fv}�^ѹc��1==~�\�Q��> qKG���+��� 	M������I�v\o�ca_���/M�ΦA�S�9qM(��09��|U6�� �O#�B�)]6��85>��p!�iLEy���e��siJ�~5r����*f�(�����#ɀ����_�)8�\ɺ7�ʻU�ޭ��}��| ��l�H�@�o���#W���Y�%��Fh�}� ��ڙ���$ȡ��3��������KQ�;����X�)Bb�f>i�ʁ�����p�Z/�33����'�E�2"�q�ԉV�i܂0���Q�Q^ֺU`�A9w�3��#NXS�0�z�Űa��X�4'P�����C��@��b@r��tS�����4�ۚ�a���G�BaI¸"��?�����:�!��9�;�8�(���}����nr�&�����(g����,����AOPτ<�ӕr���ɾ,���|��ܳ0���)�ޡ� \K �0
6��l�7�V���V�����E��$���Х���Ԉ��>�2��F�@qRufK��¾ѻ���1_G �|��=<��i�N�D"�/��1����7�fS};�D��+��l��Ȩ��%�Y��7�sT��"1K���f�1 ��h�|_z�s��J�a�؋v�9�u��7fW��:)�����?�|?c���;~�a/��	S+�$azf(qA�8�ɻ��#�>����y[I$y�h���,f�����-��0�Q�� I�QbQ\��']�������s*?;g]�Jh���ȶ�Kg\��kԌM�"�4��ˑTp�^���9��G��N#DP�~V�K� k��gǑa��fY��&J�,?��FnN�*�f\
v;���|?�[[��錵�V��~��36�s?�2a��O��0�'�Pz���!�R��4(Y�~��܈K�@��U�潧ߵ+�@*/LxRV ?Z֬mzœ~sa��k�X�����%�r��
����q�A���̃61h�[�>�>��Fe�Th�ݥ��G��c5@\�O�]z5�,d����j��TZ�IP.�V�_9���ZL=pITO�V{�b��
�zG����G����rhn�ǳW���3�kv�XI4�P��0u:�6޵oZ��n�]��F�HM�����|Vexu���F�u������ד��Q����b�~s77�2��4�[Q'����@���m/��<+
�;n��ӑB��r3�X9���i�.��K
ų�J��/!]:��ݴ�rY�|z�M�@�M��[��0�/
C4�l���_'R,�ɢ��9��bD[T��*���a�bF�V�G|��kr�`x)�� �Q~�"Q��2�b�֧-o����q�d��A=u��mV�QS�t*\�?Zl��L0y�(��*�c��<�2d���]�a��|?m)J�cK%�Fh�.D�p����f�`$,�$�QP��q�=�p)���_:�Òץ|�f��f�\2w��f[7��2���A�P��<t���B�⡮s�d�DK��̟{�H�����Y㈏��������܊��>%�5/#�����.13R��S�� �M6z IZq��F�F%>���g j*���k��C�p_�7uWK��Y(G���R�#Rn^~�V��Y�Ei�����SGƊ��ߢ��a8�H����x��(ӂ�B�\uu�DmE���we�^4�ĥ!+k\;�n������HZ#V�g����Ӆ���k�`9���T�X��5|yb�!����+������^��E�:�a�L�gZ< 3�7���Ž�e�zNG�$Ϝ\O������2:�?�@�5���tO���R�Mõ�f
6���\d�2�܌�Y7�X�l��]�L��G�e}�O�DNW~O��^�Q��19,�}J��x�UfXyө��ͻk�F�3{�L��R�ŀ���|n��v<)K�p�Ƈ�z2�MW
�r||�(V\�2�j���H��i�J�,���j���1�I�>���i/��|f��3�L���HѤ�Cu�p�_�+�L݊�P]��j� ����P��5�E�:�?�b.ъ����ݼ/J�S����0
������-N�%+&��n��v�_Ju�̬�Y{8�3�#��v<c�)����ɕ�d��>&��Kr>� ���<w�^�fnM�4�@�j	u�j��1�q&K���^�����R�CË(�=���d)�La,�~;�^ڨ��͸&.�sx�!��G>5��X;�&D�ѫ��~�J�&f9H���c�3�ZC�OTT���$ jկ�_��J=�=׶�Q0tD�N�xEM)�>|Kg��f�lS�\��C�@th�j�߽E�STe�	���~˺3q3l�p�iGw$������~�p�������	!&.k���LD�_OtjK-	�m��꽌Y�ZY	� =EE=�s�k�볁k�8�?n!6�����&�ڈ��c�7׍����Hi����*7�������}��o�r,���F]UDk�pV|I�o>��[�7�0_���A�>��g^��rw���]��ߋ~�W��"�D�r`sw{�i�2@)�w��4L�
y
Y�����E���5-�?%�/-j)j��>����f�	�2a�p�^ >�;5He�w<;���}<o3�xR�C9���uJ�,︂�e������CN$�xg��B+�ۀ�o�2h��h� {ޙ?�g�����P=n��a������̔�϶g��U�x;��.�X�kUݲi�2j�q)���d`�NM,���>��{7^@e�x����ԏY����f"@��d4eƭsW��m���PC���j}�����v�;`����y���&ŒA�ݞ�h�	�f|��i���Ť�=�g��c����q 1v�w4L��@�ϓ��fA���DP�ejO�G�~�h���<��B� �? ��Y���0�l#� jL���l�M>)�p�ҥye�^��W��@G;�C5�������e�xjLY��{gf�[�'�&A���fU��ll�ݯc����W����	��U\mQY���/��w5D悓�O�D�˟�����<K
�ho'Љ�ʓ^�Ǽ��`	�T��V�g�<<��G�k-v�߈��s��6���j��Q]W�\�]�f}]�2(|!l1����)<��&ڝyA���B~ݥ��}g�F~@sXZ1�)t������J20$Ƌ�	Jr?�w�2����L�������Yf���P!#0~��jV�#��ɏ��⨙>DM��f�IZ�����j�����tf&)��r����]m��_�:��nד^�W�)��P
�d*����7�G�9���zΣ��E����40(Q$Q�CKj.`���p*i�M��(���ukU�+z����r>�ŭ�'�?�5 2���t��k�3S�"6'թ�m��q��1�	_��%C}��4���m�E�K?0�X�`�R��ѿ�AeF#c[�K�U���o'�k!)��Yw�K;����S�t���PP���/ /����&ϔM�є�?����E�>�V�.4�����e��o�(��f&a��^��V�صL�P}ߠ:���$i�N���}	�z�Fum�"񹕅@6S����ǘ�d��y�[C�V}��s�k��;0[�����ʣu���]��֡���uu��o�Z�OY���=�����>Ip笫����6��ũ(�������p�675���t ��@p!v��@��@yo2*j��&�4�@OE���녈8���<�� �xu��I��ŧ�4�;�+(�h�*̖�m7K�cO� 
��ǨZ<2��b�Z���H+pU���]W5��c�Q �T_��W�cf���w�C����k�fBϫ�RM8ЙT}=h��џH���[PQ�900�=�$��W('��o��sn�%���>k��=W"�����?��dT4�~��ٱgR�y�:Z��Q����cЬ��T���]Ȫ�fp�G�_�e�%?�b5B20M�Òv���(!�:�0>c��I�����&=�pƜ��׎�3�9s��=3��S�>NW�l�Vc���hӶ[K���򇮭�����uLa�7���e��M�.sQ�H:˗&T���T������n�x��-%Mk&�p����k�������k�?�!M^�,��
��QY�2X�x�&O�������-�NV�bU~���#���\��������p�����D�ݬ�-�TEͳУIݧ���(vY=?!h'�}9���IwW�x���`9�=�q��M�o{��}�K�}8�=oV�&ϲ+�5ypF%��E����?����g�5�-��HA�5��)������	��^�M���(�q	}�o�R��l�"����6�S�Z,���!�
v�*M���h`0y;��%���[��^��&c�Y� �4V��XI��S\����8�q��+qg>UH ��e�E47��e)��������73^::���b���A��"�V��M�$��U�7��C��'���=��l�����L��]5�M����r��P�M`����Ot�㮨����Uh^Y�����bQ%��[�V0M�JDK��1�����>.����H��d��QU[��#)k�v�˦�h
ekFb�����)9%�D-�Vխ������ȓ#$�?5����X\G��p�I�kc�R�R#�p��سó�C�[�GlW�P+��0����Yс)������j#������#Bxrྖ�j|V��A��W�����O�:��[��u 3�\Ѽv�_^w9G��d�t�t�uh��$��e~��U���YDl`��5v�J��+o��9�È?[��-��cs�4�^Ɨ!��'6��܌*�7���ȡ/2��vl��M�)�<%�!mu�m^@�8��tQ�Ov��f l�/�"m�����FW��Z����'�N<���;pG�k�]�j;R�o;�V�N �tR�|�pu����6x��1xXr�#��"4��2�����E�>& �
8�3v~�k�_7;�C���?�8�S0-��V:wHp�CѪ�0�U�,O[�~T���������dJ�E/ ��:����͋L.�N�~Բ; ��=�D��]���m������q	�
c�q���齧X�in�mf���ݻ��g����W�+�K�  O��
{L	����x�夙� �a<ҧ�� ]�k��R@�y���Kw�k�i��~��x��G�YZ��$S���}���sr�����,#���)ՊG�L��ټ,������!iC���
H��%GFs�
�	 ��_`wL�r�N�4����w$��>E���i�$.�_�%�\{��f⮝�~K�"�Y��v~�(�'�z�v����\L��6���F�W�� Y���'0�(K�m�κ%��;G��jE<ܤ�}�S	���f���R��}d�E�d��#_�,�b�2����PF��uZ]�H�?�RV4l�%e9�>�y�,3pMml��߃l�j���� �u.8���A����w�6'�P5^=fu�C����
����ޗS��o�7ow�y�ܕ/7�a�5E'�����l�Mc�2�x��;��?�o������?4�h�����Ǹ�����.�����I�zfe�)�=On��`��×��¦y�ܣ�1�Z��k�WL�K�~6���X:��iP�A�k�4���3�v$d�4�G�LV=�s�!vi�Dy�,�Ʊ����^����Mm+���P 6��`N��������l�Σr�Rb<H-Ҝ�J�0@�jm����	���W�sQ#���;&!�hDSf]WY8NQ�D�Vm�<*��U��e�4)�3�s=��P�ݐ��5'�Ĭ���J|�O%@�2�=PXK+��K�����j������4Q�7$ț��T�g�7(ys-h>���J���~�Z<� �X�c�'���� ����������2���ܨ��7T�ҧY�ͥ+>}�T�}��-��6$X�"��5��3�@�ۀ߶̄�����Ӑ���&�6��:���3@��6����(��]jB�&u�?<�K��/?�bX�%m���|c�8$�Q� zg�	?��}��+cbcjK^���b����T��CE�=��M,v��7�Y�{�ғ���+^����}���*3���_U�T��:V�oڕ�c�׍�vŘ-r%��\�6�z���:pVl#�f_ؽ
g����=�
CU�ԱRjf�u�t^ȧ�.9x��Uvn�c�?xąPs��m'�T������Z,j���/��:�`7+�ؙ\��e]ba;.�Myz3�VX�N�/���J��Pv��*����_}�ôh��X5d��B�k��@���1��NN�2��+���A��h8����~;_�B'`[�`��U~�ۚ:��N���W�;+��hv� Jg��G��f-|� c��q��n5ě�Ձ_��X�	2'u<��PC����)�h�.���D��a��@���C@[E]Q���f_�������4WC������yB����癋�uzV��  Z��y��a�zA��������ߋj�<'7��B�~e=YoTSw�kG��)�����i>�kwZey�m��`�EB(�\QO ��o%�}d��w�\�leE�3�P�vD��������j�gK����BbE�ZQ�/���V~�ޟ�ىs�wg�lI�J.��N��#��3�I�{�,b�d�Dm.�CuYdS!i�M�q��D3�
A]�:���F��g5�����G\F71E<?�#�&��5��1��ᒛB�Sd��]'���nw����yg��F���-��Q���+sH�|NZpB8S��&#�Z��~��f�N�N��p�RoK�~�$Z�.�L�/��M|!S�V#0����pm�l�~��F��{�Nd��,��b���t�O�+�x�Ky��Z���7ʂA�j
���_$�],�J����6�+-[mu�w�lrB�j<F �A$�)+g9a�Y�*�YA�߲�
������<��r�
d>ȧ
H�.��׽#�[N8�Gq|9��f�!��G��i5���2!��-��E��nCm��R�%��F8��B�':���l��έL���M��Zj��� �=��^��hZl~��S��A� =��<y�G� ni���b�$�h�4�ǳWyTH�.Fi�
���~�B9Z7����1e�� <�ݠ��g-��M,.!Ws���mv[��X@�Y>��ou�R0�}�E>������y�����x��f��8P���GT�(��f#�X:��IJ�Zy���NP�#oȂ�����Z��A��?甙�"D�۶�9������q��TO�����Ąs��u������H/�VK���9�`������C����3+)A�Q}�3�2e��p"Ew�?uci�1nCP�@IC�v�{�\_��H3�X���'��v.�'�r;Q& ���)���F��m,�ǲ�q���
|`�����:�<ۧJ��)g[���&.H~ jM��p�7��y�7B�2`�it�I��xٿ�N=$=��j��}"Nm���ۨ�����E��&��Β�ʲ�?�{ߛ���}�{ְ��aPɳ.P�H� �uH���F��-���!���F\�4�)�cy�C�e��]�]Fd}��B+!�e�͘�d;��vn�2V�@�#2�Ot�/ujH_2��Wʦ�՗ڡM���)㠆�dG�1so��٥�VL�rj��$�/5���>�+��_��j|�X�m�(���80��*/v��G����M6U� q��:)���,t����"�SIf~��TAB�V9Z,������e9^⮮�aX�t�U35&k�5b���z�i�<�Cu3�)Ɔ(��%��ե�T_,��]Gm��d��1,���nv�Q��y�Q�׃�\~-��-O�Z?���@_G��s�ͲDs�t��|��7�C�/em�C]��@~���r\@��MKH�����c��l{^��i �b{i����s��O3�7�
vf�yy��ҵ2�vfV��Z���6PV�����ǒc��l��o5�eY��k>�UU��M�;� (�� v���s+�x���xd��a*f�7oj�n���%,4���ub��+��0��	 ���F�P[�;r+p��0%����EiB*�~��/"�� Q|��)�3�5 �S�4����$��/���ݼ�g�Ar�\aأ�8.��q#e�*��g����ι[�I J����@1I`{��(p�L����x��щi�Z�=�.��r�!�)|�F�'�-��=�P��1�O��A�N�Ɨ"d��3z1a�Bt}3ƌ�>�u��>���w�(�R�r!\���*�w�:x����U����O�x�,k�<'<mw�I3��(^B���Y�������I��G���U/r�q�k-t{�gf�����Y ��n�UKa�FJE� .�f�%=!v�2�>q����j?�a[f�����&�5A�آ�lCN,&?��?O�p�&��𭡝,n�7��I��@�5C�q�|�m���=i�U��i�
ePԛy�s���!��?%1ˍ�s\��n	�Hx���Oҵr�{�ƨ�fp�VP��{��-i�v߶�fʹMl^{�
Dh����ޏ�6���&�$��ey�n;���B�ե����n��E�9ʾA�
3���VݳϧHx��t����.17~G���]Ǭ44��1gD	o��o���d����9�ct3��hyr�e��/hI��:�<�=h���H����CF��U(�je��^�����l#��^?�R@�h�x�%�(�����``��t���Lݧ�&*[>���V7Y�D.숽�xR���0Ht
@tx+����}J���B�tmB�R�(>1�%̭�|�q�\]�b���4�JI�n��Kk&����$z��jGl&V�cuuE�&d��R�dK��f�=���;tD��qŗ�fWCe�cQ̷ht^��v�J]Zx��M�[�	/_V�K"`,;��qh�>��!�f�%��_�j�³ϯ��(��U�c�!��ע�������0(�n�N����6LЏ�RȘ���hUL0F�>��ȸ�p�5�0�&��XHY��m��=�H���sj���*-�`B��tE�����1����Za��Ii&��d��*P���}��`=�#O���)���q&�O+)�M#�#R~c]PA1.�r:��ؒ�	ZL��ۂ���� ��G'�]���j�*��$�'
�}�����f
	#Q����|X�O=����l�:Ӈ=�,��e������r��iR�
���䊷�Sf�N�@9ն�$S�v�^im(q�q��
5��J�j"����;�#��]��ah[Ota/�Q�Z��|�)�H�1���@&�����%+ݵe�>� /K��di%��,��\LO�v�ٔ�{+�΃�/"����߅3)N���|�,��ąS�"?���1w�!x�P�����h��b���#��|�+��,Nnj��#,�$ɘ��	j�����	Ԝ^�
Oؕ����TEm1�B�-���6^�����+�'�	�B����[8������*�55�b���N*5X%'��2��9|�wp��d�~���9����JI�uT5��$:��!� L�sF��,��,"�����A�/7�
9�ɈL�k���z����L�2�^)ߺ�X�p	71�����[�������r�J=�|Up��$��P���]r�g�/�w��ʜFq@6g��gr�s�q-�c�>
��t�Ӏ��z��d��Ζ�$���ߕ	i��&+�k��2k!6E�I_��s;R�5Sji�~(�!�<��]ģ�-yJ�%)AޏM�Tچ��bl�(�q����w�Ĳu�؞��fp)	��j<S�#�Q��RY�6�ْ���G�&����1�g+2��q���m+E�C��D��%Ϩ�����7
n+2��T��ݸ��4�Y%�޸'��O��8XQ��\�"D ��o�%�D�g��$kL82���3Sd�x�S޳��,Y�d�j�r�K�ߜZ77���k\ޝ���}7�Ɉ(,��kO�<.��o�"��:�|<���_���^���ce�I��%^�+i����A:�n*�H
���� ������$��:L�m��L	���8��Ϊ�W�8���x� !�Z>��G�w��̆��I��еܠGJI��I?'�Q��K�}�t$i���~F�ӎ��'�e���<
���p�a-Q�H=�x�Z�� A8�G�?�Һ.�ڦ�bj��0J�)wMo� k�S������x��`4��鍿�qw���>=��Q��rٶ�l`���5JYٳQ4��'�&��/?�^�a��¶�ڱ�6�&b~3P�l�x|�nN�(X�Js���$�X��`u(�n	�+��2�}�N�j=Z�m��� �}�Q"��F�%�#c�癄y��SqE�4*�ʈ�S�r�H�@�]�Q��p�J[�����ȶ�[C�l�%�pY9#��1|x�;,�Z_��Wv�-a\T���%�0����@��ib�H.����wW�x���jM������d���Y�"�T�Ι����.
���/�g�Fݚ���B��F�C�ބ&f���,=�Ҿ���Z��h�����d%�j�P���8,M��9�=w[�ԓc��D�!"j��$�O�k7��O1~?s�Rua��}r�f���
��7T9�J�<��fm���v���X�
�'M������䌅���V�"Q�m�C@��M�H�HM�d�Rm"�lP/F2����9'Z�Rx&�k�ЀK��G��FtT������!n�����������j��4UMd��R�ׯ`����_��I�
�?�1�Ǧb�����}u�R
$c���ͪT�#RG*u��[�������|hm窊��1�C~�?q&���3���kׅ�����SK�}���yN�gO6n�x����I[H�����{��N�[��Y?��V)I���.���0S�^�>W��qX�jo`눎���E5�Mb��!�S��>f�*kԀ�ګ�N	�t�8��i�M��{8�n���n<(�1U2���,�\�~��gZC o�X:���M`]���2�����=�[.h2������G)[�'f��t�2��X��,�g�.K~�Y~�RC=���n�]xE�͍o��{}�K��#��-K.���F
JOJ%���׊����-�𤬮
�A�UŇE1k���Ga�b�,�AeO��nUU*	&�eɫ��Q�4,@o#d��X�{���H��\�o��:�o��'v��ӝ|��8āz�`ҕ��)�~C��pCdq�Wx������;g䧢�H����=��Ս��8��b�r7zd�z�zXO'�|f@P��z��2�!���+��k�	˙��bJo�-�����,{���)X8�G���}yEa��K�N$�Fˑ������!V�ϯ%T��6��~��~��P}�|������<��uA5t0��V'��s�Dry��Jގ�g��g�,]^۠��S�����f����y`H�T~�@�7.��
� ����v��n$�����(�M=�0�M{���kFm����	ά��9q�uS�m��|���TY��m'3�.���[��A� �Tp!-8?E�p�	���>a�&59��hI�.�^n��r|�WR��ᄈʫ_�;��&I��, �L0�W3�
�o^���/����V����~!�l-�H	Ù�m�T�fa�B�t_?]2�RFΨ�Bˤ �վ��n��a�������&�7�g��y�<m"H��r�	kόC"ű�Gϲ~�G���X�2��[P��_�r�X����V��ȅ��Fj���bl��BJ���:�*Hjy�I���������}��M�zZ��9?���R
�h�+"�YE�rRS��̅���"�D�}l/b�W��L�����ڑ���Zc��'�f&�&Q1�5�R��2��ݒ����ʒQ{ܠ�24G��Tw�	f/9��q鰡:��݈~^l#�o����?�f'jH֢�]o��.��BW��!;���V/�|��z]#��|(���1}�H�[2;�= ��=�@\��.��^�c.��^�T	m��= _#t �1,|&��&�yw_F��D|-��lRK�	L.���
}b�y��Q��qq�"�Þű�Ŀ��c�y򋸂N��`�p��[�M���wAM�˔�.B�'�\[i��a/&]�")��`it��䥉U�~<Q#*L����L�:;曟���fC�uE�M�rH����R:p7(��l����
�R��6/�pd�72.��Y��xuM��e�jF�V�S�{xF�_��B�2A�5	��BX��&��m��8?�M��[�Xc�,�Á���Op��(ɩ)v�6�:�c-���>�j�DW坢I| ���]����z�����v�'ȞJ�D3
e�F�c�7�|1�p�ζ��h�4O�35�1�oӗ�2p����Hу����ޟ@���oOE�pG"�>�/Y_nA�P>�æ��ءi�M%p�r¿lnúԤ֭dG�ѨS%.�Z�V�CΫ��<iq;���f~��5��!�U�����Pw�'��m�.uLR����M2�kmjeYM�8n;Θ��+�*z~��T#c����.~�������T:��a{ք�-WZ��f�1h�}R��^��J�[w����*���iY�B��7�B��ou{��Q0��_��w���w;B��9���5���9��݀��t�Xm��q�L!�Flwy�t/�n!���*@b�6����W_���9ӅO���F�	�`���ݪ�ͫԆ1@��dd\S��p�3H�� �e/�z�,��s>���WR�H�S�\�P����êji4�|�O@�L:e���V3�����M,P�c+�����ҁ��ĸS�Mܱ@��v�9G! x,�W{s_��e3�{o>�;��jT�v�6潦4#R0�E��~c����WG�~&�5|�W�~N���Y�5I�d�g�w��7P����:�v��ʨ�l���8Qr�%�
~g���z�~\FԪ(w�7���&�=�d�2×�u���hɂ�8`��c��]����hr��^�#=r5��K���q��ɶD��D�;m���E
�ح]�� PQ�Ə5S��Z2!�k�����{��MGYu��;S�vhg�o���M�Uo�s�}�	���I����fzg!6Ļ��8 ց����0A�_�{n�M:�B����YY���>p����.�GF�@�|7?����嵏߷r�{D̗-������S<��nVWo���L�f��0�,F�f���O{��L����b�д�9�r܌���#괣�*Owa��v��ϗ����	���YKQIr�R��;���PԾi�J�xg�u�t7�əʞ-��~�;'�E66��?j�P����>lǔ�'�"�,U�egr�>>m�S��6ءy��s�v�d�}�IEE�����ݿ��6Fuϕ �ZB�sHr�"�R�
VH~��.�NY�YdS�{�S<�n0.����k�*��r�v9����G��A�?�稼Ϯ���%��ȹ)ŌW��7�����s�.碎-�m3a��E�*U8|)
`P`�)-{���q!ڃڟ5�L%b�k��MwX����E����)[$�S���?���>��v���a�A'�&��]������"|���e�L�t��� |)��9��+ZV��������f�,��W.T�(���}��yQ��%d�~�|ˍy�����F����&��ק����g���� ��ɐf~:��lX�T@�A9��_pE�R���RS�IDTh���a��S�v�u�	�`E���|�x0�`y>s��Ӌ�˕\9���i���5���n��+��9!}�p�$� �E�XC���2����8g=9~�P���d  R����Ԋ�C�'�wK�+Z���/s�i$�26�������y\&���w���Y�ʐ0wA��@l�(��[�وj��x�j��N&i�Z�e�Zn�T(��0���� }}��76Gq�
呅�ŵ�B��iX���.#Bp���骮��"��mLL4�'��iq�Ҝh/;��c�� Zf$��-�q	u<����O��;�w�t)E��l�;��Ҝ�V�]2�p�=���ΕZryX�?+���A��ϳ���Ts�W>�A?�>��Ӟ������^��0�h�u��-ZV�FBɶn�F�	��;5��L<�Z������`j�J[�0���%j��Ruu��	Tژ��Z\��h۷O���8���a�~�	N�K�i_��eMx��6�l�UV"�%ë����w��@F���`i0�J�2ֺ����P��8���*K-�0aD�T[C��o�j��&����,��~�D�C�_N�sY�焋i��{�aS�u�eYjmB� ]]Է���V�=$��f��#eE��0���˰uW9V��{NQBռ���j���V5_ {�*$��,cK���5=�o��f��O�ŉ���\�

����ڳ#iδ���`�U�h��*�٦e�YX'��m��! f#�*O-i.��8��:3�X�%x���"Af-����  q�W��i�SM���9��/��U���wh�<��\ʄ�zP@w=?��v2��N�	Qp:����(����Q��(^��� �th��������E���<�F�C�=(�P8Z�~:�P��S�bs��i�2"��@=j���-���!�|5��Ъ8��K�(���\��*[���T�����7�=ȩѼ�XğF�γ�K�{�4d�� H
��R�g�����'O���R�rT����Zu����|���W��p�W<�F�,���-1}A)Ũ�J�] �geԶ�O<aM�35���r`���ǌZ�K����tvdQ�-�I]{NO�v�<1o������E̵���I��B�����Z�^���ZHk�O�x��3R9�6����ʫѹA�pA���
6�1��`�IBN+cNqeB;�P3�ʋ6��ry
("����_�a�����
��j���(��� �UhZm�0�.78'/�{y��
����&=y�w\Ib�ȱ�����Fb^uÈuR���Z,�"��s��L�Xĺ����4��E�8Qb;v�6�ňj�ҡ���	1�U(iDJ"�n�j��[U�Jl6���:��O>�����Ѻ{G}>��o�K˘99��g{C��%�7��`NǊ���"p%���?���Y.o��d
��� �w����
/T�g�u�S��@9v>X�����<����<�;rk��s�����g'�2a�L)��ԹZ j��M�M�%�5��:��JѰl`���=���>�F V(^+����yn��xfE���H6uq�58澄�Հ�s��k}jvgdm|���»�7�vn���~{���";�kDQ��To I�*;��|�ʟ_C�d�P�$V��5�r�R%cʜA��!]��&�-�*����1A�c��n���͚��f:J��#��+�i���"(�}:.x_��nͭ�t��׫V��?qA��w��P>�X�"ĸ�/��ֱ#!��uǟ��P'_�c=�CF�rd[�EZ�|�8�����{��13�F�鿸
E_��U0.u���b�ˉ���L��r��݊�^�ڴ�6�Q"WJE�����d��\��d�jO��S�v�&a���Mk]�t�GR�^b�G7{6�*��<x�RT$jT�� �#�{���Z�9fr%���w�k)�U�2e��2��$\���T`1f�	�z>g���<'TB?���2����G6D�����A��4�M������ ����yfm��1I�	�3�[��a��1��N��cy�m�!��|���7͒�����t}����1I��s"�D�!gd�ksY]���c��N��3�Z2��K�\�R���� 6/� �zF�^[����&.A�'+���	Җ9-��`��C�����mR����� ��,Ei+Ｏ(���Vye+�1	��s��� Kk���
�M^���^�����T�!犗�CF��>�����[9u��9��[����iW�*<C���h��>C����C6ަ��@0{����GgJk&���{L�~��)�����l�7�"Xr����љw��|�?���G:�&�N�uX��v4C-�U3��%t�p�/�v����j!�Aس�}9��:t��1"5.%_Yl�
���	�6,9����\�~��Y�{T~��W`���S�#�0&�6�����cu�BY*��pVX�M��#l�b��Ҕ|[�|b>�Q�OkC~H�.nz��K�BEf��O���<�.�?��dr��Iv���z?#�D)�}��� {�g��o���;���bq��H�bq��������4O9NQ��^,2"�k�{3L|��Ѝf]��8��QKPt�\ח��"r������W"��I��IBx�B,;�΀�I�qUe�b����������g��f�mL�L�pxQR��p�iƌ'�:w�LO*r���@��9v�?�Q,��@����w��`zl
J��^�Q�7�Ө^(�'��ֳ�i1IUy)�O�3�����Q]�����2��gȦ8�T� ��Rc2����u���*�t��.�\kHLɥ>y�� ��\�:ר�UH�0l�M�<�b��ˍ"����'��\�Vy �k�����t�O��JU\C��:����7�-��e�\M3���@�S��ŷ�}���Nǳ�V�"tO�d�?L�2=*��ѧ�7^�?al�K�fƪmA�xY��w�D�H�zov��N�gғ���i�*�XY8��ى�.��b�M��M��I{�u��
<Q�]2����x`urP8�_�nGnH7�c<�bzPow�
M�����L����w8k��?~-7r�M�S�~�9[Q]|��ބ��`�R�'w�4ǫ� ���E�xx�CZ�8h�O�ρ���֦,H�����DI�~��$l����$��)��}����<�
=�v���Rl�����@�o@�ٽ.U3ʸ����g4�_尟���I�Xd�ΰ�&�%a�X4(�>��=��GKL�2�~�9􋬥cP��nғZ6TC�h���ةM�j�����Bcܞ$�]�|�~�D�$$�J��}���Q���T�'��Y�؂��,hZpv�i�h55��B�e��l��v�7�`)��k_���C�ߍ� ��˦�:[�����>�
-�_�g�����9�'E�J)�8%G�����7&<&��<�V�?D�̀���Jtؤ�ڮu��i�Z�t{��TK(����T|%������^��ؼ_��6�Ab����tW��Ht5i�2�5�?��W�j�y�U0��G���7Y��u �Dqކ��9g!�/
��2tA�o	o���$u�2�+����a�#���2�1c�@���[�ʅ�J�ş '����z�Z$#���Ƅ��@��^T���E�;��za�;�ڨ�A���?yb����m�RS�N�M�&Jy��,s�ѽ���-�#j�%g#�i�1&�Yh��c�v��	L����S�ڥ��Q���Z:(�qg�}���l�^m0����	���n��1$+>*ݫ>���
��Z��V����H�ͬҌj�B��f�����8�l��W'�z ���+�\����Θ[�%�@+���P��7O��(t�C^��:�3��"G���.B���j��]m2�?j�-�Vn���U>�v�0�#�;t8�H��ri��x�.�\��9iO���Z�4�Z��	��	�qԲ"���Q�A��dd�b��h'Ο����V�LNf�|�{�{K�F��1m3���=,2���r ��ٌ�P@�p�*����J�4��@�������������E�����ڧ7���a"S�X�Fhǘ��qD�O;��&��"Ylf]��Ô�|%@Bs�i����͑���ܦ�f:f�ֵ�9�Zl3[DA��7� y���ӹ)�4�K��z�u�k�Q�P3���C�q��颈��J�F�F+g	��>1ԊK���}52փ���KDi�*��<�e��!��%2ّ1��(3��	��tIUK�rq���b.�C��>rՍ^>]�m99j� }��#�8����m��5B�To}����Ω���
�`ů��*l̂!�x�ͥb�����m��5�i�Q#2�|��Z�s"{�+�����w��^�2�ԋ���4��{˶�E�ɮ��iRv�0���}�߅m�#^��Ap#Z���B8��o���ۺ��>)C{a��J$���.kK�Hc	
C�0З�,���$$���M��Zk�>���7��| $�W���O�Ҽ����Z#���J�����@~T��P��-"ؒ�p�����iV��;7��ac9�%)}$���^m@a���3g�=1G��8��g�]���_��
�i�Q��\(sQ��צ��\��U>�[x�@D�;�(I���"��v`�7�C�_��~d����<��f�H�P�(�:�T�#e2h��U�����2��B_�0�P&���+8���')��S�SP�U$�	ҝO�Z�i��cW�ǳ��݋%����_g�y@<��C���3{���ʁ��W�;U��XZ��֬�^�D�ڶ��?i��rq�Irk����:���K:� �7ִ�6o%�cq�Ey��=�r'�( �n��h�;N.Ж?$\�I��wݮ�y�t�i���k��@0�u6W��E^*�q��\��.�V:�)�>ߏ~�B�hDhΘ�5)^�g�:��N�]#t�;\uq��	Rk%h��x���j���d�Z�2ɀӝ8��Ԧ���i�&��\�wY��g��Ȱ��qu�p�*95�V_GH�'���ŀqb���v-[�i��J9ch_�y�5��=��^�j���}�z?"t1�1Hf&�h�<6f��AŌ9q���ظj���F��oi�B��eR���+{�� bUdj��cL����ɐ�Gm������iI{�|���Kp@E�����i���84�>��H�x�:qP�zV��- ��#\��k�F#'�3c �H��Z1n�=V��8���)��[���h ^�E4Y&��H�c�w�����q��M�A�A1���������Θ��5�43x�4��l�:ޔFT��3}�Z��:9n�r�y<���v�� ��T`��aL�Cb�l��np�'���[E�	]?,q.~�g�6C�������xFQ ����5
:�5P��-e�������[��]i\~���f���w�����<�x%�� ������H�{��P �W��;sNy��&j���j\% ��(��fT��?�V��Ev�Gږ�2W�x�7)o(b6�I�K��ᛲ2��?�[:x�����Qn\i�"�"��F׷7%�d��7L&x,�#�l��E���G�?4މd���Z�Z�L=i�hws�]{�v������5�b�]�a0x��B�sմFH��6-�����x��U<sC����ǁ�.TIO�X��T��%ݭ3 Wq0�?����n�s&�D;�G<�,�IL��2,I^i&����2���G�9Do�j��[��(��;��[�]�R�y�Nj�z��u�wt��RKL������+��Lr�V�T�����&��Nc�|���b,Q���0�S=V��_�L���e2<�To�f���<GO�y���j�-4�}�ׅ +�����괾��y�����0�b<N��v�`Q�����^�'�F
����AO�7�Y�F��nסN2��.Բ[���MW�@5���;1������Rt��u��+���J��3����l6]����x)��J���w�x)�~�^K�M�cG��C��Sr&�ɖ��:�"|�թ_���6�r���6[%�"k�p�1�Zh4���&��H�<�s[���(�C��k+�O�,0U����L����9 ��C�m]E��Y�K?�|�I�TKY�7�1(�qb
�E�+����Àr���;vmx*���ɆUͰ�My�����k#9�>���9�Z���@%��;�S���Y-շbd�9��m�WOb7Pf�����dqR�Pֱ"�A�5�l^ʒ���I����Q�kk"0Fq�Ǎrwb��z}-P�7t�%K,��7(Dʭy����3��[��5����/J%�K���o+�S�t*�v�h� ^�T�x�o64$���Q�^�1��^0��/2�Y=L�lvm�ڱ��0lH5�P_Ve�e�=�K��.N���n#�Zx���&��y����F^��du��̽��\��PR~ʱ��`�?s&�������&hl�V��~�=,��-�	9EݑSvk�̍�F(�mwK!�n�80�kE1��4r:_pZ$����
�[�?�%}�yc�@�5����I���wpD%{�\�)������O�V�Rޒ�ף+/S{�RXMy3�"�u%'֝���v<�8��E�f��u?h~j��a�5�
�j�i��5U:��jA8Sd��92���̳ek�:�WV���H&��}�M*�:d��JS�-d��#^C�;��w�V�v(�EB�=��!�6wCI�C����4�`�̏T�Ó}�td��$N<�3q�!ؐS\l��?���B�KǺ&9�ť�$��b��0Ecӯ��x�Z+����>ު�Ӆ����� ��d�!���������W-����T��L��,�� ��7Ä���n�aIhkP��c|3��֛�㊾3ewa0�V�s�0��D�t��.l�ٛ�����U�[�{V�;�pn���`|]�׵�,���!駶��g�hN�<�7�(%Bv���(�<p7�$L��<l�^�6�ي|,��k���%��m D�M�[/���˧!�uM������0 )SUS
�Tu�TG�q4��EF��4���PKE���9r^0�������c����bZI\�|Q�
9�, ˚aU�L�U�=�UK]׹�Z0j�^�yDz1و�9�O���t��x��>o����;���$�X��MW5/�̘�Z���0ݛ�'jvuŅ��tN	��dN����w^x�diӄ��v?�����}�=Ӟp��	Giԡ��k��{cB�D�6�$1��~h(gȄk�)bO�v�-n�~6�Y�2N>ɍ��V4t(z����=�!�4w��KHԶ[�WTF\Ѵ���S(e��u]U�u���Q{u)E��1)�|���a1(�՝�F��Nwj����˅&���OhHd6ɖ��TaX��*�g
7v���؞�(��U���BY�2�壣�Ef��������׮3�|�x��R%�9]���5&
��ȡ:�a���F}����Hu#EOKy;��.~�����:ݵV�<8R���}%Օ���y�,7җ�w���`��/|1�~;5;����+��v�F5�O|�yx2�&���͜��ǍS��z�D <���HL��f�$.S[1�ETA���V�E��g<�t�{���	Ņbh
�*���B�5O�^��fK��~��<{�:�^,��v�RJ�P��$2@���vA�ݙ��^\����6�M��#����(=]�.�T�K�h\{Ů��P��H1F`/���B)(3T���+rk��w6�죤U��
�_H8+b�@RT�%�Xga�ϊ�G�W"�&Kz�B���u(U�~n ��e�<��^1\��,\����UOo�3E9�n��Z9����=�A?�"����5��5�~�m/5���p���aQ�<�n�b҃��������7��B��c���Ɛ���6���f�@���6+��l��8z��<ӎ*��{(	�`�S䏈F�I%T�^� \�Y>R��^�;$v�A%��U���X�S�܄��T=��A{x�l�����3��g{m��WY��:�T�9g�Pm�{�{q���ڏ���o�LR��RJp�Fm܉$��g�g�X\����׭[��8؅�.a�ڀ?�,u���?�)�i�4���<ޢh�{��V�$9�w\M�m��)�R 3<jݑ�������b����񣃦�L�
���oY3t���@Aa�8�>�r?����b0�>�wY��|��w,j'�h�s�[�JV�D�ٟ/Ͻ�k����ՑY0��X��n��8�5��匲�%˪$n*�|"18��]˵@�ջG��Oc��@��q)ݍ� a�{j�XA�˃�3�z�
��R��R}1J�V�L�	O1��PoSbFҿ��>l��Ԥ�Z�Z��D8��es�1�J���^ge��e�q"����M�G��ݮ5�Zɯ>�4��&�L��"a���r��5�2���J/�Ve������q���YD��x�h��z�96�����ul�!�*��|,�	����dI����ඥ������}_p��7�bY6*���0�5�o1�!;� ��U�R�S����E�h��m7:��Z�n��{�(�=��i&S��(8T-�?�Ϳ�9/�؟�@�ws*�I�f`G���X�cw8+���՛�ٛ���o%!"s����#I�z$���m� �������9OơQ]4��yJ3ş!�4tv�6��.�ǙO�1X��Y����g��f�J�Q/b���%�͜�!�=��b#���5��8 +�BlU㽊����4O�F{��˻K�Gf+,yY�U��2�p�&��*Q�:�\�W4��<�@>e�2�|��~�.�Ry��4�i���q�a��}r(D�վ:s�}�3��ŏ�Ɍũ��j��v�:ލ>�^_���f��'Q|���]�ַ���)���mg��auΊ�⋴a��RA琚4)X`)b`�=�HE,^��z�n�����_�L���%���l��#{��l>O��� K�8CM�1*L�l�YG"�'��g����W����/%�{��2�Z�Hq����l����F�rh�+�M�m�Ь:K�����P�%�����fZ<ᧀH��0�����o]Oob���d���g�i���O0�/c/p=?�RX�7P×ɉ�ª2����`I�V9o��r�V)�yLq0��@�~�@�q������$������ �//��O�T���/~�!;�}�aaE (uT?�67w�������Z�4���.j��Ž�^i'7�O}�/5��%$WumZ�:�f�f�=A݋����T�D˺!�<�er�Eķ]l�D>"O��6�[*�������D4�兩�)Z�N<t�w��E<\��ͩ'��j\�Ok�M����=9I �&`��&4ۘu�r�)s��"�+�W���'C�k[�9&j/�tq��i?115�[k�!r�S�Sns>�BmZ������Ɓpri.���'��Z#�J�*��@��b�>��T0�vϫ�x[P�V�������ա]Ī�%��B+���'��$��Cj,�r���j��drƯ�����<�x�b�F��V�Ri2�r��4����h�����T_0/�X�C8���S�`��+�X���:�<�E�/�L��2�fQ�Y�0�Ұ+=G �C����oab�j�S�}Ie��W�̀�<�+��Ed�.�~�� #�2hK�Շɂ����I�,��-��W�X0�c�t��__'��U��H?��g��s�D�Z�e#��Ya�v������������r�:��	g���"�$ -��ܬF����u�{O��%�m�����A�%}D`��p�����k��r�����nÖw�x�O�|���R�*���������>؈�H�L�U2poL��O-���?۽�Z���瑖�=ٹ�e�8�p��.lo@XD���z-yXA�u��Uk0)s��M?�2,�G��ǔ١6�2��iIo\.�<�=I����=� .����]a"LA�|�KL�@��`�4\�yYvSښ!½��]��2�	��H�z�
�����M,9%J٭�Z�[nqʎ�W������$��*R]�����=)Kmv�T���Wlfp��D��,D$��"�?_����,�d���VQ��B��~:� ��)p:�$�ET�x��ǅ�X���~�1&�� d���uM��{��Ҷ�����~@gRӝX�=�BvĖ~k�W^�s�s�E���G�^A�f�zD_��Oy�l���:�=�I@qKk; �T*b{�`��,��0��=6���p�-e:;Q՘i��2�6��FH��uU,1��(��ij	S%yX�%�lE�o��|pO.�h����\c��B�2C)���Pyb�3����72��&C�>���IF��䐙���J@���\�bb��]�ew�K�`|��q�#��&�t}5�ƼN�'zFeؤ������a�6(0D�	�"���`�R����Ϡ��X��LȦ��V�uX:\�(@3��F��o�����t�E�=�F��=i��b�"�13�AY��Lm�j|6@W����R�t3�[��ʷ?�[Kt���;oש�� ��kȋڪ���$ϼ4w���@[��1N�V�/c�4���T!�>v]����=ԡ��[�H�w���7��xv�JSI�K�C�~�q������s	�퟉��X�P{�30���)��_���F;��Ó� CdG�8b[��B�-��.���$��UV��(����E���V��׋��[��v� 	�}pR���A��7��Z�T�`޲��{�8�*��s"�;O���c3c�g�ve��1i�]b\ehkv�2AvyW�����B7�9�#H��ڠ˨D�6@fr6)(�z�����9
$:����=������A��A17�w����.N$]�I@������ ���G#q����O�n�Yi�%&�b!`-���խ�nC�
�\y����l�5��{��~����)"t{K���^pBҴ7%W]]y� �k�g��yr�S���	�i�x�eh6F<-c�u�݋X ���I�:��
�����M}�=L���-�ڤ�[���>~Z`�o�G���'v�#��J�zR,�@C���t��i�`q*�g殜��L�(��z��32�Gr�:��;
�)&�V�ó
�������nhp^"[B�X��p[�i޽�uNF�U#���<ȿߧ��S~o����yU�鱿���j�y�n��TffJ腾�Iw�_R�f�aq�ȂM�d#٩�����WR4��i)X�Y����1�kD��K�D[%�qp��)��M!갉�tfЩa�ƴ�&�zL��zA|��E �}l�h�[����:So��hvĹ����n0QO��`����H�:�v��q�leA���B��-�0���X#E�i�}�84,ƙ�����;�)*iT#y�@�E�dV�(��*bhS�#�h��~��AC�'���hA�x�2��<��O!���)���m(�y6І���n����^�I߻�SB���5r�ܽGB���N\-\���AF��r�C�k�9�V�s}g�l�"W΍�Q1�_&.����{��s;?:G*���(f��0|����l�&6=���6��P)��,�k�������Us/(/���1v�~s?:��ӬHK�H��:H�ʾ7I�dn����K������߷�<��.s�rQ��]:���j�&>R�r�Oa����M���Z&2�]q��$��n�8�{g7�:�����J�Q�/�_� �c!��x�C�s���94z�5n#��q�:Fr�7�<)�W>���&*�rs���
>���	i��� d`>Cʷ��k�@x)��� &CS
b'��πm����rR-J��^�܄��H��u~����p�-"W�:��w�` تV˩�Rq,�I�Ac�p��؏RP.���W��esl���u�;g�ɭ����C%�"�"����A�	"D+}�����Ⓢe����$���-�9<Q���@���B����{��{jT����2wr��:-<0��Z��ՖR�fW��1�A$j�_�9�KߕV�f��t���B@tP,���]J�UC`�I����H
a�:",_�Nk2k�(�~U-�o��Y����h<;�@O��a����p������A�<�Vñ������U�m�'�y����6���x��~#�z�{�͔e�;����k��S�����r��Bqj�Pqʩϲy�����jc��}<��Ɋ*@e��P݁�ь�2���
T=�
�I��<:mL�,�~ɷP�7K���=:�/���7[�����!��Y/�0M�J:��=��	@�T%<����{�&��_��#Uڥ8TJ�u��m[�li��9�ˆ�����0�+ M��ś�y ��6� h@9��t��9�D�%p��D�����T!�ef~�ZI�Wc��1���$����/��`�oh�o�{�od_�T��vh��"ֺm�f��)Y�eu)vo��륍Y��XO�^����w(_����l��7�x�����.E]I����!�a'�=>�KWꂛ�$MI�j	�00��H*�tE8Tk���VL��:<�����=�m���l^��1�Te����S���孂����9���z�a�[��\F:�@�[���Z�%�z�Ot���胒�.�)�'HX��^��E]#�ܔ�A��d�.g�S��#Q\�g[
��_*��45N�F'}�(�*�V�KU�칫'��a�t�1ט 9� �m�c������t�XO���(�����,���
ns/S����J�oΊ}�~�+�߰�����	G��{�������!�֣��#^Cǥ

C�gx�М~�>L3�71	��
;�h����s�O����%]�p����#&�u�����㘁瞆�(��_5?�g��s��O�F|��ڢ3�e��bӊ.�{�MZ���y��G�OX�`�'A|f���|�8���Z3�v��6���q� r}�d4G�:�%�i�
�.�o�d��a)�]�$Z0��'p��.3@�MIV��H��|Ԏʫ�V�L�J�B��CSBů3���݌?�Z�A,�9_�_F�`JJ�HP#J@*4Aj����j��u$�N����Mo�"��o��Pq��$H���_�V�+��!%c�l�l��N�ͣ۬c�����A�k\5�0Q���K�����+e��٭$����g���lR�=2�B�e��l�������*�s+��^�S��3+i�6��}�;��x�6//f�p����x}g�b+���v|#A<�uh�r��
 
D�~ᎴsI���Tŏ�����X(�-��J�n�x��'
��5�XIz�����x�t�\=����B��>9i���zk�l�C2�|Ъ.g�f�n�r��5�fNr�$D��6g�XOL92:(ފ�'Ox�r~E����E���}�a�����bGo��VgMu?���b`ȫ-��D.��o��������tX`K���=�A5?�®u�Hע�j�>rļ��%v2b��?�����0�c��DֶT�h�@���IF�9m�}B��A����e����I�nn��/���ˍ���H`H;"=�"�[cJZ�@�nV�0f2U�9�e���K���V*�f̌�b��k`�X�!�Ꮱ���+�n�'�HX�c2�Jʀs,�oIǊ��{pu;�:�|*7�Jo*�.C8� �Dm���m�/W*V(*?�2��:�$�����B���ݡ�e�0t��Q����V��\����WT�c��"OwF��e]l�'��[����(����_���mb�L+�Xy`�A���	8�E���C���2C�����nx"����G��+G|�xy")������1&Lh]��m��g���cc;]]�z��{��/,�z_K���+�c-��׈�ʼn�#2�%��Z�����`ݱP�����������DЮό�YQ�Q�ꡛ���i�>���R�<�?�����DkP"�� ���a�t.�/3�۱��-|�\��0�|���0ɯ���q�~�!_���ȳ��e�i���T!1L�8X��@15�T�(u�D��Zaro(&|Js~����1	��aщ��<��I� ��d�m�DW~>���cY�樈�ʡ^�v���|� g��EWm?QG�S�,F�b8�N?�"�H�(*����ͷ�DC\�}�.E8�0����;cW�����q�3h�l��[&lk�k��H/��$�Q�(s��KT�L'=�(�Vs�pbr!b��d��Rrn��k8-7�Wz?��M�a����j�K��;i�ug��ҕ�J�
�T(�IF@���Ve*���-wٕck�'���/�"���+�@�mT���\����[1�����h���A�H���3R���6�h�PҾ���g���`3q�HtE�uчB-rr!I2��]�Vp/CQEJܪ���=	���<-�Q ��%��{���N��[�pD���'�#�Y9�/��
6�ckO�#�/֑�/�\?��������)�����ש��` N=��j�^Tl���8e���ICk��6�_O;V<��*�Ƴ�3 �f�d�u�;���U��]2�t����p�� ��+z�&�ڞ>�q$�cgM����
�����s�W������U�;G��kuaN�7����'�\g�i��Pt� �iE� S�{z:P6�YԮ�N2/ɫ���b!�	��$�I�t9�ϴQc��B���Ԥ�E���k鬫��,��;bD_ն��9,��i�Ͷ�}EX�'�<�]<yZ�����b��j�Hz%�j5qda�̮��2 �`0�#4���1����� �v�NA�xFw�y��/,�h>����9���A�Np���䖄#%��(y�4�PB���3u��Xl�/�(��3��V��JQc��1�L)i�r�v�U�AƼ�]x�,ᕠ��4 ǶqS�z#]a
_k�~6]�^׊1��O��>��7-/�
.�z�b�eZL������/�p��a2wﲾh��^`d�Ы�W۠�`F�	�h7]��M�y��">�#n,y��B�|PB�114,��Mj2!j㭧�8�`jP+c�@�o2q	e�iz���FݑF������T>u-�uO�,h�.]���rB��k��Jv�`�#6��7�N� ����$��JG��id߮�e�a���kj��l�ų�"�\��e��y�#�:�4-���*�F�:6���U�}�����Z�yu���_.0M�5� ��>g�c}����ӊhmo_'2T��Q�u�&�.e�^�uD���#�N�k7`w�U��x��l޻��dtѯ�VޫO�#I�L�!X)L��oz�TZO����f�Ī�C,}��}�\�p�$�Z[S���7=4֖}�<*OP���(��#v/��*�`b,��;����rp�K>@���_��{v���f���J�K9�v�A5._���_kj�Ӑ�*�g��륦�c��Ca��47AS'rȼ b,�3n"�����
~][ʩ�偞��U#}����W�.��2�B3�/�@`�p�&�?>�#��ŝV5�-���ۆ&H�~}s>l�N_���R�u�t49�P�qv�?^�2��ָb%�z̡2��t��ow��n���/Mx=܏��~u�E����Y����f�t�Tү�����͍��Yq����=�es6ถ�Z�i��s?<It<�s�$��z�8l��%0��	����\T����P3[�N��XY��a84��©���J��Ȓ �ԙ��ϻфu�7-���
�^��yWj���FT-��rC����a7�}=<������s����+�
y��x^���T��*�Y�Mg}�dn���EpY��?�����W�aꖋ��L�NԐ�s��w��u��%~�#
���	��Hl��]�>�^g��|pm�ױ��+)l�:�垳(�W7�Fq�#���E�N��P.�k^:�m�5}T�mu��=텍	�b�����T!�uw���uCo�2!ֱT�fh��#� L�����X�󑉄�����0f=� �Y�9�3��?��kA�-��Hy���5��X�2�	OOQZ�#:p�ټ��cJ�m'�wj��m� /k�<��{N�3�tN��S�����9J�XZ}Y�9$6Y-����؏�l�e��~�Γ���3�ğ��$��ݧ�3b��0s�ޒ��I�ԑ96���aM��VU#���)���!>�V�@Ә�ذE\��D��B=%���L���o��:B�2ױX�Wa�_�JQ�x0�uҶ$�ɼ�H#,<O���ajf���E�B���xe�/E�V�Ƴ��7ؾ0����&����6��ȲI�\�z�x���X�s(sc/��`i� �����t*{k��2���R�ѿ!�E�n"V���K�9^-�����uF��+�+&O������ߪW��@�7w�X~�O�o�>�|W�K�P�[(��(�"�>.�i=ԕ���������U�z��(�uݩ�}���v3ST�}X��"_?SP�+9U��}6�Ъ��iF�$oe� �st�s�>y�Ҏe{�,��qt�gU�:��
�&��Ưת9�SV]�� E3]����H3�O!�6�)�O���]N`���Cs�����S��v��>�O?��kNx����T�脧.?*�ġ@�X�v̅#g4sn&M� FPR�v<%-!ss)P&��j��;�OH��T�{���ڦ٢2����J$ �XV��hd��Gx����m�W��7�T�X�W�+fi�
��e�L%���i;����i��e��H�����䦥�^olb�&�f��dp��:p���^��pl�N��R>
�pk�T,t�OC}5Z��7���%4�	k,d��M�S��3a�]��l.u.�ZA��$�%V]��#,r�;Iw��f
|�g�g�W��ԔW�]jE��裾2�*����7Weԅ���{�	o�z�����P��b���T���G<Ѫ;��)�"v������׀̪� YAQIH�ħjj+ܝ���]���|�j_\}k�U�߆Cl�T�AT��E���Ej;�=hO�wg�}�	��	��+��C�?��}�^�Њ�uY�Į´�D`en�ɽ4K������0��A!��xf�5��\����p	8� �|�x�����/�9-ϙRӫe�rIq����in�,��T��x���806��h#>�f���,W�<Fdm-7�x�b0��y������d2\��"4i�uæ�L!C$E�V�`WA5ϳ��?����O�IIu�8�[t�h�x��sX�f�o%�y���/��ߨ��|��P�9�}z#{�A�6�Ϝ	)�l���5��B�`�|$ ��Hqn��EQ���fὕ��АB:p_Ǹ��,
>�X�j���5��ځ"6>h����-j��&�ݯ���|#v���!����5��/������o����U�L��T�n]���f�o��u���m��o��ӻp��3���sG)ĕ�X}�A�ϑd�ׯ����1����h���׌�xf�C�T��� �m�]�%�h���9;?���&i���Lc�D��I1)M�}�_��Ą=&a���cHv���垗�5:��C�yI����hD.����&����Ë���X$Ҙ(� y�jaS��|�g�-��''}%{�G���9$�3=�����x�c0���;}�Ͱ��
Z<x?M �sQ�h�o�C��d��{Wq�=o�^P~b��P]	'Vey[5g@B,kɘ53SI.�$h����'YN��9��G]�c�E/�jjNd��UR����ї� �\);���>����Y����ȯ�h�Õ�r>�>X�W$��-��h�Ve
,OX���G�-�x�i��u�.0��{L6��;�bs[FG'����5�'$8#'��!��\^8 s�TM|)��/@�)3"-���3J��g9���Ɯ�̬�y�n�n�46��mxEY��A�G�#_kU"d��>)!�c���|X�D�Q��|[��k�iȸ4,	�6����S��@�e#�W������ȆT�	�go�������/	q��:�>�ޮ��A�(CR*c�\'�H���U�;����c�u�>[��G����� �����'q.��(l|(���X�H@u�C�4���rzM)�)�Ϳ�';DnO�U{���{��6�~ըx�3�@!�r�`\.�U~j�*�7��T�S��F�ߪ
9^��>`��*wq��0`�p�
74�k�oG�����_����~$Z(��������s�;�� ��7��ľ���3��ؙU�6F�&���u�%��5f[dl��"���u�2:
�%��t�ͯ�t����?���Ǡ��Ʀ6R���oM�%��wX�����F��!�4FP҃�x_e=Ivz[WN�Jq��T���A0o����8�3�ȇDVA=���I�'�{�#��tg� �=����8������ޏ�O��J��;40����� ���A
�P�	�]��"X"`���>�cT����{e}~�qU������~��������^Va����Avo�KA�!7����Q�\�ˡ��&k^��{F��	팮C�8�I�<�V���f	`�~�H�t�u��G��>�Vٵ�������m'è�����(&�!�"{�Ϣ<��@���L0�
�к�6��!��SJ�"��۲#Dm�yAQ��������-��U�޼��x@F�>���_���`���:�zH��7B♯�
�&������C��X�I-��@��B5�]X����:�T羶Ҋ������f�A=�^>i�0�*5�I�폌����h�>hO�m ��r�D���)�S��옄�kS������~4m�R�(+�bæ��)a�06U���^^�s�ڶG Yh�B)�f���>�D�0����p�͝���=�,QUj�mC��������aB}6յ�biz%�޲TT�s~���$*G���#}�$�q��\W�^l�I�oq�:����?��g#�p`�s"�H٠��oI$���뚘�<��@cuܪ9�f����[C=������� �L��H��b[�iJP��_o�n���&�㊸'�[��qoOcFѩ�c�Ҏ�z���>�0�g���^w�pbު)�v^w�\���W�����)۵D��n�V1�\�H@��c,�6�l W��\M�����q��(]��$1�9�)�	O�1i�a]���?�,������j�I~����oߔj��T�{���T�2��� �ўV�R��K�NU��;�L���_)�3��|��R�7��mʇC��833<�N?9���f��6��O��O�N�ɺ�O��Q)Ϭ�e�A���O�&}�Z7�"z��c��c��*k���O��Zժ�'\A�Gh�t�s�D`��1�0��� P{4�M���Zo�����~����P�7ϖ�IySb�r�P�w�(�7f7�ё���H�r���Ey��R�n\t�!6d%�,���M�K&,�cS`�^P�ZcI�eI�J#Mx�'�fRԠ�w8G�Y��<���B|1�����XC�y�m������S��Q�i�E��Gb�⩁ϓ�'Qk,z�jD�i6;�D�b�o!;���HX��q����@�6kT��<r�!>|����X�JJ+P���|���o�&Y<��cD<�n�$V�y��vK�$�3Ն��ByS��e��v��O��L�2���|�� ��uS,�$��Ƥ��W��,U���������^��+c�s���(�����+h5 1���9��8B(�mN\�����Jn�Q����o4J~��n�D,wKY�NC8��F^��fҘ���,v� Wk({����np��ț�d��7��zQ��?E�>C5 ���E4��jo��^�����
(E�d4⦇l8+R:��_��p��`n�[���Uf(��\6�{�bC.��u$�@��H��]�\�w`�`S�Y��:H���E#���L�����8KR��:�6��L ۉ�Yլf�M��cˮ����(�?-X�I�l/S˕��5O3�Eo����(CM9 KTK�i(5i��X9 �^�6Tn��C���g-��_�.dJq���6S�F 'EV�� zmT����W���lG�5�����A}E�G��ld�`��	��%w�7��*��oF���M�a�ZH���M����u���V@uG�/�0�lFfi�����r!E��/�'L8��fH8+��5�
4l+��n�s��w�¯�":�j����$~�[']ī\�eZ��%����t�xr36j�dP����ܢ�A�8�a��}W�bC��`p��!�=�����P���ТuͿ��0���},3���=P�c�ކ�:��8R0%}�!2>��Ń��`��^2�I8A�ӣ;��_dvz�����Ycn�A^i#���߿��L�\����{��c�㦬xE(Jܝ`	I0_�VN�Iq��]�T�]F~
��=,�m!6ljP��XϱK[�fҬ?JO:c0S3ʶ6�{��r�������WG��斴T�=�Q>��ʹ}�L����h0�8�\W�UA7u߂�7�p�J'��X�����_����d��X�8[n�m�6�n��gw9+*��=B���4�}�(2�~��
a�PL�մ��\;�6��@�|s��c�q�T�?�.o`+:?����R�º���e�;!X����5{r�!���Fі+}-�����V��2Ê�-G��bv��mi~��9d��v����8B�z/�/,���`35c˵�T
�Q��K�D�g5��⯌3�#�����u{����O�D�B&j�݇UX`+͚j���A�箴G��Ʉ��/]��1VPh_�kc��MG�/���cJ?��h���� ��
���7��@�B�ٰ��;x�lkw�d�~+tuT��O��`?� ��R�=ۀ�{]Z9�i���l��"(�1�u��!�V]̃��������¡/a&��VKrH�����L<L{?��������R��SK�d����D\;y�5eʼ+�Ư�j�!}���b�f�(�u�f�%�F,P^~��z�;ާ�R���o�߯!�C.N\��4�%�|!���WW��k�pI���ϑ��E�]��e�9۶G�`�d�3�B�kY��J%�����l�@՝�VK/��)E�6�x��MU
u	.�'e��"*�vǍ+�#<�^)���<c��;���d�4���.��GN����@T2�*�a,��h��O��"�|�ݕ,޴��H��x��3ؤ����MFhB�>Jw��|iK���0�e"Ǫ�^��eu!����pv[�Q�ݾ�)zJ���)��$����x�@v��{�Vb�P�ԋ�����9:19w�TcVô������J�3y�&���X��pO�7:�ԠM�I��t� �V����<[Ȗ�fg6y���*�f\Ԟ�8`ɠ�&��h����#A�a���u���ʕ��?Q��T��B��
��i��¨�`�p�2i���U��9	�[�}M,��Wڨ�l��_!k�7).���<ŉ֧�j��#Ձ /�ߟO�1.���=�]&�r8������U����ۯ(?��"#�|�4�-��*e���D��;�o�@��y�������?�~A&��]&�c@Fz��O�#h�1{�zr
�����}h/ �#��V�`�t�Ѧ��B�ba3f�'��}��n�k�덳�gք�d`u�>�F/j�vJ!�ږ@�9�V����S�#�J��)1?u1�g�V��Pdx�R���ڍ�wo�����6ʤ�^�L��%�J�B�9옧q���%5�T(_�A����$k��F�/;.|�z)���O���1ѩߝ�ܲC��7ˇF\��m�!Q��(��`�j���\���Y��E�.F�>jЗ` 0E:�KI?*X0�_�	/�EP��ݡ$?�j0&�f�&��u8x�iUf,꽮�@m]5HX?Qg������UԿ��xD �1Ot����|�y�:?�6/K�S&���1��*����������%�-T /��N��j��w�6t�1������ݼa����4�B��cg�O��g�|,.�^%����w�/�;h]�WepK.���9 �|�I�������}�Q�"�����)�(���JT���cAIi�@��(�ݷ/>U	R�P�Q���;��Fg�� ��a���:;ْ�E*�J���C7i��
z��F���	Ŋd���wv��Q6XU7Q�����2�:���Ҧ�D�Ţ(�T3y�O��9�
��R;��	��5i8���܇�aҐr��t2��9g��T�\���i��E�0n��k�y)ɊH<������%�����/Ā� b/�ѓ�E.krj�$kXc� j�U���I��PLH�-&��L4�|3�$���h�犨`���R�R#����;���㖓�i/�L	��T1U?�3�Q!=�;�OuD|%2W2!G�W��C��W]�5�����Lt.�*.\~=I����-%&5,�k.`���87��L�,@Ίi^[wr﫥�=�(��]-�x��םǱ��d娵}a���X]T-�z~�0��c��2�g�	6CBE��?iڟ�j�%����0�ǔҖ���1��:�l縢��[�3��ʺ����Qs�l.B�7�:����<�|�$��f� M�4���(%���!� ��w�Il�i�'�����)�
�t��.��,���w�o���}_@�^l��7�1fA����ũ9����1̲RZ��n�7[��������U1y�ܮ�L0���0ekK^��9<�&��D6�"�w�����;��S�Jk�_�4���"g4L�o���R6ۂ��ӾP���~|�G�������%�Fãx�L(iO�3s�JS������;�T-��a�5�z��=�s��r�C������[,5�/&�>�Y�[�$7�@���Y�8co<n~�x�(�g{������+w���-�27�9�J�<�,���hhl�{G�H\(��72Tj6�\���1!zp� �G+=2���|�aj�]��f D{��F�A���{������+�N*�0iW �}������2r!aq��;;��L�c��|fU����`��`���r-��Rݤc���y�L��t���]*+!���a����k���x;�	����7^�<%F�H{=�����\�W���%�c��y4�"nl~��;9?�����F���H���B+��B�w��HV	^v]��qo^T�����@'Y?Rj{K�fx=M;���ހ���{l���#j`�=o��ڔ�Ш�ye%�}3J	���wK�'�-��&��=����E���9-A
�_t0���7��I�l+�Ɉ6�0|.�@u����; ��[�6���'�
����c���q]����w��彸������5�輰�W�q)v��	���ě
N՚a�k��y$�F)ֹ�����h �uUp��!G|��u��6 ���mW�ǵj �}J��|E�R�\��<���M=�z�8���g�
��7���Qm�V�7�����~7Z��q��4v�\�^P�v�a-��"`�B�&��7/~��١�9;�U��W�/���k��P�٦\�h'��$��vo��sF�Ʉ�>��}8!t�z�j�82]C������f�����
u�0���\����@�Ov�ʯ�+��K�Y�e-�*GQ�7�}���W��'�X$�W9��5�^��[�u�����_1x�P��U����% �ϔwu�� Z3i�C�w�y-���?_0bk�����yi�o��%h�@G�#�g�����fJƈ(:�cT�'�0�pI,�mA���C��x�B������j��X/&��%ܥ�����i�i�R�N��Q^�|���r-�PK
��)q�'�>O��]���wj_�G0y��(�|����z����Ԑ���z�:Goy��7�3�a�=Dh��#Q_�d�#x��nn&*����+��K�8?���t�Ȏi��u��w=,(�J�g���FA��H_i�6��ν�l%��;��2X�t���:`���hE�̎Rj�G��}�(U����<�`��Qi_R1�#���i!�ؼ)�i���P6�Ȗfj�<ؤ���Q����`ap�߿ZT����P�-X��jnՌ�X��q�y^�^����8��/g�M�����T�6�� ��\fV²V��-1�I����Ā[L���9ˠQ������j$�#z�r��&J���<��l���):R�������}Amle��$/u�1mpǗ��@����s��^�NQKT*����_;u�����A�ԕ
f�<Hc'%�O�r������zŖ�Ğ�����ᬱ�*�M��$V�JP�<[��$I�ܮ���^�;�ρ� ?���_�	�W���]��� 5�c���mI�F�u���J_)�������i*kj�/��GoF�L�G�y����=&t0�ӱ�L�Cx&�>+�d)�kBU�X[� �y�۽AM�Wi��|�n,l��q�n )�y���#���x��Y�<��;5V�!_���Mx��j����zFg����	g�����3V�R�2$���W$i���kH�e�267F�dGҡ�	�M.����N�j�~��"&AK�F�H��r%*��O���P|�����AJ�g#w#B�8)�K��5:�opM Z�)�~�~N�+Z�l��OoL�Dl 	�Ak��*�����8�����"�!�]���
J����c���T��?��� ���ӡF�Ƃ��>}V�&P�]^+�&ڄ����!�?3�+b�\.p-��Qɦ��+�w��o�,8��i��K.=?}8�ַǸю8K���
�Ħ�PK� ���\����+��3��&��q��j�/H`A,l���d�z�=��c%ń�z�ɲ��3��X�W8^�	]o���@���