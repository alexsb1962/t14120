��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<��4#5��
I��q��7�y�J���K|.ׁ���	����f���|P��q6�c˷(+n�C2�&�=[惢��3zI�aΖ,,���� ���Zy�Y:�$^H�% �s1�=)E�9yj��7F��t.G���,=���؃Awޥ�j��u+5�Ln0��c�u=�=�d���
8b6?�� b}A��8��]W���V�a`�%�Wk�B�N}���{�������~�6�b��i25)��vq��zVg�"�!'tL��ࠃ��L�|)=Rꚲ�%�h���wʢ�_U��Z͵Mo���4� D]ޏ�C�î.� ���0����{��N���ĘEb_�@��6�lLw�2�R���,R���j\��G� h��aΐ9JD"隷�%ֽ�{���Zq���_�(fOPNУ��p���j-;�ePBM�]y����	��a�'��UZ����uN;}��<^K=����=Q�0��@N� ��s��±+|eO��Ŏ��P�p;��a*�{p[̹��������Ck����<�NaI{�:���*���.�XB}�l�t�p�B��Nm�U��*���|t/����b�H���8otD����� S1ʼw3P��r^n����`Û�]���W��:�(�I�(�$�t����>Q��ŉ\�X��$7r�[��Ms��r��A�1QĬew:F?�����n�W���޸�p���xx��qRHd�f~~q�	}��+W8fD�wG�U���S�&5[�L�(�;
�xkϏ1Aw>���@���Ӵ�)OFPz��"��גI=��ë�$�R�1��X9:��	��	�M+1�^oq��#�v݈��eW���情�96�'��4��)f܉"�y_�n���u�?�h��Ǩf���YP��RG%XO.Ϙ�WҢV,2l2f;j7S�	�=�9b̙)s����ᇃ1SzN�E�{�܃��_�	�%�}cC�CxdC��|���=XZ[dՍ��'�m�X\@S��l[7�#Ҡ�`���Y�_:e�6"�t��L_F����j�|B�.�}υ�Q�4�ȧp�ko�a�oQ�W Xf�[�N���a����W4@<ԃ���p<QJS����\W��#`�!��U�9��Q=�s>|�,��ݟB2�`�=��[��Gv��׋���8\r��^�kC �'�#ҹn���P4⏺�ꕷ;/t�NKz*h��}3�垓�fR��#'�$��Tp֮n�[�}��$����؛2!�N����>�1�4p#�-F�}��`at��1�� ɲt���IU�u�;KI�N'����IY��D�y����3o�D�wǩ�L��H3@�D�����%�@R�@���t� ���e�4L���@�a��AK��粅�1�.ev~��K5�1��*s>����L@B�.���K��N�ʈs�ڿ��N1���?�^�j��ukJ
���s{%sv㎮�ř#��1�c��)�_K&�6-�_�����v�坜ZI�˼��l���HY�Ud���Z�v����A_�h��6������Y#b)�t�H�$^BQ�=hd\Gh�ƍ�����M6Gq�_�C�<~�]n/W����4]�Y���9�AK�4{]��w�v]L��K?�����񄌱*�7���r@����<��n�e��bѮB �T��|�@�K��D���E-3֢l��
�V�g��*`��o7+�V�`L {16%�ɏ6�ňƦ_�qpYYD�"c �X��$��e+���XU�tg����r�X��S�PXD�<����-���� ϲ�r����O���}A��,"W������ww����|��`ZV��r���Z���8����Ⱥ]�b�#��H]�`�&�Y��X�S�i�9�J�!���P|��|�U�=��7ᾶ�P�6��5����|�ݷ�,���gŅD�$�_�q�-����u�Q�]{8^�˰���b���$-��R��n�.�c���b�QI�&��y{�"���#y�>�������
���^f.N�7����wy� w��hb�m�?��A[&��g���QhqqK�6���Zѩ�r�28���5�&�i�,i�z��/c}�j���ޑ����c��s�
��NQ��&���굙g#���<s%�f�#���Q|���k	���teoN��s�r�/��(�`֕2���(���=�ɍ6K�_M�E�����6ʡ8bg��^���s�sҼ!�8�Ĵ�Sn�e�%�B��>q�%#"������ie;�f��zJ-��7�Z�Ԕ���.G7H�#;��������z8�!��$������L�&k*�"BUNcg46US܀c@��:x��0��؁'�s����2�⚲8��$��7�u�ËO�j/�@��Z�ޔrH��&9pp�u� �_"kåuN��Մb44��h�C'HC��X�
���ChEح0�~��M o)Mԕ+zʯ@���K�w-��6�����3yO�	��+���6�a��V�{���/�ћΌ�s|�x����m�X{�����B.����Eb�<�sa~Ns�i���gJ!u��W�
n��{qg<\�K�D���"�ǭ������ �f�^�N���C��ݑ��DCVe�O����]m�pu��gJ���h�����T��B���0$}S�IT���z�
��-UȖ͓1/=s��J��e�$���95�pzӶ�p��(`�> Sp5����Rdw�n�fP���)��yFӓ�9�́���'��L2�Y3U�jh\�_ly&K��w?V�Kpv�	ϥ���q�R<�Il�{�SrV�KBA�-�����1�.�[ɂaU�������Pr���8��Q�Y.OFrS�ڊ�A�Q.�(XY��A��M�l�R���E+�,^�gU����	doz/zk�%��U-�'Vo�h{{�t|jU����j��`Wàl��5��UZ,? >F������5��N���Z��K24ȫ���{R6[B-~�566^��12VC8%�m<:g1U��Ҭ~0��Q�2��J�W���Zhi{"�Q��jCJIaķ;����,{qDNE+y��c�t�NF_���߱�>`u��И�6P��h�:�r�$O�%}֬���[_�����Mdne�]#/�O�ޏ}�$��^A����Pjzc��ǖ�������>~#c��W/]s�ؐ��v���5�2\���)����Mt�ig�)�Ul�����﫜��ٸ�-wU�P�p�_񯶄�C&���w*�`c�U <���}(w<�9�9O�Y"��o�iq�� *�1-�7�`ʥU0���5����^ p����[ѪK��jocڙs�I�������		�c#��ÌZ+�x�������x�'�O�WX�c�η��$�{���2@��|ޣH���9�j~���60s��wbʁ�s.ʇ̈́� �c��4�`'��ɠV��g}�)���6����0���å�9���z31�j���7;9�i qٹ�S��X�4�n����R1Ϋ���h�`��*|��!"�0��0���Fb~�#?��j��,�D\lAK��Y*X�c�ꗗ��S�Ӫ�]����e$��K�
���ӭ읣P����%9�t����|r��:���t����4)�a���_t�D��[f�֓��<N(�Y���s�yv3�r��"$!��.?Դ��0�3�����x	X��жo�Հ���h[5�A��bw|�U��A���
F�׃�r���ݹ��Ӻ���P�y�9U��.�(�������o]?^`��Φ���wי9��GF�V�u1.���FdB�c�6��fx-�xK�C�y2���i�<��{"��+��ݖ���z[���>�ǯ�T�?���������۞��D��b#'�qʍ�J�1*/�I.h�T*KB����b�m�c���Cu57!!=�pH�{(Ψ'vZ><-�o^�F��4g����DAk�P�d��<�+�A��?�.������pt�b$�*ڛ+�����z�e�%�)��/���%lq�A�-e�Gr$5��N�4
��-� EI�sT�4WV�A��-8���E&�qT�R���O����p���/�-�@7h��(h��%��LǸ+�GM�M�:v 8��(����S�v�����1�0�7��X�0L�~�.�t҆�ó/���_ e�K=��g:��.�M<�g�*���BG��]����դ7�E�;Lĝ�ן�P{nϏ5b��ۻ|(`\�P	�m��[�Z+;��ƮOӰC����r�z�u�g e0�)T�����X:l�����)��FDuЍ;��|�?[Dӷ���W�
�+�x[�`zۻB��H�x����c ��^z��!l^V�J�RԬC	���K��`���iw�X����}3��ei���}�������Z��A��l�b�����c8񪭅����:n���F��l���	[�nk�VO��G��<��a�Q��E���I=+�9%�i����Ѝ�|{�co���7�ki����G���M�;Щ,�Psv`;7���r�fQ��~{?�5M[��#s��R�u?<�� "K騀�6��� a4
��,�ՎyR3���� 7
@`��"�[�9B�S{�P��"�~��l������B?v��@z+��X)�*�H���=�F{��܁~R6�&�Fz���IT囥ΌD�F�8`�CT?J').�jzI��0���(«���r�U��g��̲G]��e�чt⏮�Z%�X��f�%�{m�ɝl ������U'�|�߾��ߙ��׊�"Y�+�Wa���AM��S���^˳֍'ܭ_�a`���Ӝ�p�ڤ,�e=J=����*��?7�z7�i�E#���C����;.�j�]�߄ٍ��~����.�e����ς���� a�(�>oFI)��m�G>Iٛ�#�,��W�ө��e���*��m�DS��U���8��
��0�*�Y�`�(=)'+T/0�8Zc 8�5j�9�8km��s�Yo��xg�.�^��E�5Q՛d��(��O>])�w5�t�N6e, �$�y��V���6J�ƾ ~>�������~Ӳ޶��&�*e}���B �i�Af$�LB�dyE�o�����`����ۭ3����[!]�8��Q�tt�2κ��*����.���m��D2`r��UY&�N�;"b�ա����Z~<y�5�a9:�<EȖZ��[�����3h����&�������RƓ��%�l�C��L�����N*2Z)���أn�z�5�f-.�[�k��A�H�y/���~���o�ʓ*��mEXQ8U��o��z�U[:�6n߆gH3w�������[	��Nͪnl{��<���KQ�Qs���}�;>;'��w�K��RZ%���r��k�	1�T�A�'������ ���+��~���{x�ʧ�A�����u�/!!����w����2��}1�x���NܷĎ��G�`Qy�GO�3��)$3|]U�,U��ΣU^���k!s	.Z*]miY�	�#<���Y�"%jP�w��e����Ū���Q�!Gʭ��,*�ن6f�br�~�Ϯ�F�L?��J�{������3�ׂ�OF����f�!SiqL �|Į�6\%ĝD~K�H�����!]���'���U![���#�S�`%,��ȉx��A����K|�'BS,�ae��t^��oD�2<H���R8��uQ#��V�K�8�������&���*i�q��UK@S�ƹG|_�!R��S�}?��WK�5�I��z�/�͘�n�*:"J�n���j���6d:خ���>���(
3ҹ����ϱ�s�����'+��b�q�P{�(�"|Vhx�Vɩ)p� y0����qR���x�v��XC#L��D������.xq'+3_;����I�!�P&�L��r@�	��/�sYt� �\��{\u�u�_��{귎X�\������F�@��}����	����j�o�p�i���!��㭪h������nj0D|�*;��$�n����vU숺;�2R�ek�K׀�$� v�vu)���{��xZuK��>���.1�k�!�2�aYEac�+�\������5����j?�3a�l��j��D(�:Ox�:��'�\�j���0���v��%볪�I9}P�`��\��T��	�l�7m�(O�7�����o���;t�w�d�\۷�m��4�����x��-ן8u�:k�ݡ��?��g����s��S�Ю�k*i�@��/�����Ti�E."�gqX6@����j�=����{�l���>���Ҩ:�O%S�}�B/��/���;��P՜��F!&�F�ֳ^Q��o���
��Q+`hR�y�:�Hvk0]�и�Qt���@�k^e���-}^2�t�������5������c�����f~z�鏟�b�^�Zk�5~S�L�Ӱ����ϻ�~jՙ'�<s�u7I&��^5��!Ie�c0�$�������d�m�5~�CW��iF����E��Q��eE�A3|���X��usjFmO�6m��	��!y��(�}32� 1�x^a{��)�A؞a]<Ԕb7%�Y,=�$6��%߹�g�5MA�����ÇP�
�p�WJ�ݻ�~��	,/ܬ��Ey���'k5~
n_5UP�����ڒ��W(?��2�}��U����*�������DyXu�W,@�NP77���\�Sv�޽����=��������c����һ%�^�e�e����5���<� f*��:�d�}�>�#��6ऄ�����$0�������V�-�� ͊]U	/)�,	��^��`%$���bQT�1������r�@=�p2�T8�I�%m���?�v�Qd���,�2g-%W���7�I��O܍���5���&p^3��p�	lL��wuR�S�G#�m�o:���;���Ǿ���iR*��)�G��K'��e��nU9̲ը%y6����� �!��e�/{`��dv��5&���
� ��S���<9ڼ,���m$�Fex�|�k[8K��}H��0w��$j*��Op�ˋ��0ی�<� ǅL��24*3�4��}Ag�	s[�ä�xl͍:���{���}d������υ�K���>?u�!�Lb�EѤ��b��6rm{���Ҳ��>=u[l�v5͏RR��2]d���:%3䃜�b�/͡A{��ɕ4ut���|zx�-�k����P�dߩ�ic�Y���w���c%�-t����1�(�5b	z~��iG[p����e��Q�W!{�e�\8?���L�p�KW� r���nܞ�
R�#A�ޭywJV ���go:�ε14�4�%I/XQ��d9��s6k�t�iI8M)}GN"�����S���Y��_o��O){�ҍ�r�i,>dۣ�@oz��,c�Ԥ���w�8�dp��"xN�
��԰��`��;��aHp�n:�2��A�T���ս�/��{UĊ+p~�^8�E1�l�t��]�>�'d.6���$W�� ѯPm�(��b��)<L�'� �@Z9UR�bZ&��2F\[�X�?ˤ�r%�#g�4�56� �����7�S�B?2g+���
z�Ttd��������*�c?M���	|�m W��R0[{�{%V]��Y�H�z�i�[pp�o-g��Z��9;�^Qd��.��?��]������Nᕸ[q�I)LH��G����|w��-,�P�y��!�?��
�[����?��o�T���-[K=ʳ���B"O�d��z��tJ����`z�1�d��[q�t�b��@jp^;-��4C�=��6S�W�M��{c��;��(XA��
��*Cmӭ�@�<!~+Q�U?h�A_�^؉���v�GMɵ��\��&��&�v�r"Ab`ZU�tZ/��_L�wwdθ���V�V�:��\}Yk(�:p(N>�Ȧ�*;����n#)���h���>U�/N�I�^��b��v��O�_��z]��v0��������$���G�B[�'>�j���Gc����9��s���	WM%w�Oj�ր���s��͒��:E��N��CJ%��|]�S��"E0��3�5��ôkz�YKt��n��1	\�F���d�����CC�i�і�9�e��^�br$��'g��d]H�n�<����Ye�$I��Ь�/���i�`d�˔��A�Cߋ��9�3}�j?j��y��SG.3L�z˰��� gk@{��m�삢��=U�(j�*q����(%�̭$qD=N�v`UQ��æz-qa���,�V�l��Q2Ct��[�g���g��Dk��4��~~u�1��uř�p@'������U��X�JMU�U�_�h��&.`�a~�g:8�w�`��[c^6����x�N��0��o���A,�9O��N�?�(�^�zm�\|P���������+��,q�ƀ0�S��[O�4�qY:���[=@HJ�It�u�@f.���˺��g��ܵçe�r���njx
,���[���V\���X�zS�����.�����x+ġ�|��I�Bԙ��$Z��M9�l�q^�sYd2ek*jڛs@D�c~FQq1Ż���*�Ih_Y�Y�A�$7�����O6�!�{��\�,��-yB3�(f�~M�ǩ/�9�7�VF�5�Q��\u��u,8���~�,X�	�o�|�yx(���P`9��ݺ�*Bp��N�\���[�C�g0�އ(/x+�0���	�-���m#Ī��U]���Bb�K3����]~����|L ch����$���iX0�c����5�&pj-i@G�<�fa����G�sR��=OK��2J����p��*v��������o��^Z�Ș*��[Pr:�jmb4����?8jA j"M�cy�&�9kF]�K�m}�P�s����=��9E����#�2���2���ߣ���>��P�m�=z�pK��=��0dp�k'O��Ȏth-w#r��������u��N���;Kp�s�'����m�2��,�`�at���%��p'ߴ�!h��S
\��Ч�MpO��S��:6�5����k���g[�S8�޴��ԘaFÞ�棝�E�v��=�ʓ�a�gbޅ��o�t���)5�(�_��x�2-BNx��R$8�m)�$z+��"+cUGʁ߭i�ҝ8i<MX=1m�`p ��3E��2��J�<�I�٤�\�js��-��iWK[븕����c2x�~�"�f�#���a�0Os�C%�1���z]rp��v9��<W�e-�U��a#��<W�6F].�O/���"���f���T>�k0�e=�� (s�B��5��{N�B�vuŚ�_�=I��i�v��H[7�խ���h$r���:1�Ͱ��=�XvARM�X��8�?[�.��q�=�Bg>n2k�HBUAPD��.���o1˯Kr�g����=�������=��ͬ�V��-jR�;�6���p�gp��O�����mF�xM١�^L$�[2K��X���~�X��!oȻ<Tciz�U|���ɽOԦ�3��F$VȺ L�.����D������X��6 _b���S&א(�I�������}9qoJ�haA@RC��a�����"�,Y]�pHBL�JV��90�!WuFȭQn�
��#rӉ�*�=?��zf�6t�h\* I�+��܁gasY�\mL2*]O$j�0k��F�W�u���ֲx"�Eܥ<B�47k����O�O��;��,.T�*3ha�nl@������%��+�q�>� ��7a�uyD���ˋ���|�a7��{�G˛V�:��^K4���¡�L����h��NZ��+l�g��61�b�t�bb�&��A��⡊��LJ�m�>8WZ�N}��D���mTI�#7w��9ok���un�QK䧜�:�ZS��V����Dg��M��$����'�1���&�b{h��k��J� ���u�o��MEiR�$�𭳑�/�P?A�u.���x=|��d�n���l~l0<����-)w�1\�r���ۑ��j�����z����Ki��0-W�^�Z�����4^A��F��Uq��N�w���p��M���m�K̈wY�U|�4	�KP2L�^�Q� fyky�����dȣ�O� ����x�Nb����5Wx`y_�q`O��vq0¥��#��j�"�ZQ�myVay���L���~���|M��B�]`'�\����XU�x?�մ`Ю$�J� �c��[\����c���i5�6���I�A�t�1��X�4�5Mp�O0FiM]��$��G�vU�D��_�m���!��5��ި�훟�n��M��X�O����YT���8Ȩ��A=Z��m�,|E�!��9�9ֱ�߾⾢H���`w�T���\��*>L��@A�*�b5��ܫ�xx����6p�_�ސ<�h�	^9������]b�1*=g���8�E�?�!���(d����A���x��)9M�Y�V!Đ[�$��j`�Z���#�=ՄGD6�
� ���<֌�b��� ���Kj-��;F}W�4���kW�l3j����"ؿ�!�����j0i��o젞�FyQSm���.�8��F���;����lc��-ZL��X��#�x9�d�@�:o��/'V_��q�Z���Yn�@������>���Xc�EH���T��9�կ�*�x���*^��4�s�P#J��x�]�u/�G� S��(�&����"�_J��h�����u���g���"*�s &"��a��Q�W,.%�z��v�m"���,kB�!�b�e��������?�k"��C"{�ܻR�Y��q����O*�m�N�hP%.���X����u�x�L��`oR��a��29=�Y����Iy����S$j��ҋ����'$����gv�)^��h!N*�!��o�:�:�oܘl��6:��*p�"�h���j��ҩݖ��G�Q���p�=4[��-u�eY�PP�n~!��ʧ��=2)r�(�������:�b`i�D��Ϳ��P.���k0+(��̣�w����b���S��3x��B@��'/Z���*�s!�B{λT/�xq*�9�!�$��Wq��>Q^T:"шY�R"����S	!U�$dv
OX��z�g�9X��k�Ķ�>��h@J��þB�W���Ns�m9{)KKis�e(�cK�障�[�OT���F�fd��Z�����'O����.%�d��f�O�o�4}��[;G&���yk��������H��;s�};Z?vjl�]9������\p�<��������J�2ZL$�eMl��.���i�{(!ZTڰ� Y�<H'xx�c�u�T��!�^��u7��&^��ֳ��α�4���r��<�������Y�k�;�g�����7=n�
=�Bw �����c��-�H3E;�q�����b/�/F������60d
5�����Z�b.�C=s���D�	�}&A{��8�{J�v�+j�r��Ğ�����Fe�d=c����kW�|�&�g<D:�4������)ϻDP��x˳���S6ڐCώ�B{W�ՠ��A�������� ��KZ�h�o�oa�c�h��ܷ�$&�x��	9����__�CH�,��*��(O_#ф-��8���_�K������Z:��Q:�jO:��WR�X�������g��rBM�[7�;i2�9:;:PXu	!:/8z��o�Έ��u�v�э&���k>���i��/9
������(�fޔ��6��:�澊�w�"W���)a_c����X���Й`])�=���Y�%�X�=��,a�o�G�ş�#�CͷB���!�߉~e{������`Ӥ��$I�+�g�״��u���k+'Ja�dd��+�&~ 6zP�?{������S$g$Ԏ����0?�:.��@��|�7��F�����s�c�dMn޸K���J����+X�ꂾGb7�(_viq��)Ƥ:�^G�����G��y�$Fb)n3it�2�.f�A^��3�K^���Ct_��מ1
��.��Ȝ���S}��:�2����Q�4�[ֶ;����Q!(�Om���d�/!�i�W���0R��O��Ժ���D,�;�IH��<#A�Y=�e�@���0F]z�b�)��_F�����z	�Y6��j��L�J��1
��Ԯdf7�>�3��m5����V��0%��=�K��� c-%��%|2[�0qR�H^hˬ���j��kd�tv�3 ��M�Y���ľ���~�J2��=3O�)�7��Q�S���M�C-�؄�&�ܶ�6��G{19 ��Z�˰�R��-Sa�$ ��T������/�E��	x��{�x��sxBd7���qcv���ܞ����9Ӯ������ق�J�s�8tf�8pSƄ���t�=��# �j�LeG�:��D��V��=�,�w�p���m��"H��U5��;�$���t�uxD����ܦ��1$�}MVK����+�ЭN��M`#i]��Y�Qg���h��n�n2+�����:�,��Gv�
�2w{O~�>���ɯ^܎�B�&��U����4,��JL�I�;|W?����N�n�o �vj�	����x�y�0�M޹�o���1���.�oxNj���������y���M#r^7��ؚG����b�#랝�8c8p�ъl]���&����[��ȍD�[:q�y0k�f����2-;� l&n���#�2�3� �?�߿�Q����]7G��7+�O_�y)�ß�2�_�:������eɦ�BJ���=�ťt��$�7�m݋��Z�a�M�̒ݰ+3է�=S�B�N������B�nA�{K��Pm�	���%�b���Z�F�sPِ��J�[klG�q��k���1�h
�I����["#ήu�|8|�S��|=�YBÎ�c����f�"u�8}C& ���P �;��!�!���zx�.T��f�~r���C��j1�K�0^��s��ȸs�K� ^�2�A��q��Α�F��N(��+'��A�堢؃rQ���T>��Ir����V��F,�I�r�2�s��"Nr�t���Ԫv���w��?�҆��(�v���Ql��%��_L�Q�X�ه�;	W�/V�V���ۖ\\��'Y��`�]-�aS{F�;�h��4�|��~q�'\����m�6�XS@zG�E�ꅢDv��n���4��#-�і��
����x{,���?^�i�^䩃>�F!�|^=@�/��$ؘͩ#�f��)�@R��v�!��bh#.d*�����t���t��L	�d t[G������7pH�qdUI)����M%B�!p�}	���_��4�;T�+9l�(q�6E��R�;W<~KbH���R��I$vp�-��##��\s=NB��NiLJ� i�+nic�&���X����M�n��#�N�l��Z�ږ�*��&��pʝ�$�,utii��W꾓���7��q��:�R���8/P͠υ�>-�و�&n�Q�=^�W������f����B\����p��J����b�iS��N�)B/_b�w_����F�[�q"�X��͝w<�{�i�8�+�,��,��wm� �y�����,gH�("�c���/�^�q2�%��>�]Y:U\��SY#�M�j��~�:��x�G��-e��lᦆ��%aA.\;�坅���9� K�{҂����vuN��r���#��=U����{���u�����1(��S�Mf�O��>��z�z�+;�V	ĩ6֞�u;"���h�N��%&�ncR��$������(ql���Ba
 �w��Ƶ�<9����GHK�j�I
��f2�n�%m���5L�&��Ѧ�IG=�ާ) ��\+Xo^��giK�{�S��˙2ѩ�	�k}����Od�]��ckkU�q���fp�5��C�g� 8�f�Ň9����|��Wʚ���o0'���`�e�w�S��Y���87J|�L�?$Y�͛�(�?]h2��ݱ����n�̽���5�V��6M�^��Ў�:n�}
@�a�"���sٍ�%m%��l�f�*��O�G�Á�g���~O�����6�F�KpboS-=K{S�"��3|?5�@6�|`3m�aG�i�N"E�J�9Jg4o�s�-*B0da ��7���DAa����r�$9�4�H��B��u�T"|���g� Q�@�����+G�Wb�$�K ^b��8�R����������N$Ɍy��s��g2˹���{��U;U�i�o�<Y��R8�Cd�&f��W�ږP6+i���a]m�(g쥎��h����	�%VWB�Ts��P8V�pZ��]w寐_������_��]/*z%m�N/:��8C��l�d���7��Ӂ��k!�D]G �95�!�졷7�R�|K*�:��Y�}M��F��u5	u�>��[v����9�e��Z�UX���5BGO������K��߉�E�C5N4���m��v���_�M�kȟ1��ܜMFE՛@W^-�O�n��p!����tf�߭����	z���EW��=�,
Hя@?�Ѽ?w+L�{��j;G߲�w��m��}k]�Ǩ��%���������j�n$P����+;�Jt�uA�\�n7�lLDG�Kd��B��I�it;��>�fUf�aG�NA�}�Q���	?� -W��Sſv�9�n���L��x��i���D��Ӫ�8ۣ���?�.O�w�C�:� SG����.Lܡ/��¯e�����d,5Q�x�0�5������ʞs�U��o�m��]9�\�B�V�֎��;��1$`����<�f������`��3䅝u ��H8�EF`���o�
r��-���o,yM;���7ߊe�Ņ#�.��Um���T(L�\���ꭓ>��m�n��)��@j�ն���<�&]��Q?��%r��ӍO����0��7d�>�ۊs�	dp �j�Z�
mx�5-u�m�d6��4_4U�f?�M��[x�4ETg�d\�1�r��]�b; �	�b��I��Z71�27�ˏ/��!���}�B!�=7���߀�rOZ9|����'�I����r���c{��{�),&w�8�;��P�|ﻔ�cl�l��-�5ss��4̍o��!�rP%r��"���a%�
NO� R| JZ���3h�x�TӦ�86�]d��6��K�g��-����zcg!'�ԔU{#�g��EU#a{��i'�%0V���z桝tIX���;S��UP��>.*=����f�ne7���c���Bᢻ� tyv0��nk�h��Nz�g+Đ�*9�h��`x���2qtR�&�H/��\,w�U����^���%�F�
Ԏ�BeIvKE�.-����z�A�:8�����y�����Y�_[)#p�rln*����Y|��b-�Z\�0�iP	/���%^u]+�*r�#>�įQ/(�'�ew�Ή64QR�ӵ�Ci�՛1��`/��Pʃ�UA'1�f��5��u|>H6̽��G8=�*�p�O�e�e4l�*B�%$Aj�z��+��l��f3�ɏ��}�_Txe|"�gǹ�)o���0�{�q��at�j�n��z�l`@�S;���j�@�Aԭ�N+2.����/.��"s݄!w�6�v��o>,���G�C�(��:]·��YV�Sd�%O8��x2��+(�M�lt�aNm��SD(ͥB��!�{CC���6�p�%a�,�?�dY�Y@��m_�h���ۗ�m]�9��'&IG&�cXr��~�̍B'��t�7�ЖƊ&x`����S ҺDR}�͘q�)i��:P;fY��ZkW����ܩ绻��nBil�A�TW�L30�B�L��Ip�
x9�x�4A����"�m: /�Qَ�g��	��e�Ε�^_��u�&�v�L���U9�� �@Y}���4��8�Q�w�@��og��@�g��.i5C�?��P>9ז�`�{���M�Ld?�,r��<|'+w��7w�a����w��:ߟX��x94n��^�ڟ�2�����X��ZOY|MG>Y�n�*,9:yӌ�֬���y��1�*���ǣzlP觤N�3��tC��4kK�c� G ϒt���]j:/9��]��&��ܝ�({J� ��d ��}�TR�<��>��U�[�z.rJC�ꘛ��mD]j?����#Dk��?-h�
�+t%
�&�>���ڞK��3�AO��h%�9Jl�Gb^��|򼧖v\�f�/t�O������㍱����ؠ��'���x�_G�]�|�f'6�"{�<��)���%Ȁ�f �2v]�Q��I#�QS'���۸#�W��z�ڡp��}��{�T���H�:��G¼5��u�l�"�zo�6�E�v����=��a��}.�F���6 ��>�'�?����8PՇ���V��S��һ_��8fЄc�����4G3D�,���~����3��auhV貪��G�2��e���>U�|���Q6���^�n�6Uʰ��A��(x��U�%�p�������u��3���~��3�UrC�\�	0�حSH$���jX"U�������!]��T�J|��ϢV%��Y+%�P�xA
cB�$݂��ڞ4�"��s���H���6��.ݿ���)r*���_՛&�	�u$�J�U� &�~�}�R�����ɝ����nK\v@��
W�����"_9<�K(���oz뀑o�������I����DOx�ocamS�.�����tZK@�x��x�HJ��z2S#z��"�iU��'�Z�Y�ӢR�_e������� �Ȩ��H�`3�^;�S��~��XVntrMs���]�Y(i��Jնm�@�a<;EjyPv��8(֊��
AN:Ⱥ͜ە�ս�|�#%ǅ�?4d͐������*��\,]�^�I8]���A�e�����1�'(�yGШ l��}���M������NW��].�<_��ܳ��F�{��}���#~�����ܒ)���S(�Q�)J�u�ܳWL�H_���c~��!���b-�Ln<���@i8�X]�w@�<���e|)�_:�RF���e�js�% �+��:��"*�e�K7�G��lgǅ៴e��b�c����R�����PQ����*���藱S�*t�jm}�INۛ:>J��]�1F~�ԉ������<�!�9$M�c�)�ի��B
sX'Ę�z�q�YP�R'����?�kI�s�b��('l��WlaezzL\�U�Ps��f�Nx���a�6��_����S���Q׫;}��!t�HS9�o��|%�}��џ��r@7�@r�B�R�X�C��c�	��,���L�[�Z_T��Y`Թ�i��8�%���6K�ͬϚ��+�XNn�����N.Tt�kfP��)1O��{e�;iI�����-=�_(�����L<��TZ��Y�rq#<���&���+%ϖ��[T�;ݶ�i�2�It��_OX�<�^��	���������x;Q�yC�{�m��m!�D���<�鴍�e�3u�n�q��bm��J�(��(|�i��R)������ōGS��f,�/�RY�F��")@tCxq�`	���J3��]i9���� k������`�b~Z�t�]-�2�^|8�VY�2�c;����G��l�l��ϰ�;���;��ݫ|I��:�-�8 �����AS�0&Τ�(��=�ӡ��wd���@D_����/}��J׼(yN�r��;#b����?@�H���E����X�����\��
+4�<���xnD��o8���~jы��k���,b��:������!'7�\��C0��56�(�k.�:.&2�j��o��icj
S��?��h-s�����E�������f��K��8 x{����ͅ�dU�Yt.�eXBS�&X�=�]���AX��~/��
���B͸��vq�gr���
�rߘ�e`�)$�g�U����og{7�r�d�Df�=L��W͗f�gEC�y�0����A�*�=�v����I���^.z�v.�ї�)��&����mib���:�!#��G+Q��p�D���s�������Np%�K����i�<��IO���V7�[��#�M��3�����?V*�&a�����"��.A��bQ��v��FR\�8^2�e	��+׸�3`eW�Z��`SO�yL�z�9M�<��g���T���!F�Z�s_����b*B�\�#�<M:� J��C��CGvǲ����}�k3�����Bp��W�'��mǗX��2y�`��|g��I����Ӳ����c
6jD�����!���^r��Ŀ���1Zs�'����j�W&'��;�<�W����=s��L��:c�x�Ni�=�j^g�	4�q�9Ύ�r4� �K�a*�mx/A/���@˨�@-�z L<��˅W�c�(��rԙ&٬&L�Ssw�uߠ�����=�Q���Ѣ��Dq�Ȥ�# ���<� ˊ���M�/���~B΅��*��eN	���F���s�����S*���b	���.H�)M:�)ו��#��:�fMHfר���<��^���jG��7�]ْ0�!�6��J�)/��'8��A����QrbQ�JŐ,�<+��?ꎈC�ў�l�0����a�d���s��Z�j�=� Ϝx|Q��=�#���$UP#6*Lh|���KP�����q�����Ot��c'����쑺���%�X]\0�����$L9���"]���3�r��#��	8T^n�d=KKn|�7Ʈ��������3�eJ����9�vW������N��G�4�V��/orJ]�G"+]�.j܂��Vx�mG�dhha�<D~v4����v�Ee�G� ��1u֫��ܥb����u�u�غ��kD���M@ϖ�M��-�$h}u�lo9�����pÝ�o�#i'�Fu@\/T�f��@�Bl'n88��w�i��Ӊ��M��U�g�pi�a��^Q+��
) �#J��U�����gw<	eu8P�5x���9������M !��s�u���������%L�����S���T��_&��m#nw�Z&�
���������u�f�����f��DcU�,��bvĚ����j]Q�>�W�\�Y.�ڒ�D셛Ù􂯩�d?MķL��V9���R�����9\:?9��Js;��K:4�N�� K��W�Ε��^�:i�,!��r��Ptt�t��/�h��~u�`�!)�� �����E��:wD�)�9�y�J�煽���Ǎ���Q돸�\�f,��$�(�����G>��Ԫ�EU5�f�`��O}���q��w"EuJ�G�aI{��70��!�gcC.��.�����:���a�|�wB�e���S4Jy`)��^eY!�Z�զbȯ�����v67�,t�s~;���膯�$����;9#��I���[A�s$���!�.8�ޭj����S�k���B��:S�++�Gfe��d;BTU�x�9de���X����JOz�#^%q��;������[$R^��Wǂ���R���`	� ����~z���������W�r7?�" ��{f#h�@J�7��|�Ք��'ǳu�/`�k�Hq�%|)c�~f��v��]q0Kn�Lk �d��3��,n��:x���j��>�N]�\1��~��8�h���qQ����[۱�)�]�Q��0�Tl�'=�,�dx��a^2�P8�G��b��oa�WP��j5���3���ن�i�8�#�>_$8(Y
��YylU���:�J,��FD�b�h$���$�QN�aP`���cP��h�}a"�q�nÁfz7�J�llS�Äw�T�z��թ7(��lT�Mc�
��m�.��2��8���\��Jqۃ1����ĵ̪W�y8
Ϗ�L�d_�􉫕�LJl�Pƻ�R�0`QD���a���wOSC��-�G�a� ���,I[yRֵe�����ڌ�:����9;�n��m ��**���J4������	ߐ�K�E֐�Vr�%Po��sA��K���M(�c#Z=�"m�+\��?�E	�u���N��,γ��)�9���$�Ά���g �WZ�?g��XHc���z�4�8��RL�Z�;��E����gykSz����|篛�d�0�|�a�K���hku:��g�)Y�bW/�|u�B����ܮ�MsV���*1��)���
�a���t��]E�7d���q��p�pŀl�L�͒Uű���̌�?E<�K��h6U�
u�J�	.ż2RQG{������7̀#��=ઞr(�}�����S�� d)��4�zPW�P߂��z�g(�U6�W�3L¹��R�KSa�t���r�rf
�<�i�T��KqY���:�۬�%��^�XÀ�:U(D��dxxa��8� u��eew��ɽ6��ЈOӈ�q����y�xp�HO��
��P�)y��1�����̾Q�=�#�{^b��拊�[�.�֐$��O��<<͵h�И��=��K	�O��,@�&�<��� p�Uz��׭�����Ǎ�#�>�}�/�s�i���+�m"n��H<k���s�
Vt6J_hp�?� ����YL&] M;�ځS�[�p��m���l�aFm��.}���~R�Z���v�a��3O��8�aT-4dn�)DYE�(i���qs� �'
��WG$�əꙋw�$=��~6�M��c�.��Ћbe��YI��0����#��-[4Y��+�fvn\�v;�}��y������
~��)��NԪ�4��{�	B�V�[�������%GO��1 ��Dxk���ev7�pk�#qДrםbg���X�0(�j��y��
(���/��@�U��=̲���7�6���2Q��y�j���C�����Y���a&�uU���*�Q��W�h�2ť����9n&��efV�>��ۊ��Ց��(�{�6���ݼ� 9�+��v�
��X��J��^�����{��#�V���u@AG�W�,����i�v�ܵ�e��:h�;�~V+�M�L��\�̀��}I�<��N
��=�2��{�S8����\��J�1���<OK����lUp<�2�������R;�fl��y%��j��ZP����$�⊤�
���}-�{Å;/�c�לɛ,�
9m@���+n��k�S�H
�_��}@����F�f��1B�{��xn�L�����5�o��&@Mʅ
+�o�ޖ4�����}.��^_�Ǜא�#�D�U�D5�	�I��"�	�ն�3:����H�Z��(ֺN����6	���:6�IT�B�3�>���������wm���UuU�Iƹ�Q��;�fz��{�NG�1P���JC�e��kX�Q�AF�����IZ��_�C����r�|(�s�h��CT��ł�CM�O��^��;a}�N��\��\Sӈ�����W�=��]��#3v[��I*M���`8��.�m�$�£�N뭹�r�*����
@�'�&��]����u6Ur�EO,�S伌����լ;�Q��wB�F
�:od����	륓˙f�Aq��c�ɉF�9�Ω�Hǉ)�y}�h)9��������
���2z^{��`��$Z
G���U�� |<��=d�s]�`5���asF��-}1�e�O3T���ߕ��h�W��cJE�4����ao|����/j彷�H��yx��X�4�%�qGv��9����o���ֆ�[h��j0�^���!�ń��J�L]�ٖ|���&�jf@���`���.-w�g7��։������I���l�8��Ռ>O1Ȣ�Z��FߕT臞t�ن[2o"�����/��tb\W���##`�RWk���������� [�řp��e�M�Md������3�(Gm�˃a�[�>m� ����s�
o���Vt���F�l-�e%�'N}��A�%�� ���R5�2J��zTZg���80�A�9|4]����-b��)D�鮉��\����*�D�g�iO- ��_�1��e�D�шa�]5�૫fBMb�>E-a�ӌE��Yt�>��1��?��|cE�C���>���_�����w�T����2�N D)�7�'uLJVB�[�hҳ�p���1���RƑ �7�b��YI�	=��,ھ2%.�yh�M�m��R�+��w�Ң%�w̴�fkY�4h��.�Τ��6��cǒ�X��0W�E�d�.��2F��/�`�_��苓� z�R�t���v)����Q�k��k*�M۳���mKf'�>Ң���:�K1�DͭJ�#�W���n�4�I:��۾���J'�8��T��+"6�Wح�w��"��Bl_L�vSGh���'P�%�Fb�����`���{��z(�b�A�;Yy�����Q��P�6���/A�Բŗl����AYܛ)\b.��~�{�Nφ*��sI:x%[ZV�"^���W�M���6���,'�1L���)N��q)�mS��/9���7�`��6�-�x�<�4d]��@��m(�F>&s�.6ŏ��57�� �xO�5�����+�-�{�=��a�;YC	�
~d�4Cq�� L����n�^��&�=�qL��7���NU���Y�yIY0D�˼2
b�R�
���{�8i*s$�d��/eĩ[E�j�Xt��Y�3�����7=w�M%��p�t8��x���{�9��uX!L���~$�#b�'�4�jɤ��^91f1��g�_�V�H���./���-��e(Q�FCc�J#�/��4�v4��X�M����t ���\	C:�T.�	���.GI+���>5-�c9Ȥ�"�3��NQ�:�2��tq����2�ÿ�ġC��1{�sc�ub�貭�N�H"Q{�F�+� _,��Nf��%�h�,e-ITV����w�EMj㕑��ʨ r�{G���C�u|���G��퉘��I3*�����t�c�?���n��"��n�s���I��Z���M��^Ņ�e~��&Ȝ>Cm��>L��0�,5�_U�<� e���k{3��EcsHIBB]'�j�30,�9�`�ς�L�i/���f�{��:wXR#Ks���w��>c�wsZP��*V�Y�i����O����s$j�Q��v% .��aA�B����|�ŕ�«�Ѩms>.���
�-ԧ�ώ�!;���5�O��bA�R��鈶-}?p��%�2K=9O�b�x�����e/��sV}ap�˲[^��X�pm����+����n(:R-=�=_�\����7.�m�X�.C	�.巰6̼��H�ȗ��H�?{��;���t*#dmUr�b_�$�x��+�wET�TMfS� gs"�eЛ\�y�#Þ����z�7&��{6�MA��.y�j�0����&��L�}�(ɲL
@k�{M�j�+�?�a^�m!��_i���o�BCh�,WzRۅ<F4�	<^� ti�P���	q�����M�g� F�������a��FC2pP���*��ӂ����)��A��>�!�%�{�! �k{��L[�Tr/Դ��n��R5t.�v�$��|)鿮%dFt�6M�BϕIq���L�z8 � ��ͶՊǎD�
���B_��IG���3��K��'�v���W�w)Y��/��G����^��y+��u��~`��4\��O��"�؞�9ր	O��f��σ�~��0r,7W����b{��N��2:u�=�W��� m	��a�_�b^�j��g/�6���嗳x^{�Ɏ�S	�`���dUH����L�e�}�>�x�D�%��rƕ2�����Q5v���䦭wV��r�}�
%�V���ls��Ymǰ$�̥�]��t�J][�ۻ���l��[5sR���[��h��U͔�����ױ�h1�%��Đݜ+(�	 raD�խ��A��S�6�I���'�r��G����G_�o��D{�a��)� �?���
�	�* ��6�d9�m�}#%����`G1J��3���=��ZU熴M]�!r�-��H����a؀<"���%t«��l�"~�aB{�p-պ5%���l�����J�s����b7	�#H��#�]:�SV����v/Y�j�⚢�H!��W���!��o�:R�d|��z�`���7Oѷ�c�}��Lko���PĮHMS���xb��$�[c �ә����-�B�*j
�$RSB*��O+*%wr����kƼB��eПR����SWsFi���^w:��i�M�#F�c�����ymY�WJ�Z:��c�Q�~<	ԑ�n�4����I[ 1�,�>Ž���:Cה�rGg��Z��@��֓���〢õ��ӣ��7bICo5E�#/�&�+j@� �f����>�a�{ޙ�6BUƸ����vy~�o�y���KY$^�	RoG%�_�o^\���{�z)�D,x���f�l
�ޱ6*ۗ�d§ɚ�h�2�`2K������s�<��ʉ7edRci#� ��G����goQ('V5�u|�2[�W(��T�R큨4���}�N���O��,� \+) !y����o�^{�@5Ph���+��/�zw��>��5E�\������������`&D��rkx�� �7J���w�xaQ��+BN �8�ei|�:�8�O=�[���ό�o��\��^p������t��A��x�
��칓������ޗ$��6~[�?9z����%�&n����Yu�_�P��P��̄������l�nI �M�\L#s5�һ��}P�)�4y�w�v1R�"�Ht)S44FΕ}t�~�]�<�~r��R�8	θ[�V��ڿ����1��q��Cu���P�@.�����a�1���T���4�9TKkZ���h6�K-pr�ϛo0�|�g�*Ìr�7 ���v=��R,uZ�)E2�mj�������N\"Q��
����"l�U3Y͇5�}�V�nEY�`�-0q�I-�1��/Ë�sL�pt�o쒂.aG��y`]NV����=+��ftqX�>�/г�9�3֝�>�h~���N�A�a�.����ձow�)��)2�Z4��25M��#�us5�o�LW�vٮI̢4~r��ӏBx �i\��'� ��?���ɔ��������
�3�b��vڪl��vmQ���0/o^tk涅o\j�t�g&�*�x��Ȯ���Z�{?J��
�*��нZ��3�S�ͣi�8x�D8C���F6\��cRO2�����5�#v�*w�V6�����'Bb}����{������d&��T_����8�$���h��]�����)�^��{�0X8�xA�H6
��굽Ml��r,H�nq]ߒ8\%�Q�ITB� u�Я��t.}wB^�t��C�U��*��ԁ�I�m�ne� 	(?��	3��i�ͺ!b0M�9�(캝�Ή��+����"r2L� 0^k��֮�bB*jsa��h�2V9V�V�&�iA-�{�if�m9�`��[̎{�i6�O��$�|ϼ��<��o��
�SZ�5�xx�$GU1�����ݏ�=��Q������S��~vƢ���KNO�x�-N�]<���L���:!���
�o+�ȡ*^�?��9����4!D/�K�gCc��ӯ�3簔��꯵|P!��/ә�Σ��˅��?��J7�<�s��S�+�b�[�zv�;�!�S��E0�U�����W���p�F�hɢ��U����Q<����}�ӭ�8|F6Zt�I��G��T\���VrZ+l�G|MP��O��<�܈�Z55�Ԇr��QF�4�����Υ���v�>�wF;���7�_jb3P�:�sg�E����3�nzS�'��`S���1P����Z��˺5g�'\ ���B�U�0�l��j��ń�E��L��O��/���i���/4k��4VU�d|��l�*�y��2z�Pwp����B��B�	D��$E5%�~_X9��@+].���@�I��Z����8g�����׀6��k�t^�S��Q9�܉`��Qq�[v�f� ��k�6K�8�G5��#�=�m�E� Ȍ��bR""N6"Γ�� �P9�W��I�~��H�bƞ{Y����+�q��� �[b�?ͱ��7��4��4�[Մ�M$�Nr�_���}�c�k�dR��"��& ��s�l�4x+��iE�x}a~Wl��Q�#N#�aV����țfp����e�V*� ��E��Bv�����!�GY6n� ���Y򂠛y���!������Z����c��d`G��Yf�!F�g���RG⑲���0�#�"�Z�f" '�=w�$��c>U��������Q>��YXrg���2��U;�9_{%� ����_�d �R�0��`�
�p��{p/��͎�]c#�Ё�����J>���x%�žE�jf2s���谱���2
�\����@M�<>�W�a�'�2�C��"��V&�YF[;N��'�][I��WcH��o��x9H�����a5�n�P��Av��D����6�a�u��q)����WEÑ[�˹o���HP�,��v���ک�	SfQ�A_C��`����n�i[��;��KlNs� ec�3���8r߰-�ʊ�4}�Pq]M�8B�t�Q�a�O&�d