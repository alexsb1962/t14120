��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~їZ�8M[p�S3 \n�Nc�p/�cǗ��p�c����U�
���	&�:i�^]���v�bB�G}�\#�S!�HM�x�y���r��uL������5��\�����[�CƋF�nX�KHs�0�<51>�9N�I���U��|-�C�TCT����V���f�16�p^*C���6¿����CbG�^��o�zwU���+�r�2�G%:M��\yN�g=��������Aj�1��Dj�KS	�͗M)I��|P���&�g5/ok)'F����" r�BҾs{r��Dt�%�����Dv@?�v)�*v�B�z���w�4ko"����]�X.�l�~�����0����m=I���T9X���ؙ:���t������F|������L��xZ�xr��og��y| �
dHnͩ�#�إ��$.��7퓄��H���\������q�Um�~����f�A�7]1w�Չ���\�;�٠� �1_m�C��4x5�������|_�U�B�8�������c5׼z��:Es�5^�o�>�6x�pK�lt?2����[g8���������>�J�� �
�eQ<�ZP���\���m�@mM[�r�&"�_bƝN�/�6fS;n\v0j�`��ݛ `$�7����
��y[�+b���WȊ�ʰD�3��t���H[���64t6��x�Aכڠm�"�`9�X#Hl��`�"3�xp�JJeS�J���iU}O�����f��6�p�q���aċ�D�v,m�d�����КI���&s
K����r�9	@v������*���:@\NqqN�4¸���7���&�W�sC+��%���'w���K����{2��LR��'�=��nF��%$ވ�Z��u��Ҡ��g��(3��
GK~ͅ�Y��Q��!��Ǳ�C]êDr�|O�K��U��G��_� �c���!��Y�<�s$�w,�Ug��X�w�;�]n���5����F$h(���E�㻨�L�:�2���s*�>�u�W�5X�m4RCzǣPU2 @S��2��
��$��D_\iRȟV�����H4�qQy��R�j�)�@�7�w}@��(�J���8�%��u?���8���3o�L���������]/����zsG�����NJ	�a��0ڪͭ�����a�%����͐6Wl�\4ɮ�f��O��ax� xP�J�y�����>�89 ���ܩ^�l!'����_=#�F&�G��`��U)�{�_��yn���N68ݟlo��`0ǮG�%���V畷���' �{��7�B����̞�������Qy�-��5��P�\h,4��w�-�4+��xO�œg	�/��i8��-���Ջ�ڒ�u�뙁Fu	5��ؔI�Xͻ�CR��$�Jkf����ؗ�p#o�D<{��Ű�1�_m�4�o�j:�U��E9��ΎH��n�M�=[��X'1~d�-�~�Q,S{��碣êX�]B7T�MglX�\� Yk)5W�=,G�3��6GP���%�)�M=�V̭��h�3.-�*t��A��~��;���WFs�f��`Z�:���Nq^����7��t��QZ�I��=��$�ys����j�gd��H#h��+�>:h ���s 	�}�m��|�\ǣM��oA襸�^iV)숭���4�b�� {�:~>8�)���ĎG;;�؋=��8��J��a�'��]kҺ4��-NyL�%�VقD@���ܥ���%��'NH��B���ܪ&��b��N�xiN:4�y��g\�?z~{ED��V�a� #f�̊�s3L(Sʲ9�Q��XZ[�^,�f���������h��L�15�#�ű%�"m��lzf����J|���2bZj(�Q�ድ�%�=\�Nm�d�B�F(���ʞuG^��u4%$��o���]chǣ����Hn����]�3ϻ���+˒��;�m$Д�BxU!�u��쒨�MaI�~�%�\SG����uxu�H6�Ȉ�~N���i�f�z�-���j[W�~��͊^C0{i����+\\S��kFi�~��_�l���ѧ&Eu�#q9��?C���=a�����pA��Rmٌ���rF�`�믌�lʌ-��8�P5i�Tl���y�mMܫ�����}m��W0���00�f�X����g����0�0�]��J��m�אpWrm�*�f���XB�1�	S�l�o�.=5x71u@�&�AP|\�|R�Җf|L��/�46�[��%(j��H��� ��ГD����,�U�f�[�nxM�Ł��:�U!3��\��;��(�|IqYV��#������1�Hh��'�3�2�<?,�[���P?>:�g�r-@w�0ߤ1-9.og�="̈Ć٥�~/����B�S�S��Ӓ�ǹb�h�2	/z\�Gi{��!v�<Oq�z��^���s�o�U�����=Rr�0t�zr��L��.o�81�k�� ��P��\q	�	��lP���*����q^�'�~��{�d����&�|A��I��[d1{��4G����9�p�5�Q��T��AF4-}B�9���j&_�< uT�A�o��^(���ےģ@��(�
V��q�h`��P��y��ML�'��}�w�k|;���l��[���\���>�醁����w�����P�X���BO��BA����R���gol���{T�U��� �R�Dɼ\�^ ]��M�SQP�Ѽ!��9M��� �q�U{�K�:��_C(�7�,���~K��?�����0�r��%�&Ҭ�Hĩ���8����b�B�>߇�(��0��A�)�KB=��e5�W���.H]A�&�W4Qt�X����#�Dl���=$�����S߫�cO�vX$n�kn��,���k�hs��iT���X�	ĮW���˻t:8�%Zt�]�/L���6���"5��[��.ļZ��Z�vf�JxՇ\������y�\��^s�+r�nZ��~�Җ��g��+G��{�4�_��"@AϢ�ƣg3�;�$���ը�ߗ֙t�}%���O��'r��3�"�`�|�PɈD�?���&��fI�����@��k//Y��h	��7�y|So��kfU���^�������^1s�h����}��#p��G�󄀍�&�.c�������%d�)��K�8�M~�jy����q&�p)�|��3����Ần��ê�k��#Dբs%T5t�z[$5��@��L��(��+Y����F ����=�洛�&����وdP�C$wv�M��<��c>��0;�K�k3�,0k��B����O�T=��0�4�k@�Op� �kYź�T�Y��Y+�����+{�߉Ȭ4��x�̬v�?�&�I�&������هR���A�T��,����p�P�N%�+��yE�@s)���m��Kb���c԰nӸ�1b��F�R��3e޽�W54��R�<*���
<�ȅ�Y���/K% �_�Ɓ�A�G#\֨,|4���)��3FG�Q|fB��	�d��o��z�z�Wǭ�s7��-��!���*��.n�JO����az��_�ݘ����X�4G��-`�iR�jY�!<��±[�����^x����9_%�%����=z�:�/ԠS��O�$3wI jlM�፵���Z�n�[�4�Uu*$Z#Ѷ�EҘTcXJ�p�g�����Ǿ��W����o�D"^C"�Y&��C�_��L�/X�׺Y� 3#?��Kн����ڞ$��m|�L�*F1�ɀ~m����5����C�gԸ�윒��ׁ��/���B�0Z0�J�w�[l6�ďǰO�,�0G��c3'��1��mL5�a*U4?3�]��R!�[�}9�tD�*iEEPݻ��Թ��u�UQ(b�1��E�b�����JD��k!���ª� ��Z#~a�̴w�|��p�b蔮%{}/��������pJ�4��"�$ǨC�w[���镩NE%��'<<����-�R���?)8��)c����0&#JwF��e���׿$�K�zQ��t�1L���/�+�>,{�<^�����u&��d�����u�� ���YZ��h$[���3�p��v�++�rF "�n�^����L� ���|8;�>��{�'�C���\@�qQ�5[��q�yc��c\Qh����_d����������6�P
߹��|M�k��Rol�+� �E{�ԙ�)7����\,FA=��@��4�v'_)Q<�t�q��)V��<�m\�zI)��*�.�f΀l��ɛ��7Ҿ|��&��T}?�^�(L���r6�!��,6|ز�4���q��Z�\��0��\3�=���R}߶�t��U���ΐ�{l:��R�+� �!>�[��%������OB���[���r��@ӻ�Ⴌ�OZ��	da�j7yB@1dE�����������!4^�S�CL!^�>�n�T��<�׆_c�o��om���4"�q����ߟ<���飈�cj�Z->�o��D����<0�7�ة~ӥ��N>�O�ͷ�N-<�LI�4N��,buY����aT2N�(X���t۳����l�9�d7���"�m�H�7��B�-_���-mvq����{��>j	z�YN��e!��r��f��aMV�Я���t����B7ILk+N�p���7��`�l�P���Ê�]_� A'yT��Jg�GI��y��s6����n�_����vn������og��K4�{Q�v�$��S�<X�a��%PG�5IH-f�?~��ߕ]�Zy�)šo�~���]K2���Ѻ�x	��pz���ʉ	>JĘ�x"vV���S�G9J��Wb����L�%~7���f▃s'EA�3�m�#�*�Q;�rtb�-��8��<�mn� ��aq�%{x������a�1���K[{0?���B���.:ظ�5�֏J�D(<�I2�R7h�Ld�Rl��w�T����т�H���}�h�>�La�{!PsB	���9��WN�p��%!��' �g1���N(�����&vnd�,{G�y�7S�����/�M�	uHKf���N�D��T�ǝ'��?~Y���n���BO�'��7_ҋ�\A�&1�fߺ�Gږ��`#���"U��>��48U��;��ج�8;8�s<W;Z�����87}Q�x�=����_%4�?%��*��x�2L���0��S�j��Ϯ�ed��ßyO���Y9~P��3��6��&����q{��U:�t:C����=����y�d`�� w����l,,���+#CG.��C�Ώ�kT����릌�^�t� �TUCP���"��	Okyع��IG������@"�N{�K�Z�E�?�o�7�lҼ�t�_	=��� i׿&�5o���գ�?��t�qqg%�ŧ�E�ȍ��T����|^A2�Z[%�	�~��m4"�j�؁&��d�W5u���yY�F��k�>��vЍ�!jp�ՐE��V�F`���J(�C��̦��Eڑ��,[MJ\ ���]���ҒG6��e\("��~<b�[/T��\�k|"dJ�;#I�����+�����ԠoE��x�X�9�����$�����l,�Ë��� �FR���'r���'9�#SL����٦Gʞ��I�n`�) ����ex��{���j����"��'䄷MӴD���Nm�of��z���+E'~�$׊��ֶLT��t�u\�s7�r�O�j!6��)��3y}Q����P�vP*|��:���\_popg���W~�A�@�L`�I�m#R�%�a�]KXd *��oc�<��O0�-�K�2V�x�4�j,s:ǖ����f|�Ӎg]'V��f����zs��,�G�_�1=��BZ��5��ݏ��㊆=u��c1�րV�k-��}�?��&Dt.C� A!��!��b�bn��8��Q B��y�����c����"ڝ='v��ex�!<W,Q���itfJ�Ehoy�s&U"�E����g�)u��\�eUy+�ޡm{ z�e�+��"|�c[v���_���T�6N������ֽTB/B��{I�E���v�U�֌�@6�iͣ0�J0�T�[��e��h����Z�T��� m+�u�`��P����^�Zv���z�������9j
N�{
���B�~����%���-�ػ����[AQ�9��2�u��@A�ZbMx�$��H�g,g��0�>��mv�.ު,S�k:ˌ	��C����4>��CQ7-/�( �k+�&�^���l��/^	�׎�KD�]ʌ�4K���@�;��9�\� ��I�(�~ďS�V���x�R�EF;J`��*�?՝���S6ؗ��ck�:W^�м�!��V�]D�c��ӛ�`�ѬO6�-)�>P�K}J2ɥas��MNt�Y�ذA��6ڇ�z��tE"�Zn��zb���М�
i5��@�I�XxA�B��G��o 7{81��$�o� H`�{24����dݏ�K��{��	����G�3��W�W�n���㴇� =n0�!Sm{�b���Ԟ��Zp���n�C�����7�ܜ�̭)yd�+a�	x�-�U����B������3�ɒT[m���#9>����OB��?������U"��KT�Q�R�˾�`�e��c�n�h(In'6�zEyO�	���_~�C�5]�|΃~`O�8�A���`?���~[��9t$*��ލF��%>e�:y*��IP2���Oqt��r�4d�FM��n�`���`.gud������P����Y�=��bHْ�L�\VImf8ZU�@�۸٨�N�JH~h�~��x7H�>�>Af��"D��?�i�B�]j:ƳxJ��0���nJ��{4t*X����{F��鮸r��U�>$ȱ��	�S�3S��K��8-ƷB8�X=����X���㬘]Ru���\�F���	n�+�Q�ye���:i��!�Qٱ9wG@���q[� �!�5�(��
ﺓӳJ� ؙ����������<X:a4xz�<��i�`~;��EG�BIZ/.~���k�j��#r��v1��:��Q5Р=?���G�e���"�������3�M|�|097*o9���-�ZHʙH�||ί"�e�u�!��ŞO"˔u�	CD��G&��|�t��?�<Վm_����Kݬ��۵��Qv��������i��g�òdRA��	d�Gx�[K���������t�;�!U��ׇDt���i37�����㛎�@�źl�r�S)�+�$�V��8ET
K�/�-�X���+�¯����K�=�,eA��t6�G�����}�%b��S�NX|@8E�J
A���q�������;�VA��>�?w�`�%�0����R��Y��������L�.8i�Z��l�&�rQ��*ձ�|"^u%��5W�{���f�W�^�O�aO� nxV�A�1\���E���5Et��}oR�{!�\��nl�Dts�x��:.�H�B.�I��L��^�0'�4g�����Y�J�a�8�d�D��QQx2^hf�e!��`�p;��$kz���B�e��Z�Iyc1T�w��9d�8S'ሯz�
��E���as��3�=v^��i(|u\1sB-BHӮ�?���I�����\5~�RB��Y�7�X���m���\5L�:Y�KV��Q����}`���+t���їy-�����<�Z�g&K��/���2�"]1�
��޶�/�uȘ}�̺ky�g��to��[��'�k f*�S�������{�l���)�׻C��'�V�e5mq�zO�xv�Ă�[����A�g����9Zf8����b����z	:�Y|��(*>v~N�W�^G_�;ұY����_�j�v�"_�g@�z�od)��	�7��@�[������>e�>����'������F�jg���#ͨޣ��7)�����?>q�n�f`�=����?�jD�%ϝ��2aE�"}�x�9��R��y���<l|z��%e
���I��ES
j@:I���H��-����Y�j"i���n���'���| ܬ�B��H��B���-'�x32�֚pZa)���P%jM�9�x���r�R7}��3r�Qa��<�6����
���4�u��z�8��ƹ�Ȼ�h���0����^]�P\ D�4� ��BfNv'�'&RĨ��=�u�a�ٚ%����ՑR�}�)��\��+*�`�"#q����ն� .z��_�Le��?�G;��Q'c�N-��S��"3]C���3�#��YM8����3��.�o �wK=����� �>��c��n�k�c���t%��OL�6��)M�~����d��~3��+����[�C?3���)�T#��"s?��e��|���g��e�N�.Z�	'}o�,�C�6�Xf�6�	C���%
8E�%��oe��C^(�\`��U ��v�x�I:V&v� �����"S�>��P4|��s=�F���"/(P�AI���/p{��{�������-K%.w���'�H�������uKH�0��a�bƬ�CЫj�jؠy��h�S`�8���H`C&�q���g���ș���sՀ)�(����h���{<.M�W�݌��0m�~.�Oo����3Q�0C9�R,D�5��4��S8���o�E|EG�<[�|��k�2�M�nq�6o�k_7�<��6��l�J��<���r�Ɠ���F�gm�%�;[d��V	���壿]��f���j��=�"e�Y�ي�	�S�X��FQ��RˆI�yq�&��:Z �;ǙH�rp�;����7�
\X��������V:�cs����vpT�C��R]]t0`�)0I\E,�8�&��Q����g�B�k�u�s���[�m_-6 -�����瑫���R�]�`��]#���3�~�Z�(񻨕r���n�M��|�#�+\$����� �)(�?�v�3GK���BZ�y�lj�����/�����8�<���|O9���#���`'��`*�Å&9O�?5tg���^�H�-]Q78�at���d0}� ͷ)������,���xU~q��9�9�V�S�"3n�D��wBwe�Tо���386�K�<�a(K.z1���v ��W���w_�7��F~
$�~�� �����9Ee�����m�����Xz1�sMw���T��Ũ���%���E���n�"|y]��	���$���8��R��E�[ �+6�L{zQ��Je��S�rsDc��R�J���u�M�0��{�2�O�L��h�/C��q��F�t.���P�*�����)R� �;ʔr8�Y(J.���.��@I�RԒE#4����d3����{�S�����yfW˗�i9�ob�Pz�+���tm��R����M3 �2��Oܻh��S�Ίep�\�1瓋cn]F�:ý�4�ߵ]�֦�:$��`��K��J.��gF�>~�h)�&���&�U�
�Ut�Vb]Wñ3�ئ�iyѷLz+8���t�?>lIDJ�0y�8����%���7�ʙKV]4�����MXW���e[-�`�1bZ�c8E�� �rlv#��(�*�0�E��t��L���g)h����}����|��шZG�b�j^DzˑpQ��$!�c&�QB"#��b�b�#�>�_��%w \_d�u� C��ܿ���_x�8��]���
��ɘ�}i����&P�' 	aH
r��n)<�$��$[mѯᕬP���z�◉��t��] �G�4>K K-�l&�i�dɹD��D�*� �P�t���¥�A5��<�0ɷ�h�<���;��5�5'��u/G*C��?���QL`����E��p'�z��Fa�!X�f�������00B$����l���~�#�Z��D ����J��m
#kT�HK$�OM���������:�U��c�K{��K�>��m�|_{ծL�(����J�yZ��(�^z9Yb2�.�+�-Ҳ�dn��q!ý?�X�&�硧);l�~�x=��[A��Dida���7筪z���m�/����i)��!N|�ГV��)�j���p'1>^c�������6)�.Zd9�k8��
���uጴ_-$���������t<��dB;��"y`e�����v�o�n��4��'8o�/_(|��[���������ms������dr����N���:c��ޘ������?��ʥ�ƚ;W������*�s ������@��@�%�+�x������터�/S���h��a3��8g8�fM�9#4�y��'�x���]e`�S�+5�M�pL�	����(H��L�B��e9�\�`��i���}���X)��eՒ���4?5Ki�;,�8��;�F�_���S�N-`<���qaԓ��_�N9߽�*γ��������� �p!ؤ��Uh���K~��?�?��7���,T:f�E �E��oZ�Y^�7���L�I����K�ˮ+�$灙ݐ<Kt�f����"������r)~�񫧲ݱf5��4�n"�Ƈ:'���Dd�����ӷ 7�T�XB���#x��5i<��J-�.H )O|J.�"���^��)i����^͠��b��8q���B:��x�(�!�":'��xd��BU��e�P������ ��y���ٜpj�X�i�h���^1r�v0=�Iȸ�ܫ�������GnΜ2�Kn7�ܾw�,�e�
M(-��N�w���1@z�*������+LǋW]aW�c4M!W6�d)�/������I.0�/�zX���}V�ǧP]j��(LT؏`�?�?�A_���8�rrhe�R<~�^:�"��XR�P	�U�(��Բ���l�.�l{ad��F����qa��;�.ĉ�����A�<��|���(��ݚK|4�s
���0u����P�ՂsĜ#(7�mzf��w��
k�܇3oS�|�C�-F����\����Xv�?�A�^�Y���x����\�8/.)���8�G�&mU>bw�s"���;|-<jʃ�) xD��B�wl*�Z̴�Q
s�LǞ�5��^T��'��IЂ��γ˓�T"��Aݑa����l��)��z���pnC�eS��ǚ�B�E�1#�*5B�6�u�E=������6�dO���O��� n;fU��ې�߭�d�y�VO��\����q�˙�	e�'�"�|˴�.BU����� J6�i�$%l3�޷��A)�m�����x���ktҞ@(�^�&��_P~)�$w�3��V��ф5�������Y@�C���*�]�T@��~���(n�
���tai�be)����7|4ځS��%Q�c�}�Z���i�0<���ۨ����r�����	Z�>���6�R�} ��n��]d&�|���U��Q��)�a����L�5)�	�zE�^��ڭ|fR_�JB� ��N'0�J���N����m}܁�'˦�c�-Xa��N>�Eԧ��o�f�85�m�E��_�ޞ�H��׉�ȧ���V;Իڹ��K// b���Z}/_�D~��I� �R�� ��&!�T��9�!���dn׸� 论q�!%��[�^:Ͱh��+i}C�������a��X��%�8K��Hm���e���5^��*D�wA�J�^ޱ:-ܵ|͐��;Y��-\��|c�6j��X���E�`�R|:��B6�"U"���߅J>7�,�ɧLI�5l�!�V�>u!U��hG���d��	˖��V����"�Z��Դ�6(��L+b�����~m��C������rJ���p��Zu�C�&̔e�s^���2�Cơe##��X��2�����O#Jz�G�B�b�}��� ���?w,�	=�x�/�H�U^��ŭ�)�npՄ�C���Ib�߁����!ZC,�ڗG��E�eWw	���������9�;i�(��E���yIU��_�l���?*�C�:!�'�$]�Yh���5���c��S�O�	��`��Zmђ"���G|��qB��|,�8+�W��}9UH]���D�T��_�����>��i��D~�\z*>^��.�< �����z��QZ�m��p�}�CǢ�%�|�W�<y����|z�ګO���<�����z[��zڽd��El6�AϢ�I��eQ�m��X�>v3@g&��hק�.f�HG#L���#�m��k'�ED���-о�X��\v(�A9c�5P�����@�Z�j4Q�^�Z���&۔$��.i|&=��vl�2��w����n`^xlY�������~V���*h�[}u����a�݇��N��� &J�
�1mĄ3P�e�#	#�K�c�&���$^y�f�E׏�2~���Y�N�-7����傱���V=�`�݂W��,3"�L��e��F	|�_�M�O�T�|���UɹM�L}g��k���)sG6�'w(-���џ1�![S���7�~w!��#WP�?7�Wf�����%fq��ҴWN�L�x�=~����t��%���DU��]��܈����9��[1|�ٍ�Ugp�;�h�gU.����2�5T�����	y���*�i�S�Gg�jy{�E��oO�&[}$%���&�Ί���a��n~���W�O�(��!��.ńq�$)|A�Bz���@�3��|u^i2�j�w��LC;�:P�d���Q���H���$��	����_ˎ����O���:�тS���EZ��ͣ�5���Ӡ2�>��W�j�1�K�X�Cڦp�2'#���ˌ�y6p���S�8Z[W��VƆ��yƕ��-*�@����s��5��o=R���]���{�ϒ(��#�E��A��K�ey<�N�U�Q�w���1��M��6k\%��5]LN����@@AJ�wA���h�3I��<XYU��S��q2����6{�^�ȸ� ��L�9�tm�7�q(�WE�y42�G�>�
'AFߢ��_[�ۗ1��6���^T�2���ٻ+�)�caL���J0�'-$z+�#��j&c�f:��qykR1~��ˁ,�*�٫���NV��@�+�a4
n�{�4��I�U�~�C��3�#22W:lg��6,�*s�l>�F��������cֱ�x����:(�$tW�=?���)B�h�6���^�@��=IE�j~-H��MBz(X����tr�GƵĺ���^3r�;^��*�ke{�S����?��t$����M%�y��8�dQ��3F�LM{����Y�ܛ������bA��p����1�j�?���C�m;Po��/A�Y5�}a�D��,�Z/�\�d�"�t��z]�����8�>�Xb
�F~�#�	3�Xq�u6��7��3�����l_����9L�{iiQ���0�^���}�:;^�d�|(�
������BD �ܫ�)���a��:��C,�{rb��MY�e�u�T�[*�(/�*��B$������?�ϥ�܁��P�ރvzʽ�������k��U�U�mRD��$�$�D�@����y9̟�u�� � ?nJ/<�m����U��<B��a�~��Wc���~�OO""��Ļ�@��r+u:*�|�5�*�,���G�Ө�,��|v���&a.��듺jK��\-��<�4�;���-��5i��p�ru-d��^[�"+�_�Bn�VC����? ��0�M���_��ӑZx��9��xB�2���Ppr���H��U���@'yJ7�����,҇7M�V�wGI��P��lu�mu��p�?!<�kn|aF��_�5�,Wx��T�\FP�|x/8�������*X�&��Ȇ������d�~W,v*���هŖ�T%�����SG��s~=l(����\�v�69����7p5�Q��Q��B�ل�����<G9u33�3fOk��{9{<�F{�'=6��Fcy��F�����������~^�k[��1�
�s,(I{EY[��/#聝ɢދ�.w�]�۴�P���K=�����d g&�ƛ&l�ء�~��J#f2u�"�" �/��O���"����ȼ%/�=�~�n�'�iݳylq����8'��5�3-�lr����m��xmy�;D+09G�V7��{a^�[�~[Z9I_n�
��4�-	�N�ѿ�(ټ^I&��� ��Â�d��$�3Q*<;�:@�&�|���G����_ӻJ-����C]����T=���mq�#*����Y���2�����;�؄Kn��4�P�r�e;�ft6���,8B��}l�����ׅ&�ފ�؋a'�`E���T�#��.��n��0$T؂f���x��8���OCL�����X�����`�i4ʄ��'{z�����A�ݵ�/�x��qx|Ź��f�A G��CS�LJ���NZ`'m9��%C�����_�'����4�3�~"}Ψ�E/@q�/����;�S�4�=�(��jŻtR@KPL/,�0���'ǿ���
�["t=4G�$&OzW=�d�x�r� MF6(�E�Y���@���V`?o���d� ��]��at����ΐжm���H������Z��ز�嘤lh��Y>8��F��帠#�w�z����2����H�(k@�쒽~��/x����_b��2�9����/귴���<�3��Z���q��2���Q����א�^$��{<��Wl�9c(�x�= ,{�ĕ�
��b("τ��4��=,''�KiX<z��|����rDű�� � k��Si�rZy�����*+ь����I"_r{�*xB=�ߣ���9`��+�%q��p�	�3�\
��Dѽ.'Yo(����ᕤv��1sc�ёhQ�Ff:F+�Y�C�X���/bT�L�7�t�U�M��T�0RR|���'>���h)����k)��7'`�@=�-�7�-+iIq��s�)�Zr��D;�C����	��z_�f���/��݂i��\Ϙ�m´���n�u�<쳖�V��T�Mg%F�2��l�q����Τ9V�� �^U��>$�{}V�)���kx�������f@�f���>f�7�ͬ뇶�����)v�'\�����H](k&�����Z�]pWI~#���H�to��a�W^����C@m��v��P�ީÄ�i����P�!��6?����7��j��D�:@�C�m����v-M�C �i5
�ٶ���M�@r�4����R�ٱ�G>-�H�CP�"'m����I��d��C~èn�*6%�'��=O�o����4��{`����f4��s\����
�0˂�, .��i�o�v۽��,�� �Nvm�O/\�4P8̂��C��r�m�
����a���6I��W#��͂8Cbq����9I=�:�2��|���|n��i>�r��|��˵����S|�O.:MYl�T4�|��V�5p��Y���0�T�Ue�"�<�;+}�܉z2�)���)TjJloF`�j�U��Zc]��f�o�'wL�U�A_����4I��ͨY�7�����R�� �B�Zo�ʑ<U�hY8&&\�}���bN���m��Ctվ:�h�s�����p����"��@���8�I����Y�X���{'f89X
r�Ύ�y�i�������E�%UFE8Z�z��0(vH(��Tx���xu�u��⡰�j�;���Z�Ds�Kw
�a�f�b�za��4���؋���6��#A��1ӭo���z�����f���m_��	5`B��8ʠဈ`���r���3	CE��[la0��0R��\������?%�p��0Ua䶨=�����g�s��N�t�<�����s�ʭA��l�w��#���w,c��j!�|2>x�"}�.���￢I�:8n#�8�/�;bd�a�i��!�̰���u
Fv���ɨQ\QZ)�\�*�Β�k�;�����s�x����lӦ8�q����gG�=8���iCD��0Ӱc[F�7���*e��b��!מg�����l���.���.8�A�N���A;"���O^ӍL�9J��R�>�,�\������v{c)��%�t�������&�#ƉG.j�[t� �U8lS*�Z˲g��ŧεwq�EF�"�nhKf�4�=:�}����������1�l��/���l*a��kVn�
����/���6e�c��PYۺ�#싎O,���~sn3*�=��;�Ț&��䡤�[�����7���p
s7	�K�/�y;�?RI	�<�#B�������Y�!������n��n�.7ՏYy������Q��a�jk�T=���q
�S����0����^��_$�j^��~Suۜ�$��%�������kp�E���{D�t��|A���p�l厈MI�Q`!ғ"�T
v|� ���$�@N��Ia?qv>I<��qz<��{��Kc���':	F��\�?��GnW5m�%=D�����F��u}�0p�&O�I�����g@�,
��=X!g�j59SH@�#\������g,G��	&'�(e�Uc�	�ꌐ�J_�2i�Ij~� їD!�t2���
��;R���y���FK<�G`V��W"7G�|��q�;a߯�O�'+�J�u�3㜏R\���5������5�U�������_����a�!�����-*M
veG�O�����᪠��&����q:��a�e2 ��T��{	\�/}An�ta��V���r���9�F��G���#���C&V�8���6lT6�ߊ�Kf�`Qk�C6}5г�sR��źLRTk���3�X�&�%�.���hk�@�ґ�'��J�]C���5+��4C3�m�3�=��d�����Н<����Bfļ���}����Xm��������.]����f�Dt�����VG7s�ѷ)�$��D�U�� �S�U�pO�
�L�һU�Eb�4�õ��߄[���yy�d�����J$��^�\`�J���a'�\(5ِ�@�G����^�B d�F����˪�og#*����_�i=��ɸ���)��<��URGs��o�K���<$��O�~���}����������s�!�����0�`f�&:�I�?x�	ۯCk��pl�ސ��I@��|W�u�y��7����?��f(��w/3�U��+k�-djael�L�8s��E�����W��2���T7�H��?��.��1����BF,[�Kc�Iz���y�xy.Tc����y
PM�n��aA@��OX�&��{��[�����QY.���\�X����HפT���ה��F?���ա��L%~A&iD;�T����	�{@��I��;*փ�JŪB%S�#�?��y��LK/��]��Ԉ� W���ܴw���gN�~�x�Č<;Y�r������r�F�����O���������!��YP�qր�v>��G�|�EÇ�H�<����K���!VSVK\����TT�w���|c���e�� 6ӱ�m���^���ΨqE���2�͓P�PR9�&n�W's�6�Ë*������VaFي�,����@�"H=�q���<h�e��)-��x�b̻��R;F &7#�ur%'�Tx�W�������Ǿ疏���Ж�����<�q��Uo�Z�Lk��Q��'@E4�����8칾5|ޕ ���#��{����>�a�Ҷ��S��P�=�x��\���D����cل����� k��P2���̤��ݸD��&�r��uV�1�����a�칌�r*7���%�`���%]�/��f;#���u�
��Bմ�o�A�L鎱�[z)����iU����Wc�q���+V�Gs]]�RC����*H�N���u�G���u������bA1�>��ͬ�0�-Y�xy:�>�B�
�Pݰ�vX�vW�`�P[�At(QP�=�ib�|����kF���� ���FoTUEo�<!�\�[��Цg�5z�}	%!��Ս���Z����Յ�����B3����<A�,�TFe{��z{4�Ɍ�6<��>�� _�J��A%����H�.6_1�o��C{��W5���Hx|3�\d�:�Z��s|��;�ڦdQ�D�.&j����k����*�m$x����v������ք��[K�b޿aW|ֲ�i^l){t�T�iMH�f�󏄦�-)���P֬�
��F�d�Io_�)�ed�ǿ~棛�c|O�\H����F=W9MU.0m�/b�쨅i��T���9�0����d����^�!��I.�)��M��K'��F�������h���s� %�s����9����H��[�͇$ O<�H�p�V��-���؜����d ���K�w!r�)-�?�IKθ4�D�ڿJ�d9���u[����|�w��4����M��d������� !pʙ+VR憚Fos�y\�.����
��
�dj9���7� 
�G{��In�q)�%���V|gۂ�]�f��ĩ�t��q�n?C�A�&k�j{+�dV��)-01hD�Jg.���P�I��?�d����wMV�I����+�����
Q�79rb�|�6����qd5�<5<��x�c-9�8�<��ϟ�POߠo6jF�0V��h���z�����3�y�k?����@ҷ'��,�TM���n�`?Ѽ�/��G��W��+�3��-%j�ꈼX�#��
���U��F��
W�(�*�g��Og�Z�۠�q�_��C�8"��4R���o,Q�D��C��DP��ҼkO������b@�
钹Vh)���x�G�5=/Lt��Df��#j\ڰ�ZS�7=�1.aJB]~�❺z�1�aH&g��^+�{w*�q!�9P������f�> Ic���V+����{�6��9<�X�m�O,y�Ym/]C�L��8aT�HCɱW-M;�\_��K��Q[.�E/��Gp��A�P�Ch6�В��rc|���b�
����h����9f��2-�BE� M�O�,P�;�@�` �)ª��i�,�,� �9jrp �<������i�� V}��՚���O�Q�<?+��A����f(��z�W��dbM��^@i���t�=�H�S �x� ���� 8y�d[z�>��g���1�(�����	Y||������f%oʟY)P��z%q�����q1���l��~]���bsԤ�ӽ��R�CJ)�m�sy&�碄w�&� ��Ǯ;9<՞9�Z͇}A�ԟ���xerK�a�����))��3Z�ǏT�;�d����IF^g�,�,��� ��.����H�����+��3Ql��}R���(0vC*�ß�tl��j�݆9I�P0���jkȰ��S_!�(�����L��P�jcl�=�j
��~8l?���倨*i�����ж1�F�-Æ�,j����3�"�zVOHs�Rקnt^�8_���TuF�m�; �-/W���M�a�oo��N��u.dc;�U>�� �I�Y���=�'���g���Qn��[�ڕ��!�*�?��7��?t�����%e�U'7T(�*6�B��Cpx�m�	��~n�f�][�M�D�����B��vƮpq�J!��{�LCrW\,���28��.�S��i�LC��!�wKpz`��1O��-��������R��R sE$Xa��#M'8ԯ	Ko%x���3JM��_;�gހ�K�n��Cp�LdZ-Ҽ��#�Jq���=��|��		z?e���U!ON0'Ƕ����
�Sv��2#	]�
m��iU�g<���U�a���V��n:B��A�%��tA���1�_�t�{��գ�a��T�n�@�\;������b3���$[�N����6[%=e��L��aFZo��=� �|�?����+�o�o��~k�b����I�!lb��kNGd�|}1$���p�#���iئ�n���[�[�a[<��Ϻ1����@�q��q���U�Z�6���$�d���.������G�n]3�Q8+��f��N��d�=|I����p|�F��E���s����T���&"��!��--�Wpj��B�!2�1�	qE[U��{D-.�K�2���.���d=m�sg>]hk��8E������a �[T1FG_�/T#���2wM�D�i�b�P�	�y�������)��OJ�r��+��m�9��g�/"K.�v%Tm�"!��Jtq�}�@����'�4Mڔ�g���i:(ܧ�"ls��_�����)��E��6AL�a����{����x��88Pp�8��h��O�=�R��X�w����4�'���j�Q�����cN=V�E�Q&�79�ʛIH�����	���MǤ����j���}�(���M-���Vm`a��O�6S�'�~�>��@-��|�X�~a�1�1p|���W����Jd�@��焳���()�Kv7���;��P����XI�&yU�CUU��_�O�;]��6���U�d%xk��*e��q"��,�L�A���[��{��5ο�8u���f f���2��@����Sd�p�q�͞l�pb]��[�t6X)G[����z��1��ƶ5�Ǥ�n\j�k���g�f]�!Ǝn�CzRks4$N4"}q�@�F����m�Г�
=i=0�����3$L�g�i�����:j�ܬ��d����Ps�����u�Yꈽ���iK�����?]�F�{���&Z�_YDb8g���lN�����Z�,�(P<�v������jd�����$CHн�=�$�Pv@�T�;�?�3�s�)�0���A�Z�G�SP<Ǚ��5,'�����/����\`���2g���/f��3�V�g��o�>0���� '�QЀ���?Ӡ���r��.��Y8�h�%g��Q7�n{@��E���Ϛ�Y�}� �ތ���q��SuWbj�#���6����O����0?D�"��m�ס��'PƮbdx������(+X���w��kK��.����.Bh�7�N�c��<��2W��p�ٷw�`�)��:��`������ ��HLonRO�戈��hIÍ�ܠY[3tC�#Af���S���(���9\C0��A�n���)(B;�J��o�%��&f�O�]Kz%ƢK����sXd�3�E��[����R����/��#����BH[��Qز���Q�B�Ad� a_�����6T�l��S�c����I�2����: 7�aJ���	�BZ3�~�(L2n�R�����R�q/W�XďA��4�w�*�h_c�cΧ�����O^�C��%а����W�=h��"�~}J�ή�2DM�^�pU�Gc�AQO�k���v\��z���eң��� A&Ҷ�|//��1j?�>1zُ/����hG��Ks�p.ҧ�]%���_}�6��#��z��{�B�#K�(�U��J`���`9���a�(�c4o�\��GUL����Տ\r>4Õ����E��G�2�b�\�b��fT�f���ϑPn$�hjP�Y현�@�kks^z*D,x��Kq�Y[Ո�f����l*+>n����u)���YW,q!���~�W�p_��ڈ/�$=C�ml�<.��؍��nE�%<���l"�Ph��m�aD��񺓮ė`f	X�,j�:cޅgB���1mp^�x�DF��">�BvA�I���~ȿW[ϲm���a���y���h�J��3��3�49mS���b�9H�JdO�VM�!R�C��fҸk�{�	]8�G��ȓK���Q	��z���c��E�G7���Pa��m�i���E�1[8N�杢Q�1�/VQj4�0��$��݊�W�\�|��;��1X^4ͫr���>A��;m��9%+�ّ�j�*w�q(�j��'5JG��U蚊y+*Ϣ���q9���"�Q1��F� ��[�T�tG�Ya����!��)f�~��[�|ħb�T<�KK����( ��.k�tq���I���¼��&<2뽳���"lǻ�&�@dɽ�^D�YU�Z\Ĭ��*I7��,��[!�D�$V�O���m�8e�)��Һ���gC9��I�V��Ӎ��a}{���,�I"�����6:i�;@�{�釈	(ǣG��-) ݀�i�tw��b�{y^�Y���fs,��;'P�ϱ�=�_�Χ��9�8MȒ����g8�*d� ����N���u��?����ޚ���������>����\�FU��pl����d��:�X�Z}����WU���v����'�S�F����n�?��<���Wl����q��)'B���m-�x��{J�v�8�(��]v����Lݙ{v4z�1V�E�T�8��Q��=:Ip��q׾Ș�������{��ͷ?��Z�좠Y#�
{i��9�~�Q�<��n��g,�9��[-���*�)�=K��u�x-7�����@K�-��v8_B3�A�!Zx��}͘�EK�dF1E���v*�΢Z5؅��Cf�Lh/��ޙ��`�'3_f��ns�H�0b�sΛ���1����d�����+h���X�K�����M��4�z�&�?�����k4$k��^1a���R�EYG�$�-��8����$+eM��<�U����Ȫ���i����w��u�z�<��D�j�Q:h�C��X�r���Tm���N!>���]ć/�X
֜���\�G��l@|�̖���� B2�����h��&40��5"VZ��>ai�I�ʩ� �����%`��-�(\��}lJr�!x��-��1x}3�A�`9�"<�0�i��u�
��m�d�7��~�2r�;\ς�i��R���7��'���F�>W����9���Ţ�n�&G��1_�R�z����3C��g�p��w� �t����yd��@������hɆ��w�q��!1�b6G���e���fS�1k6�}�$��N�A�d�F�vϸkIw�T��,�����'�L�"M��6񑱉i��
Җ�f�����h1*[�h8�{v��/
ߥ�z�5=Ч��#W"�f0�S�����woE��/s��@�/M�-���
��A�DHK���F
�5@& �_H�t���@-��=
�^'<9���{+��oE��[%4�4��J<�L/����D?6P�)Dk8F��/t��r�<�S�p�aknN&XKg%���ܢ}8'�:9��r@⁷G�P\A��Ǭ>3��bNܛ^E��k���y볷���f���К�2��`N��x6H�j�ep���� �Ԉp��n���'��Yֈ#�.�k�ͦ=�O�)t ~��`�M�ȓ�=���Z#���]+�Ų�JZ��!4�� =����t��;�n�m���Ly�=�ęYx��|3��xH&i��b��u�U��_�)R��L��(!�;k�)	����|nU̳�S�]@�7��h��Q��
��5��RB��XC M�?�=�qϪ�~���(��+3�@��5.a|��V��?��/-�4�OC]�L����ˬ�÷�<N4d ,�W���Qmda_�cy^�A�N}2B`���C�ꃢ
�B�����s�4~6����>2Go���I���7]�����B�̋�d��W)Rе3������Nzoɺ��׺����f.��_+���������2F~r�˕u_�v�S�&Q�
2����R��4_�;ۙ�Y�T��`��=�:�ܷ;�YԊ12�6���~_��o �{��[50d��K������꿔��Z�wJ��m@~ |��;(b�W�9�II}Fs~]�y.�Xq#|�m�_n���Q�����9�S&�/E�I�T�����@�+���7�۬���&:!��s�[��a쪴��7��k,S߽����g����C֟��,5I{6K@�8c���N���;�ok~�����&���4�X�U�I�53M �ͩ	ݺs�E�������b`p����<L�ܱC�<�[���ҥ��tA,�<y]��SM�Ҫb��ZaqF�fH�%jT���_F%��%t�o�J���6|EuWf������!3�rK�3����𦼬��؊�ï1*�q�P�6�32���Cm���|�F�+���"�+�u�.1�V�d-#8����k�@�a�Q�-i�y��z�^I�->h�A���s�t0��~�i�L�8��R<v�L-�����Rc��g���������
����mMG�̻��� 3�[ˢ�w'� Ļ6�6�7D߸<s�@�N�.�9u�[w2�k��B�����`�m�j�}^O�� ��"�U��3(����t�cF5ɀcӶ?�b�[PqX!k)-�.u߽%I��}�J�Z!"�9�����!:�~
p�"�mWt�al�v�M�ı�_sr^)�Hq���ũ�";��~(9_�q�������
ͧ�0����W����w��a�|As>zu�l�2�X�*�X`�0b���_v�K���Wl���l�@t3��"(Qquf��w~�-�������e��N�&�'�Q��]b9����.u^6��V�S��\\>+g-�J�l������� |B��E�ײU�N+;�iZ�2T�Ęb��t��V����*�M�	f�+�έS��\xJds�aesT����H��,��N�ا���M�* ���������*����z+�������h�3[	@�h�ש��M,g�
�:${���' R�a]ӻ�c����#���b⇃��.��,?؅��A�l
�k�/�<������yn�=��D�·��Z��3��c�t�L2���E�}��AJ��TO�Ν~d	�3%�[���I�V`kC�d-
�QYm�r�A*���-��?��������N$�G?���uC�3��wc��GR�cu� G���N�������hqH%��<e���(׍YE�=f�O�J_��޿?���E�o�c ؁0�UZ�$d_�>��4\��r�˔���k�c;4az.w/i��{n�q�2zK�2�Y}	���A�y�<����@�?�/kI�n'5/J;ysX�y��y�7HZ��3��7�h�NK����J�'	���8��٤O�4����������ؑU^)�t���:��w���Em�tN
ɶ|�5\�lcn�$�5�]�C�S4Ҧ��wk�>�\5�ĿyZ�X�"bU{���UU�h 0�+�mES��C���ӡ�g�xN�`|l���I7-��ŋ
���a�M\l��eݖ'�.�Z�(by��u]R����%�ͥ���]��+�����K���d���)��qZ��a��@
�\��Ln��w�H���1��w(Y0����J{��V�uqf�T�Pa�l7�=����g��KS��p�:E��x�T+-ZE�?H]��h�:�&������ЄN|�d�=���	�Ix�1B�!�3P~�u�}���omX�o�8W�o�G9��n��Z��t	]����v�YM]sؠ��켳�%��y���4��g�^c�u�ۡ�aY
�m|�"bH�<�l��P]3*>�`im1�7�m���D=���)3�x-~k|ؿ5�N�(1V�˝*��5�&Gq@��5�`V�,�NÇ�� �p��yGn���ѿ\R��(l�ف�� \7|ُ���ݚ�kjb]���Ё�S����B�IcBǑ�=S�N��9'�;]��ܥGE�3��mP�(�;-k�~(!�{Os��K��]����V?�Q��|�S{n�x2��q;��di ���1�_Փ�I������'�H������hM�.���8��<�x�i��P�G��N�f�hl�&��<P�_{�]����bP��@�F����c�0˨�V./���!L�.M�OCwB�K�δ�T�s�,��D��l5�pM�/�1��)���ﰂ���k���ӎ��7�M�'���;f�(�	������R1�H�Cr�:���q�שN�=m[�K�ıu�25GF?��t�h�z�`�R�#���ѹ �� 6���^�lq�p�UBx�0L��r	���\͜?~ǘ�bЛ,L����\�X�]΄:�q#��HdA�/w���-6�Xq^F��T�~9���?5&���"��{�:y����WɈ)e�2!�uH� 9J+�Ϊ�=g����=�b�S#o����)��~��G[�g
`�n��%5]|�|�!+5��5�$�B��G����7q��z�� Ks��1����3�j��4v�����[���|�eR� zDI:jv�p�jZ�	�����O��J�9�C��J���^B�g>�� ���|��Y��a�*sv�R{m��X���5E��0�s�CG�+�?�E���%٠���7��Wd-�m��}��6�z�Cv��@�QCFL�]�sbad��T���K�����{P��K�l�P���䴈��c1f@m#Ј����/��p���"$���3�		*bS��~�\��8mM6�e�l�ݏ�gL��Fp���]�$�_����j���a��?@)>�QڝbА��s�n��Ad��%x1���[Ή&�:����$p��n�������'��C�4�u�v���M��I"�&�����է�uĉPl�)M����G�X�hWЫ����k+
j;�'6���(��`硐3�<��'�G�)�Pٌ��r��O
ٻ��9vx��{�{T���a��!�5n�:��� )�����̗C�ͬ�WuC���qo`Xj�QRW�ʤ��H!IRv���L>�R��#�9(� �y�F�nJ�&��	8��F�!=A�����{��o��#��HJū`D��''REX�-��e6�?Й���)}/qLL�ҝ;��/Ot@7���q�i�ܲ+p��bP�)d፤�O9A�#�.��,��!��R��z���M��K��v ��+[��j�b��t����[)��f��}��D���7nފ�����o�>e 3�)��cHma�:�Mp����{4A(��Ļi\F&�4�a^�� ��vR��7�b�����z�߆B�y�d�N�.rJ*��xI��M�K��+���<��VU��\��_M_�؇vX=������-c}Ž�� Ҟ;G�n�6L�)/}�p6�X��҄{ܙE����w*��r��y�Qj�s!�-��m~�9��҂:j��r{�+�?��	����������Y꤄���ͅ*φ�'%�o�s�NK
d!(Vx]��?!�$��r�"s�g6��հ�����Ȝ��BiC�]��3=��y\��*]� ��A������e ��ڟ�J�{�~y��_�́]Uƭ+��Ȳ�!���^J|+8����W���}˟�s�a�!�x�G����&�I��=�wmZ�٤���\���p.E	%�F�`}ҥ��`�;��;+���h��V�x�*�3���³BH�������2��:]��e�R
�n�htU�8�C�@h/�nq8NO6)i���n^��aY��D���*���N*��W�^��T�	��M�&*�L-U)g��$�_U�GV ���X�3e�5�tA�t։2خ�2�b�";Ԇ9�e�������AK��K��K�8�	u��sL�=�[�N~�� ��4��x��\�c�z�(Oq��� ��s�JX�\����-��o�
��+��@-��o�O��~X(�4�C��P�#i�Q+���o�Ԛ>H6=�j�u�7�:]�:���hi�n������v�t������O{�c%蚙(Yd�����U�CXQ�����x��mfd�\�K�qh�`E�E��F=�6���J="�Ӕs�3G��&?�&O�|��
���꒽���zw���kѣ�O�
Z+^��NO��M�{�އ8�*u�^�;�v͞�_w�^�6�-�&�=C���~cs��Ic|x�Y�"2��U;��~w�G%;�s
>�ɳb�쟋�|FX�"|�#��=�ǥK��?��\[�������?!\I���]y��WĴ�0�߯�0S���r���������<Љ�A���g7�0��R�p�׳.�M��v�5	y+gG�X&�9��h��p�.�`[���e���ܘ��!9v+\b[(�"0ĕJO�ᡴ���ᑆ)Z�C�ѪN%�u���-yE��gTO��-��q>I>gt�lCu�p��}q@����b�%�t��S?�`#����t��dJ�!�U!wF��4���Z��N0�ί� 5y��u[�Z����,_zr�
׆�]�*"��:xx���7����41��H�^"#����֬���͗�xQhJ����v	�!��t9+���"���2Wa��ej
j`lrz	�v|�W�Ƚ�'��1����To�$�l�i-�<�І;��Ah3�/ǜ���/±$6�0ܽܖ䪻3e�j��r� HK�#T�ےy$�4*܅ϒ�#��������WT7_i�eW���E}�._.��HDƔ��Gä�q�Ȝ˲���~�H�����c�C ���{����	�c�X@69.�Z��`"79�{=��;�}dI��C�B�,d�D1��c|���Pa�1��.y�V�G=g"A�����?d����
m���b2�q��]��V5�D�_�ɛͼ|�M?�T2��H���ʎ0�ce�R{�M8[�.Uc�=�
���VN��&q�JPA�Ɩ�TgݦO�;%鈳���K3:v��Kg+zv}��S�7�>Ԏ���\���c7�Uj5�P��?�ƠټjKB�	�x4�׬���v�x�0$lp�������BqA���v�l��ȥE�fEe&�M����E��7�<7Y���&#�`��P}����x|�%���m��t��'��p�H��R�Y�58"m?1R
�y��������d*��ή���ȅo�~�ܓ3� �<�pa�h���7q��� Ka���,S����-f
�K���><��m��U����1��N��{������ȭ��:R�&�K�{WPU^~�˔@�p��hg~ٝA�\A�x-��91���὾1`)Bg�}ۡf��5Rq������G���"Kd`�kQ����1�e�_I�7~�!L��u�W�ś{�]�����Zs�K��a�۱��t���#ϴȫ�����5�`�S
��ȏ[����I�%,��Z�xq�W,�H
��~H�����e�1��[��>�-�����R'~�g,�/�M2,Z����O=)m+��MC�!�O6�9���i�!:�eh�Q�a���o�����hV/�s�`�-*���Hl�syUk�U��q~0ӫ͈SEiI�M�D*���A�[K�>{�؄�MS�P��H|Re�6���C*��� ��#�mO��;AR�<3Q��Vd��A}X�AZd[�r$Dٮ���&��)9�:F!� K��m|?�������`��ҩ�C?<T�gDA����I�����l)i9�D�Y����Ja��[J@N�Vx��*]ˊIb��X��k���P���=yq����eb]�G�<G����(M�vuY���d�ꪑ>�2�ڵ_Tu����
i���5�>IY�q�5�g�r�4`1�
��21�{v�s�ppW���^Ƿ�X#�<+�;}Y�"
Ix@lش|72ع�w���؋FŌ;��|�H���Ʊ�ּ�_������؝��WS����B`|�Ue=����v���X���	� ��Ee�Ё+0��`A�ffO�T�uX�����Ȕu�A�Q�_���]ҟerV��o��ЩW�q)�	�F}�`������F��u6$�>����Y�.��R]D���i�It�ҹf��z��q��ӛRb\�]d��K@~��C���t\�6� �J�(&ÿl��[k��f�h�����y�)0�Ir�O*�!k�Puw"I΍W�2W���zD�뿡Ŭ
6�yE%2��7#-����:2��a�٬�;�N�@��{h��
ژ�~!����|5\ג���//�L�;�@4�k�ޝ0�w��Һ0�v3%�(�Y�)6F�����]P�����4��^��7� �P��Lo��xK��t� �o�l,Ky��y�}���Zc�^�$\�1>���;�����ip��P��	�CL����*����}$���4B�w,]H�l��]�4	ř��:����'N+㛏j/����9 ����<A��
�Y���[Q-�7�!�v�0wr�O�f���M�o���9��{ZY;3F��2�L�0V�+�.[�o���7��jCU� �#� ���*�V��Q_Q��S�0��fGy�mma���/�[���"&m�@Kf69$��X��&�P��g��T'v�͗�'���?�A��\�Jw���ڭ��	Z�������Ҹ&LS�Ikq�v�f���a���%zҐ�׿t��X���x�����y���8[��B�'8�E�������V��bY��=ۓ�Z�L���OEC��P���V��������&T��pHT�F��A��_�;(��U?E�|{�E���p�Y�Ew�{���T6���g%��bۀn����w���1g� P��<�f���y�R#ԍ���)r�|m�hF[X��m�zq���d�G�f�Y����ϐ�4n��P���!ȣ��5�K*�)�3�a���pJW�	�jϟ�N��M�2���R�$k�H� ]]�;@A\��k��q����; �{���x�Rzw�ia7�A�=��r8ƛ���d@'��<$�PV�@�3�֜ Nr=�S'�N*�Bj)����z���wD�B<q��`K�r�t�����j�WO�P�K)+��UF�[��h05Y)���O�aj������©8��\�K��E��"����:�$ԍ������>��ۦeǴ!ٕՄ�K����\R�Ϊ��M�!��d8�a�Ֆ_�*��SE[�v�ɽ������?��YEAT��J�~���HIj�6�C̃���W��X�O���h�������Xŀh;�l&S.�+��!�B�!���XՏ�0C�����{=�O�����w�]$�'�;��+>爈�/kظ|�w~��4�Y���?����2�q;����|�F��z�g;xa�| E�=J�l�FkO!��bg�"�������"ø�J�K��l��
h���a�'0��5݆�U^!��B�dq���5�	%�>t�J�z]c~���5�;;a�o�ڀݳQY�G*�I�`�r��8�9Cge�����V���&Q�Q�G���+8�x|�P��7�^�"!�}��[Y3��ڠ�@D�r��[I�xB�g����߳85�T��( 7��N$1���Iz\�)ӟ֛h��Y�����i�8���2�{�1�~�e��2�$�H�:�}�dw�0���Nt=��V��~/@�׉�6�T�{���!�t����T��~�d���A��ȝ�`�#�sl8�=É��b��NW#�Z&0���|'n�(n��-�M�ك@�\��6p�6*	�G���n,d���	�QSÕ#w͑����wۙ��!*c_��p�Us�N���hV�j�߆	Oi~I&�;��$���
#��[z���=�A�^>� �*���m��ðԯ)����
Լ#�XS�e
���&�����k�↻G�]����Sz'X��bx5�X�#7{�yIuWQ��X��%�R�`&~�$tk����2���"������k��&X����8�� �Os\�\�;��DL��LW5y��J��A��xJ��.����3���T�� Q�g��m5!�=�����F�`�)s��2�c?]^�A���}-��ܓ�	l ��C*XEK6�v}���F�U>�A1}��dR�.����y	��^@�P�[9xݹ������3���ړ~�ȷUj$�'�^K�	�V!�x#�����>*1�|�I����N�KMՃx}@��M1㒰d�f���в����p��F�C���R~�������н.��v�l�B^Hr�`��4����x��"J���	���~0��!ea��<�^Ra�ʶ��(�1� �X���2L��GH�[g�
؏�0|�2-3γ���9��1"+�뮤��n<<@��׼�Df��Х��6�I}��3^�O`�v�=���e_��g+|L�e��bo�-I���\����&4�1�]��8���f�B.��k�B��m,�I䵸l��'�j�Gg�&���D��@��U��/�w��΅��gk@Ʉ*i�shx?��ώ���~KM��{$�>��-�I� �0��W�1AQ��N�1{�X��>.�:�'b��Xs�~; a>N�/�s̋p
J��=�fĞ6�'>gq}n]�V�ʭ.���,��꼝F�B ^�/�h���/��Y��d���`����}� ���B��Ī��x��_��Q<�F!�a1��<�8`��O�ʻV��Eׅ�д'$����|��l��o���@�KP�f%��'�l�N� ��-cLP3�K;~��-/g��I�?��§��Ѥ㑜��v�W�Y* �nϸ��(�q}v#QG�чC�3��������W�X� `���?D�	������C�j�d�9�0�0V+\��@q2=�W�O�>J�<ژ�JX��������M/���M�5?H%����r.�|[��(������C����ϥOW�G��=g_�lk�5��r�2U��gF�D�UM􆲡��"���T���gc@v�r����!b�����2��ګz\,�#0ecVLx&��x#=3ݔ&tu[ѺЎ�T�[�+����X-:��VĖ;{��*�5��6+YKu��$~����o������f�cE�*�X'�7͜9��0�5������sf���2���N6X�@nr�:t�w�&:����v�
����o�g�U��]ł�j����^�А���O9�P�$�J�b�,�X<��(Ɣ��8bn��Q��j@��|�>�ꂽ3
�ym���W>��-�������<��̼.76Q*�0����A"�{�J��/��?B���w�-i���Ww�mK����%c�W�v�}(O-�<����6VR�#� pqe�b�2��ǂp�l ��v?�'HmQAR��p�S����P^×����#���5˄�J�����aa4*�(uՒ�?��6%����Jп$��"���WWc����؛����
�|\�/)<��7�;��1�Ną���{��)�no�)�JA���2�q�]'�WU`=?z����)�r��R��S� \l��ߗ�M����S��>2E�Y}�\�j�� U��e+��t� ��;y�j�\_��-�*�3��W�;d��:C��S��[pNR�:.\�CJ�S �/Pe��|���;v�����Ώ7-R�eW����-)��w��)zE��rԳ&�0����6R�Z�`z���BiNOM�m���m(�Y�wv�����.K�g>?S(�ޔPf쑟��\�~IaL��	̀^���D���gD�3I��Y)B��8)��_ꁢtq�#��i��z�B��:P'y&�E?tR{h,/	�ʵ�6 �jkp��J�,X�=DY;� v�
��������;F`s߻��1\#h���� ��v�
��	
,(�����W�A��s$ҿ�*�V�Q���g�ho',�u��QR���Os��8ݷX�W�4?�vLp���UjX+[h��BtMܑc�)vD1]��(ӗ�yz�Qb�9�?EkoT�1"Y�l'
����fj0�?4U6w�cdȥ��vU�c5�g��"� j���0o$��N�o����!���۴��,���̓�S=��߱J��K��D�|��E�����"�c��x=h���(�*As4_�b����d���)	fׯ�lj3$d��\x����-�{�rT�1�F�������"+(���✹J�/�F�u����:a���3>;�,>/$o��A`F��!�)W�&g4-%�ݐyʕ
�A����#7P�wU����
��^����u�f'�pΙCe�M��o�|&
$N,	�%e�Ml�|�����;&��b�X���$A��7�v~��sG��ڭ�+]C�6�xR ���c^;���HT�C�zO���S��d�\/��"$�~Ӊ�*���" ���m$@�r�g�v����
�dYhXr�H�l�����O:����ԙ�z3�`��h������ǡ��D/,}7go4�/��T���3�}oh@U�Pϼ=�{L�O��ME{��0��i�'b'NV�$�T[cNN�'�m���)��&�Ps��8�c
�)4�gi�D�o�޷�������d�p�ky3�D��кG�,�Z�a20�E�1�E[�����ӓ <=VU�����liƆ�a��V�/!�S�:ܬ2��fAQ]��հ>|HMj��RQ��Փ��K�i�h����7_�.1�P��gq����F+*7�͡ŏtg�Ԕ|c'�x�E��:�Lĵ��]՝�i~u�)��O���I�j�K:�������E_{�#ck`� ?�n�����o�Z�z.d]s���Q+¼��>��)�w��Q/|���x#e�_޲�n&���|A~��'����hȝ��6��Q7�E�9y��@��:�(%��>W��P��4L�\(�e.!�o�.(-#�8^�&��m�q�C4PYd��mm��dwg�/�Ӥ��D�V��[�Ńo���`v������G��E/�������&2*��3� �����r�.[�|⊁�Ҽ���m}�E}$ת�:�Y��4'�4���@GB�ewr�ф]�eT��A��&�/����3�M5Q�F�ZلU	�RD�NI昗)���_�h���Y���*/��*���ՊCe0��r��I�j(w�E��/uxi��{������+N��y)A���yr{�:~L@��8T%�4�ǫ._S�X5�2��H�4���2TS{�P��{�� ���������X���k �Jv,y��:Q�r�V�mbg�R�޶wB�1�������AۣG�ש�J�B;��ȳV<���Fj8a�p�<)��:��ñ�x�67���@�U%fbb�)9��G%�L= ��Z$�B�?����!�X���П#�P�(�s��o]��=�aKkfm�@�M}�/�RbҾ�=��ҩ��i.����<�['�sk�a�����&�2����k���ە�BV��6R����04&��y"�:8!�B�n���=��
z9�k���.H-�u��.�C��w� ����q�D"�����>�Q�g	�AO}O�
)�	�æ�,y�6�9S�d7�)��\�v�8�;��GL5A����=�,q_mH����b��S���3�*� ��AmǱh��qo��-?�?2��"��Cft��u��NCn�����cn�3���#�Gp�rr|���h�{(�#b�z�]�Z���V����D��Ա��	�j����Mn��V�� �7un��~��ej��(���UB��~��z�A�|P&4P�a�!���%�r���ػ%RO��w�R��@���{���G.�1B���*�����w�&�:j^�R��{��.����b�[����0�h[��XT�O��md ի��ʟǵ���2�����3zuЕׁ��,A�-��������b70���������0岽ʜ�d��������f@����d$m��<��/��C0Kt�~Ĵr��C���Ic��� �@r�MHh���O6���G��M��M=ee��5�I��+]�g2ζG��R�6i��Qv|�wItM^,��/�ʊ�����xAg�V�	7N����f��I���.�1�55{���}??u�a@�w	���r��,.�$lx !�F"�d�h�#o2k� 3r�u"CHp�4jxl�W�v�9T��R� ����9�u�g��յnZg�7�YEA��	���n�^����NYV�v4�q��T�\fVwJ
�@�7ӏ��i.��a=iXī�
��'�M0BBo�����呵�*�
lƿ���(BL2��K�/g/�2�Oʲ��W�f�� �17�]T��ˬ:��"�ɯ���OԘrPeE�%��39�_�nV�ĲV���n���7�k���!��#�s�����i�W�뭗�/Zws�ڡ��Ij�$%�[��|a���#I7sCEJ͒Ƿ�}m��x�
,��<M�-`��(��N�]�|G�M���	��E����1ƿ���(��w��T��nk4Zn�@x6��ԢR��3����n:��(sh����]�N2��W������x��C��y�d<���h���2<��!���!@�݊J-z|�|2�I��ʼ~��6W�n:�T���r���>"k��J��]��7�1�	Z쇪A{���,�,ie:Ω��`K#;��;�,�pKEUy������e�h��R�}\�<xȵ.�)m���iW��#������ߙ�Yv���q�"�X���<&��K��r��ϖV"+
-������y���@�b�؍=�3����bT�C|������3�ŎG.$�:Ө_���A���wWA�Wud`�gG�/�].ւ���1T��,�<��l��nP�l����$�L�FlS{+�p ��txA���!��TERO�˄K>�-#�lbg��Ȯ�/����p�9�e*����b��Z���ߚ�C�)�1O�zloTEuO��K�J<�*Z���)��l��fy����Ӝ�Q�M�8;���0c'�dK�\&~�ъ��ꑇ5���Ɖ�ҝE � ���Z�&��:����	ͮ�ږJ/�^ECi��	��l.�tc�m����ˈ��2���E�vS�.���d�m���< ��{d?�����N��nޕfa�]�Vitw�|��	��z�Y4��¡��Gr9�����J���I�rRp�����[>��G@���9]Q,��()}5�$;�+�� �j�z'k���^ik���+(�p�h_N�bq�=�y��R#�!��r��b��ȗVa@X����+R�е��Vg&������;<*Յ;��_�x����-�*[���(h���4vW�
m/<̃�_sq��+�y���ʵ�FQY_�T^��7M	Ј#�K�1�<k3�׸�)��݇*�����u�)z��|��qF��/"o㽂��mE�~��(���cw��~\�md��m�q;�a��qu>�
�_��$��'�cȲ�_����$Zf��c�Ľ�埏өcH}������&<��au�h�*���{d �:NfF���Je}���֋@���;��Ճ�O�NF%m;\tE�b,�t��>s[ ������Tʞ&Msj��2��i��"��O�+���m�&Hܡ] 4޴���PCv\ˌ+y�=���	s �mb�'��8��,�V9��ڝm�����		���BW6E��K���Q]�?�wԫ���c9���;���sB]��qbp$���
d樈��C�����;��z���0���ȱc���_�J��M�\�u���we��Eds���	O�y�9Π4.�zn)>
W(��V���6D�Z��{�Z�.xθW�K�a��MA���ޒA"�h�cdOv�F��?��T�#�JĐ��2s���i�ݠ� �o9�gu��o�ٷ�d�&:�oğs* ~�B	������z\9;��Df}֍��R�k.�iůI�Mx�'`�BO��T���w�(�2�~�"�$(>�m�G����ep�oA&�҆hJ؂�ٔ�^�����]^`(.���1����Y��l�1�����L!l?�3ٝhcPLHHSR��?>�d.ۀB@�.^�9{L�>���h���1�Y�?��U�N�t�z&�g"H����b9�t�ݹ�/t؂2�	�;85���@iꈛ/U����f�0�D/B<�����i���p�D����b����{��Ņǁ����	��7z��=�� X��%�1�Y�z�V�E�3GÙ�̜��$��A����P�xܙ�Ma��-#�	���I�C� ���1S���7G��]�W���H��l��JX�nl
��|A��'�â�{C��-���ܫm	R�M��#Ճ��λ� U&S�����C���1�Tv�
�h�r1F�����ę���ڠ��]*� N~,"S{|�B�����A�ؑ��P}�	�0���J� ����6���¹��Go��z�Z'ط����07����f��8D�%�{�Qhnߪ4�<�M�l��Y�0��A�R��SL'��YȥBj:m���~�7��4��a�?��C��|��#{B!�h�J`���"H�sۗ4��������@����U#Ҷ[���&q��6���
��I�A�H[5u_ W9q>��0����9���Ӣ
AP�"�q�1���k��by��q�)!*�չ�w�l�t��(�)�(�^����p�i�T!�Q'���N���x�y׍���Z���p}�"Z��]_�=�����A��kr�)�,H:DW��6Q�{N�v�p5�?������`��BU��r
��WT�aXr�0` �	#�ߋ�&氘�C���B��Kֽշd͛h�e���/%yI�MfZ��@C���T����!�X���Қ��n\#�,L'kۃ����.E_�l>S���!�
���?R';@n�G_�Od��3�n�~F�f0P_�y���/A��4C��1� ��纯C.�1O,W�J�w�%�2T&Q�y*1��m�-Ãj#м�Ku�3=%���~`] �`VłEצ1	��Ns)>�S�[kŘo ��6�r�#�A�x���R�7����%�zﳏV����c�{y�O%�H�g�&l*����Dt.��URA���kr_
A�X�_x�
:w�F78@"��g<����h�ٍl�����:�dY��=bЁq�Gdj:�� (+��q�{�v]�w�� *�Q�~���װ���Pꈧ �CR��:v��`�����f��J���w��\p�A�P�����c �o6o�����ʎ��ܨ��c%�X�'.3g��b�[��φ���t?�+ۨ̃J�yO�^u�O pK)ff��6�%�_�.�4�I��~_�ݰ�����}�,f�(xҡ^pp�@�+
&�s�-(�����1�Y���Ǻ�"f��MR��5���N��_�J��]\z���_Q|�QU��е�(z��Y<T�����H�2`%h��ҕ�,]��.��D�8�b]"��u�S���K�',�}��Jآ�����6p��]ɲs.������Lt�b�ej����[�mۖ{�O��P�1�7Y�'��9�Of%]8��AB��p?�x�������}�k�#�@8Z*��U �\�^'�mqe�O̔c�P�Vm�� }�@��j�W��5P��{ '}eeн����LI�4�h;����>Rf��� B�[X��s��B}�cO�e���j)���0Ь��Yu��ُS8�[��J�x��o��ay�t��齸Xl�s��i���f\!��
kd6L�{h�N�F/����3�ȹ���Z�0A����F��t��pՁ�[{�ǈ�_�BVGҕQV�a����N�o�[̦�G�Y�Q���5��#�Fv��M��Q!g��L�/N�?�L��=e�<�d��=Ux:Z���'��
��Z��`��lq��Ѓ�Ǌ"�O@�dӣ�T�ѩ�ՎW���`�=���|}4��M6�y�ȍnK�E)��֬���Vb �2�T(���O���M��M�+�r.���/���&�N{�t4��ÇuV���`���G�}PXSTL�ݪ6|~j��1��=�&q���^� ��f|(�V�ey�=�&@���4k�β1*���`f|�Бs *�����?�Ў4�>��H�)O1���h�W����ĝe�����)�E����V��ED���Q@v�va�g2b$PY+Gw�7�ާ�bL�כ��M�m��+�"{�)�wƂ�
u����P4���w�)�3�'-*���Zh��'��O�BN3'���;���=J��9]U+��L�}����s��<��	�]�W��F��n�{h\�� q�����ȭw L�`K�L�����dڔef�� :�SŽ��GR�ʝ��S��t+^ ��T:�z���0�C�R�}����YwyEC�l�Yu�,U��x�E���I+2��+QcC�Nէ�/�P�o@��H���j�h����q�����38�^���v�!U���0��qb���x�a6ڂS]�����(o+I	E�nͣ��a��P<che�*���a�j6��r�n�v3�%LD�(�a4�3���	�%^r5a��M��T��/� ���|�S��ȹ���j�*�F!}�	PX['��'����y�h��������!�܏8Ž�kr��Kt��3�,$�7r�Ёe��-$���#��F�<D��g��F��T`C���I0
5��E�?
|zr ��爻���sq/=w�6�}D��.l����9�@x|�]9�b�C,��������~��R�gN����A_	%�k���Dh��b\���_���В�Ut ץyu+�
���	|PO>��;��6�#">���7�
�\���OaS̠c;4�9����p�L�BR.e�:�c�r��3��D�{�D7=\wH�rĜ�O����f �!�v�J���]����xp�FL����J�����p�$�8�JC&1�����-V��.������ɴ��F�byᯑ���T�O̻���z__�dPm@�YPY�{����Z�g�;�c�pb�$q�܂9��ԫ�@;-���<��/ZN�ސ;��4��
�u����Ѳ�m_ζlК�J�g��������s����B^�T��:��[W���.�m� �̰$��q������	�zW�z0���2B��m��u���7ч���V�pz�{���9���HX��q��c�8<_&���_�AT�|He7����:1� �ڿĹ��E!W5XO��-��J��7"k�D�=����Sօ�ˮ�~����Q�/�F�#X$~�v}.��L��wҨڳ�۠��8���(Ͳ|�Xg{9��W[1e#��>*�BG����mlUB-y�xn�*g��'�_h�_��0�anJo��O���؞�D�Y97[� ov�_	�t.k�7���Y�^���撣���^�S�ϘW:����a��?l�U��c>��=�J��zVuJhg����+����=W8�]��@,�7�_���ZUK?��I\C�v@ґ��?P��4%)����D����_�7g5�ٿ[��|H%x���x5JQ	ȳx�,0��)?�3�Q2Vr�PLX1�A�E��Lyz���	�p���0��j�=���W�Fd�ƓLr�%�p�p����S�{u�7 9);��v��$��hX'�R@�Ob����";�#����]�i�_���ں�X��g����˒;톽�F8		jP�O�]���m�vշF����A�@i���hؿ|B	8���n��������1*|Nl�skL�E��x@���HW
U�}0�>�|�\�
%��H�z-�U�����E���;�~�4s�l�r�I����h�a^�=�"yHmr�����8�?��i�#\q�&L�'e.��zt����T��D���8�����x�t=�Cu��Ҭ�}ߝ�E=���.@�bGD%;��E�nY#C��n\�[��Ƌ<!�A��!S���V"}�}��H9�NC}��ҀI�h�<�e{U����Q��4�׈$2��S���4�t3Lk<Nou��Ї��׃��]�o��|�)dCx��i�3�N�W4jP/yve�'���{�,��X�=Ŋ9���w���2���D�k��V��3&d���F �P�����3�d̽�M���sslNUe��"�Ql���>��B���Kk�n@Pv�@��Q̕,3FI���R��$���}�Z�>��nIu��^����$������f�~��]�k����֨٬����2l�+��-����f�#��_1�d� v$��^j��!T�%:y���v�|ދ�)D�Q=�!u��;����kq|T�Z��:V�X#f&�U����Q)�����@�l��e����Z�@�� 9�{t�BbT>�� ��D�����y�,srgo�T蔟Y�9���\䝱�v?���F�.�p�Y�`�����B���+Nhz�<eL��+>�s��"ꉵ��,�;䟊J��+ڍgݺ��o�y�����K���ߕZ~�naf��@���1�	WT[�����Mv���2��<Xp�9G?^�~<f*4v��B�?�k_���%��xm��vpC$#���Ö}
"u9��� ^�k�ȃ�4��#V�yˠ�y��r�˜�U�wzK��?��-�J����8㏈��K�?���O��,Z�v�6e4(g7�yD���{6x�;-|JW~���ǹ08�q�iFȡY�h�V��_|��m$:�r���ㅔ)�LAQ��o�F5�s�L�O�(+=�<�ѐ�����eP�AGo�n�S�`4��
a�8yx��u[û��ڄd��Y�X����68�[g��?��h�j�;=��٫�p����l���a��-F2���HJ4n#1�m&�ZOz��W�q�����w�bim��fQKk��'=n^͑�ݖ�	������}3��|K�A��?Nv�x�.�i[�D�2h�M.��u�6�6��$v���B���S�p��K4�r�-$�`(�1jt�4�����g��GW}@�t�DdoQ��ZhGg�Q���)�x����yK��=�)58�ސ)�wQa:�QAn���e�#9ă�y��$z���R�$0�4��7,l	Q.�8�^�V	�ރ����Eￌ� Y��V�+I������׽y�](�m�����X$6���k����\�e[��܊\�}x�]��gnm�:\J�+bp��?�a�"�k�W�]��h4s�9naV$b��	�H^��O�R��YF�8R�[�]��-���,�:\c>���	R>��kH�Cb��ʡg�x���v7��� �S���<[VG���\��/n�ߞ&`�-��;N-YB:�si��~�< �	��e�8l�)pE�l9��7P�q����@��t.��O�c	>�����ӋRy��t�c����w�����Io\������ݴ�z�_ߩN��
�������,Bw��$�Tb�Ǔ�2 ��l�����	q�gN5��9m��ѧ���GȲ��V-�ek��,{9+VWT���)�5��_�j/��S[�#ņ=� %UZW�{�2�N)�w����4ڦ��ш{�U'h�r��d�"Οg���>s/ٷ���[�w�}D��h�6����Nq�j�*v�,ة()��q�Vc^������
��q8��C���"�8p��2������g�]"D��Xڵla���ӡ+���!ty�S�Ʈa�;��o�nqB�� ̫�>� �㞦����w�z�
�uF*"6�]��ˆI���:!;9P�Z8!�pi&%(;���%�۾4*���X�'��z ߨ z~���a8׍���y�I7�w�ވ���ߑ����(�S��Ho��ƑLc��vi��4�n	3աYQ˥�
،�HE��B��zC���$"��1��z��+E���x-	�@��k���p�Eh�Q�S�u�6[ep�I�(�;�!QnE�?ֈ_�A��w��8	�YM�t��p ��(�w 鰗VH��"v���l=� h/��3��5Y�$v�Ds�'Au�ʲ�J	q��VC��e���#��<`�x��T�"{76n�����sÿ ��O����I��A����V�.�~�׮��
�w@�nb����6�����qB�²%q2󌩔���J~��`-������6&
:qslyHf�ϧ�~8v}���4�N��pA�� ��c
��~.�(�"5�uT���bo�=���QA�S��uԺ��� ��u��������y;�����C��,��p�7���U�`�S�?ڍԔ5�K�>���2C	d$~{2��菏Z�ķ���Y�ʵ՛Qe㗠������݃�aܶH"Y4-�����֢iNʟ\^�p$�0�8n�9t��C�2�"D�������d��>�c�-DY�Ѣ��O�Ӫ9z�'-P�'���;�i�3���'V��P
� �D>v��U�e�a�v'�ۘ�۟��Iq�	�m[�3��kv����w�*m����p�;�X:Qv��N�i��*)lES�RK]��� =��hGx%
~z+�i�b"��D�����(��U]�VQ�G.�$7(�%��z�n�B]&�B5K}�9�J�����;�A:����_���H�-���C�;d�-��N\��K���}��s��	�xg�,�l1"����'<2�Gq��}���v�NaJ .��	r�������)�g�y�7͹���3!OӺ��UZ�@_�-ġ�y�0?�?j�;�k3D8p�$q�K����Axy�d�&�����]�aR��+��A0!C�A�n�?x��_[�B_���MCns��'C�����8:K]����i���]��'_9I��ť�S����s�6�w�������d�������d�m��A��'��[G����o���S�h�3׻��H�*X�M�r�X��p�krߏ�]��2�٢1;�ɼO��-Q\U�?�6ѿ0�'�����r�)�V�op�h	e��-�����6�I?��tw���?=Ou��UU��`����6235�"�^�����х%��S�<�Z+�6�R�.r�1+����9zU�h\�|)W<����r�T�x��WG���8�H�u��"�޳C5�����J����D�`�����8��$�U�敒/�8���˔��|��!q!�wB1��Z�u�T�R�h��j��&f����ѹ�M�},&B��$���ߜ��u�U��*DY!�z�� ��Y���(�����c�Sñ�>�!��.����B�QF�mR�~������DK>��W�P�R*�j]X�r�/��2��Y ����4cJ⑥����� �q2o"�|d�z��Jr��s$C��`��0�Q7���p�LD ��J��}�pUܬU���0*�3>����{I� ���7�p㳩qZ��5���JJ��-�e.��a3�l�gp�Pi@E,:!h���PEIDy�#�'�T�*��/X~��Z{׻F#���
m�\L~X*���do�:x�gJ!�j�\��2L�b,���4v�#g��G0pb���V���=�;#��\��`4���'�-�7>Ck0RyTO�^�@�9�MT�D�p�kT�.��z ��!OT38��;�����ܰ�t�ޯ����}����)޲��A���Qe�.��=�p��鑫��hZ.�d��&�����b�А�%d5S��Z����ҙ��j��?*�{��8H�w �Χ&����fR��'����J�eF0���"�[����v,8�/�[ͥQ��fq�Խ)�3�n���������^{Pvp��~,��7�B~�������AȈ'�Z����4�7p�p�gPҌ_�hp'���^�u�T9G�o7	{�a�;�WX����^>ى����[U�����Ǭ��{�\"��"����J�E��Ƈ���N��1K�E�?�����[�1�.!��
��'�_ u+�:A^S���>\.�t��|gx-U�j����Ѡ�
ҵ<�r̤ru��4��*�����T�Ȼ�B^��̾]f�U�A�����(�~����q�bJ&��Qꆅf��.�a�n��H'Q��~,��/s."�/ޚ��,�V)���y�VO���ōd������4����4���6Fޓ���5ऋ�
=��Yv��f�˧M���bJUܚY��8b�����KXR?��O���r�O+���;����'��I#�>A��?�%�@���&�s�F�����.�3�9ʱRX��1�V�9|��r����R��l~�Ё*@`+�ב�����(��[�t�&a��d���w�qV����=G����\`�M�6��R;R��FJL����<-��c*�Hg�/u��p�����p��ɾ�K�:���rA���fZeZZP�[����;]�+�K"�XdN����u�p$(�n��ښ$�-S5�WA���H)��q'��팼��9u]6l��{/Z-L�f��PS���jbi���G�~5_{$!������l�3R�:�=�������"�q'{�Y�AՍK(�x��=��3�{�n3A���_Ȫ�}���!��k�y4���B����7Z+o�y����8^Xyt��&�{���w���5�aJ�"AP�6	���05�e����=�O� �=�0�J�~c���T��J*���G|M�Դ����'��%8�(�Y\)i�K#�@���h�d9�ˡ�;�M^�%ɺ��jb�����7�E*o^\)?���~�'դTS�xHx�ղ`+o/���Y����yT��K������
�%�IM�j�SvP��37J�{�{W}n��P���v@�ژ2���&U;~N�4��6۽Giu��}#�{{�W��$p������ s|��!Ҽ[rز9�>,��D[Ļ��Q��I[+p�����ts|�M���s�Ёu���>Gjh��� (�'�q_��_�ۀb�ϑU}�ʤ�vۻs��7�+vV�u��H,��+�[��2���%�F�wCM���To�B	�6M���2� ��)�"�0�-S˗�:6O�
  �wh������jxJ�,I�Q��u|D�+�f�w�e�SݝJ��$�_��]���s2S4{���e��H��Z6�,�/"/2�m��0V?��*E���W`����v�%�H���[�[5A�G�5#�#���~7.�W������ppĻ��kDMwA�v��0�NV���ۿ���������QRӌzA�z�_{�vv�vO�A��y Y����`
7��&IIѦ����T���p���Z� a��䏾'��%�YDBF]C��_����c�щ/��D�dH]�3g*���!yc�<�l�eH��=����?�͌�|��D�X�Η���Zjӗ��Z\ ����6-���>M冥cHh�cb�2��?�ʆ���\��C�҈���\�3��Z�2`�ٟ�1���Y
~��������; 0�������"Q�;�+G�=�}�S��n�ZZ%Ya����j�*�*�qClf����� �h�t�6��!�[��~��DZ��U<A�r����Zk�K��^�*�z��ߡՁ:~��[�:��Jc �����3t����o���>s�:��N���S���4>sx��^h���$v{o����/j��������9��%(��<�ݢv�yʚ��.3�L/�p�8��6�SJ��}��鵖�����D>bG�:̒��]F�׺g
�bd*�����(�TD`_K���e�%�(��p/�"��˾M�Ծ�]+c(^\�_p����Ɨ/P�g�'ēsL$Q��_���'����o�.���t0��BU��zJ7.�i�g��(��ٿ��;%���38�����~���m�->�h�i����#�h�������ҁ��xB�N\��r�����e�(��/I�%���c���'n[ Φ�5����tҀ���H��>!�X���qg$E�����_���!���g���Tm{��r�(�F�V�m��B+�
���
v݇bd��R����k�@V|q�ڻ&1C&�����+�F/3�c� ���AS@%d2���m��?D�]�(�8wBy�G�(�0k:��D�9�CF�AB����B�[���C�#�F���Y���ݔ]h��r�1���=�\�"T�AB�|㦒��l����ie�N!Fީ��7�UA@�Ԟ|��ϒ!�z
q�j�p�*��%.ќ6�-��X6�s�*/��L$la�q���#
��j���7���x���+��g��<L'�����!{���E����&e?Ѯݑ�=����z�5���>�"�'F�%���[����P�L�E.�jI?�/td骝��X����&������V����r�r����}B��1�%8��G�j)Bhi|XE*��,b����.!G�-�!zgRW��*����w9jzYK�F��?�<V�V+k&�
�q_���Z}�V���&��������m�rJPѽe��:��+��q��R�A�k�Q2�
��+�!�����D���PC�E"��i�u�v{&#ͭ>�k���B�Rt��ᤘ�av,�81�?�za����<ۨr̷�^��4�h\+֋q��_]!���n�_�im��S��iI\��c���1>��*:�G��na(�%�H�B곫5ʗ�ʵ�����<愢��mtX�EL�4U��~��MP�&Z󋙈���,�����2ޮX���l�8̈́�D^��w��?Gt��F���������'B1;Ī�����NTvƗO���8�A�B���i!%����}�����������= ����8T��[�6�Ly�(�"oۣ�ݒ��$"�{}y%7��Ug��kNV�ĕ ���ʖ�B�z�Zw�Y�:-W��ng.U�mn����7[S��2��?h��*5�MђJW�h~�*ez�%��Ӎ�H �=��.ϭ��h��$��(��b��Hj���v��ӝ9,����Z�98��0���x�I���"�����z�N^��"$+�Mo��|<`U��?2��+",�\�HQ�1�-v^�WJNڽ�%�R%;��U��Y(V�%Y�Z-�u��H�)���~:��1�����O}��ßl/v���D��&�յi���>OUHC&�q6ԙ��Y��eO6 ��j���>�M�����:��I�mM�qjj�5$ЗN▶FMQ��Pk�.ǔ���J�3�r��6���� �W�Pbw���w�>�<� "`�t�t�i��I��
8Ъ�w���R,����҄*���)Jrh����64ք3u���b7��K8� �ȿ��,(GǛqh3�J��h7�{wDΐ_�F.�!��¤���{����Cl5l�K��k%=��f`�X�86[��~���*�&&�[搨����؏yw�oTC^blZ��V�XnE׃��_Z� �nO�C.�	�A���Υ��&������4��'7-�)|{^(���!�9N�� �uOw&Gc#�j#W�8͎9ƥ�u����`��@��DzQ�v��A�3����z�g�.����J^\g	��	��9����VK��lB�Rs�
ƫ�jO�G��Id�R�H�Q/z5�\+�Z��ߛ��P#�j�ɬ%g 7h���U8�+�3�}֍�X�쩅��Zk�-�@˝,ǰ�}���Gx$a��ժb7�:�g�k�� X�2�t��k�%W�7ks���������u���R��d������@g����}�Y�N-��$Y�*�LB��:z2�[q���2`�Y�/ �\�g������r���g�[�����#�Hq^x%D�#T����%��蓉[�):�/c�x�:#�`��}��K��|�B�V4��Сv
��h[��ix��V�?���-���ײ@�Y���4#���	7T�N�N�	���4�0�Pŵ��1�/[�,��7 s�>	���}]l��#N�W>^X]�cH�tp�(Z6�dtǩ�8��)C*��`0��U�.��b������r�/r�QD˅duR�K_�1������� =	|c/�8���y���4������ӄ������\'�C��؁��	�G�4�[��	�T� �\�͑��~�H�#ʦr�B��R���eLo\�ܪ����Ø�n}Ԓ���x�¨-o���) <���熚�t��('�1� p��"+��e�&/���oA��,{�ƣ�LY\`52�:���X؃��`9��@H��%H�.�_@�L�&��q�����[1�XQ�aբ��Do�q�1�In%|��X�KL�V�O y���tG��^��0'H���Q��6y�G\#�t8�[�g��bۜ
;��Y7U�:��;����S��Ņ��Ӵ�l��Y`��e)!� k�Q9���!���W���@�u:+|��[Խ/���+FPp�%D\}��<^(K�!�0��e�h��2��"Z���0��{��9ߤ��*}o'ɽr��]������~SweS�A���p<+�Dw��P��uW�0%����1 �A33-%��@Eӿ�u�+\�u��h��}g�M������os�}iiw�����X��_�8XgJ�����MH��R7HJj4tG�d����	m�H-��D��
%t5����<;ԕ���� �m��4�Uv���n�����B���U{�\���Ù�#�*��p��SwZ�x� 3���Ho-㝾�� RKXh��;�b��Ɓ�>���YY�VF '����V���Q4A�:��hi�����(#<o�;V(��jc��V$�ʊ��N[��R���Jf
!�8�kT��.�g`?��pҵ�#��{܋ovYG�k���J�����pyf��35�J=11k}uG�I�|�9Sz���8��0Mb�.�Fh����a<�5g�18^��i��.ϭ6�����*��v3�j�6Tgӗ=|U+��6���BӦ4tǉW���<��٥e�"S��:�?���U7��i�z���7���)��U����I�x�j���M[7�b}|Et'��l5B�;j�����������^R�%8���M��5�sx'I�.��nY>�ObŽ� 
f_˯�=k *��5�UC�>���y?6�ٓ]��؆�U����D�z��?�eqT�)�F�I�s�L�]�f�>AYi�����N�$
�`��7����d:�K-�J����jذ��EhP�$�B~�,`�0���O�*竢�Y��h"GߜsX�>jR�V�U��E��LQE��Vσ�}�`1]��SQ�4���h��+h mn��$+��d�J�:a�/�RȤ����JB� D�\�6|�l*��O�=�i'��-o(�9�q�y-ISK�i���z���۸u`��ѭ����ݼ��>ɣ�e�A�\h��`e��X��VxV8rqP��ʟi��.��z����A�c���r"b��Sі|.��������~"� 4�$�k��B,�[Rr��,�Κ�!�C�������4����t6l�<bΆ���~��~�VaM��f�f:��7���~�b����œ`?;�L^��d���vv>@�\�>^�jJW˕�J��/�T�D�*�E���܌����L"u�uvFE~l��1kg���5Aא��� _v�����`�'
�r�Bo[��ܩ�A��,`��� �d�%7{�H��W���}�u?RcL
ّ%Κ��������k���Ga>5��l*�-9�E^��t��!�4�>���[�)wS��@q�/&����צDP�!hFz���I�aSXr���9ӊV1�;.X��N4�O{G��$����Zi� u��k�����_� E��˶�xY#��������R��9�M��0&{��1C��)7�:(A	��z���t<�r����7hGG"X��n!@g8��A��O���-/�F]���O�3�[*.��i/�&ϼ�с�cA����8uj8�*�)~���XD�I�~�8�7-@�
�)��#�	Y��pM��w�<@^e ��f&V�����_�����ᆧ@V�j��Vh���B޵���Uo�7g^�W��ن���֗߂��FrV��}���R���7�J�>�;�.1&�z��DI3[Oǅ��=6������_Kf�XE8~��1A:#v.�ӎ���Qp�0��u���M���x�R��Bɜ$��s7�e��_-؜� n?�S��\׌ʹ���K?uiU#~�,���1�*łm����b� 7��B_ҧ��sj��q�l�_UI�o�Zm���ՠ�tМ7���m�H�V���'���P˗p��u:h ��s��B/�?�D:{Dg1��6�N����3��Y-8��z͎xs�c���x�%�B���>p������P�gC),��)���fC�1��F`}�Lo��!���^Ǳ�B����8�f����l��2��w(�a�s�	.���~;��z]����E@����{o˷�q��t{��4��W�$=�7�������g�-^��ٝ:���'�v4�f�uϜ���#�������Ep1K�
7d)w܊�\d��(V���l�}���kޝV��׻ˉ�hy��9�ȍ,e^An,��;��_�vz+x�[���-���b����ţP�����̵� ������=�k�¨�liW�
�ַvq9Ʉ��|.�?5�f���nn�k�;�n2��R�5����aR?�
)Z7�TPr�5�#ӥk�
�:�z�M.L3�;���s��#��:�~�����V~��L��G�:���q22� ��Uf������
	����������-S	e����QZ��'M���g��R�|�7���mJR�_C�-D��{��ĉ���q�tJ�ju��(�Ӯ^�g��1�v2�,��]��J5���­��(3C�jk��!���]�}��A�h��<���(�Y:��]��b���=�p���À-,Fp���'�?O�r��=�e��,c!�:�È>R�?b����;K�2�5�D*;��Acb�iW_l��B��KS'܃J�u P�90�7{��	9
z\Q�Y�b�wpL�g7�28眒'5F���HLh��@�h�F�P�Y#t�3{�&�9�r.u�A��8�v0R�LBr�f�pJ7V;��=tZ��Е9KJv�:���aU��»�=e�Xn��b���C�K(�(��`>�ku;�Y��~ʔk�u�ϊw@�9/��D��Pn����J���hԆ�8�I�K�j#[��^@>��pF_��X�?y6�����Q{�)����Z��E���C^ˮ���eC���1J�F�b��@;w (��c���z�O��Mk������D�ގ�Gr�X�UE3A�`<�͔��&E�P6�˚���;��+���\��Qɩ�f�q�13�![<'�P]'3⋟��VFI.�@�>bNAu�^;��~�~���<5�
��E}��&���&g�N#u5�}���w�h�*��"�n�f�	'�M�*��@5��9��7�&�C^�gl�7��xA	0��\Ř^꘭��7����曟�R�V��ey��k���BTĴ+�+gy����Q����Kk5���1T⦋�;1��1!qnf-�A/&2r�ԓv�j���N��=ŉͻ&%��SLt���I�K"p1��Aܛ�?�H�����"�i�L��K��n�̏>8���k��	��{?Dֆi�K9�^��:	�ÒCȗ�+`Y�K������KN	~��F=�/g��}�|Zx��mC�(K5�_�&b�uW֨��⧎�V�M���@��� <�Q�p��/sH�\ Z���G?�&"aVy��S�9p��Ge�m�}��TP!�/��A���ɜ:V����G,�����G�0���sP�v��(LpP��d���w�T������2d)��'!d.���D^�!4tU��*�������"���#:8�wjÊVy^��,k��{իO��[�W�����3]�g����	�J�3N��:�Ut,�	���%`�o�n{ұmKg:��z���x�{����Ŭi�!τG�9A���AP�7c2�|�Bˑ7|�fM��F�!i5��>�������L�K	Xl�_��eg GS��O�Hx��3Q��4.F,��v	x~�h$��iJۥ(߲h�O-o� "�C�g�E%�v����-$�x�` 7�Oy�K��ܲ2^2��ÍN��ݙ��9Eʷ.�z��ږ*^��IN��CXq��Q(o�˥���;:[��Y���{k@꽅����ԭ�J���&�չB�u0��)�O�����Be���e�tыV��҈8B!�3l2Yg:�uT���v��?��]�R}$��3�`-�q����٣_��kk�{-9h ��lɭ���ňF���6��m;Vdl/��v6�#O����Spf	 %V�bhD.��>�����b�	
ҋ�r܍24��O����,t$�R�H��a���� ���L��Ɲ�K��2}l��w�sWg����cUU�JU�����y�ogϞ/���z]?^$��*�"v?�����@�z��3F�����t-�ؿ��%��	�+�ڷTӧ�2�f�K��9#���z��Ov��%�n*���9
���O3���F�CU����*��J�̙.�潬yѽn��p�����5r�e,���B��Zۓ����=v�K��q 䁛�����C���&{ܔ/����9�v�V����]GI�]�ά��G�Ԩǹ�HL�:)A�n�\�������	�GU��Xk�h*���n	�i��K��R�~\��������.�	x$+��`y8XuŎ����?6V����x̢%��x��sLz�4���/S2�ܮ�򢘢߲��*����ނ�`�a�2���������Jq7X�C�?�ժ��V�'3tW
�W�6>��#�1W"�궄��`)�TOV����aZ��MĤ���G�c[�Y$���$��^���L4M.}�o���O&I�aIA��l�Ƹ�����mס���E���H�3��/�m��ɠ�-M��{nL�:R�b�t��0�ŏ�_O1�,@Ť��&GH��"�'=����d=lf��R�2���R�k.ٱ>�dq���V��ƺ� I����HS�ۺx0\���
k���֙9�,��At����n�* S�ac�w��>�'�ɗǔ��9�Y�+��{܌��d�2���I1!Z�꿹���Ń������µaG�l�
�R�1y�<��ut��%o��u<Y���|��h�ی!x�����	�W�FI����T,��J���pF�`k�*}{�]_��Lnc�ڿd��1v��qg	�hG@*<=����7P�wC�N�h�{����w4N�~��o�8�|$�򯪋�7���Y���0�0ٞ�jN�����n��} K�)b�Ƨ�KH��YZ��3��Α�̳��M{1��J��^�v|~Cb�EX�?���?Ϻ��9��:'�@f��"��2$A$�"�.1!gN��YH���5SMv/6�:y^dyo����k�.fwć8q����` :L<�ꗀP	q��ti��;�@��a�#k��7�nڑT
M�N�%�H����T��7ɪ�ɰ"��_d��N��g��{yY%�ۭ��do.n�5k���Rٙv�a�,���P�nk��˚�DA�*s�A�}����$K��D�\�m�4/#�̥�1I�r����������g�)O��qzg�`2���	h��l�m�?��U��"P��_Yۆ�$˴�M4�����J�n��<O	(�f�;��Y���Q����Ye� #�=�S׹�8����w^t1���9���Yw.z�Sa~Cȸ��{��u<�(	������Ӗx��yњ��mo* ��^c�D&.Brx\)[C2k�a�y�FUk��
HD��l��mgBE���qnb{"��&��d�R���Q�+quQ�V:�X�U���k/�LPcD���;++J�0��u��Ŧ��(zV8�=k ��L��Kt5�Sy�7�1�nbL�\/_xq�!SL�n���ỹ4{Qx�i#�߂}R͂9 ):��G�Զ
��s��-.
��$?����E�w�=�Nh�� ԝ�m�^
!��,���¨j�u��-X��_:��Z�L�4��.�%�H��1��Q�|i�K�����j%;Ev�>�Uk<eH�ޭo��+�: $�ЌXN~�Y�i��� �R�d|���L�vl�?t���5VA:p7#���;��%o�:�Aø�d�Xa���u?�ެ]�8?4H�hn����X�-�n��ٔD�V��{z�{�t�g݇g�1nMm���	uvr�8n���dp��'9�}�O�Z5�3\���y�G[Ѯ�3mRƲ!����"WR(�;w�l_C��x�C�y�#��!J�V)o>N���|�5��n6�H���a9w;,Tj &�*�U���U�'[+��xV�.#҉X� }F���z`�e+U��@������Өu�Σ[����e�^a�ܚ0���m�a��982XFr�6cz�F�7��U��lŽFɮ�=%	����C0��B}c;՗���磩仃θ�^"9�=s�N9d!��)�� ��1�Ĳ�����q>��S�}��ӋY'��y =x9y>{2d)�a�ڐ��0�h���)H��h1��P��=.�4d��7���L�*�u�����`��T�������E˼�w�C��d�>uңG�x����,���K�Hi>?};���c=��9eL�N�H��&�[B�pr��.g� �bQ��#���d&�Vݐ����-���ˆ��;|�]_ZY^[N�yy;�Џ*��fA3��1?-x1��i�ԡ���������Bd᷍$\���'��r�an��N
�0�} �\w ���ޔi�KE��A�DOQ��O���h-	@���V��^�@�W�(� }B���@��p��뤥$��Zd�����s��a��tm�W����ɶ��~����^��W�+e��p��N�N�@8�~��|�}�V�냼�+o�7�2�y����T����n�?�N ��A�T���B���H��������e칷*�	F�f�]W��p�͠N��e���h���Ԍ=��Q%�	+'��2^�WĠ���ڈ��{�Mo4'�4���i��P�tf�ʳ#^ALl��	��6� 	�p�<�G�1�	����d9d[�+VI,�4�PY!^�ؿ��8Fnw>�� �R_l�z�Su1k����x�n;s�%���ORB�4tB���+�Q�҇#c�oRcs��s�c��H�B�q��/�d���v��;(��z2"��IN���臛��b��'ᯈI�^���0P6Pvo)F�f�ZQ��K4�-�{^K����4juv�}Ɗ�����pJ9ԠY�.���!��Y'�4�����e��O­�_�j������& ��ʍ2����?�8|�f�?��&�ɜ�>6�惙�8Ԉn95�\fϐ���<\��d�RɆZ:ӣSZƫ>�;��o���#�m��{gޜs洜�~v4�Z���+���&c+.$��=/�OD�O�/|�w��{%�c���L}��-�.1�������r����l�v��Lo��vX��\n��2Y���8Xg��{���U���|��9&�Np��r&lc���8^�sq�ӂa��Sr�!�kv}�:�l:�.�l��).��aQ*��B;��������m?����e�W7�E�aM��s���G�F�Nx�Vosb=����L�>q��&�J<�&z����J���!v�����ϕ�!�5�ȍ4��Ae��2#ts�%k���e�T����$&�doݑJl��^����?3ϯ��Nʑ�3�K���&�+M�iVM�^����']�#)�*��V�	��p���l$��XB��Yf8(�m��e�.['��yW���wd$w��b�6��Y�@�b��5���3t�u������4&qO�_���\w�Hk#Ƒ�;��2�7+�5�uJ��0��"s
I-F����K�?~,��g�d�*�-
��/	�j����u�&]�������Kr�������M%������s��_�y��n|%z[dt]k��Q�?���'үZmۮ�~��%g�	F��18R���k�9�ײ�_�o�>�P6��
\�)HP������t%��R�|IKK��:V�")� G�`D@�F��A0��S/t��/�e�X� �wc�!�%�;b�0�x��t�O�I������l��#IrM��������
/��x'���ZB�䷞�O%�. qرϲ<���R؛3MDAKh�eR���":���h�*��}?α�ۚ �[{��6�}K�b/�����C��"����	�]��~��k/61�N'H�F1���u�_;ȧ�U��G�.�1�ʘ�VU
i�������
(�<wQ�sc�C�Г;?2Р�}�/�����affk�7�f�
&�Gɹr�*R����5�X��-}!�:���4�0w�DW!���bw�^��U-��!����y��n%�1Wݬ�vJ�����h�1e_y�!1KvE��`��ō�7|01M��Gh�3B�0�<F\�����Q�cs�u 4����rV�9������h�WnyVx�$z�.�O�W�s�Z8�;*�x[H�U�c;�m��e��J=7�nEF��
e{`��G���qy��\H��z�;�?���������L�P��g�iwJH\�t�e-��5ؾ�/]��ǊTgc� ����d�2���'4*�G)5qA �>�Ƶ"x^�`.�V����G�	&h]	_�i<{��l\z�q�%EN�A+�]�`t��Ӥ�31����d-#\/�*�2�2 Z�o��6��=8:��;�>�}��Rڟba�D�p��,�*ޢ�C
�H�':��1��*i�- N���6�8n0g#�H���Ȋ��)�ȧ|@�-�*���\�O<� c�|�������B� �A�M�^����ُ������j�M!��z
��k�Έ��_6J���u?�Z9���	��X�
a�#W�y�:�A��.�5�(%@�ņU8EU��!�i>")��n��2�ߌ#=A<���l���E�2xk���Ǣf��J|A���
�u����M���j�0��mV3��+U�,*3����@Yf���3��,W/�P��&���V9�CC�I"+����������1mD�M�z_z��P�t���zs�W�
z��e����B����C֡��$&���	V��7sQ َ�Ŧc�u!��nOT�8�h8�^hұ���=S@z��ݤ�3��#� pV`H�jZ�>�iG�-�#lP���*^�����T�tRo_�[�=�9b/�`��0�ގm�#�R�G,þq۔-	��PhG�~>:�ĪO�� �����2�hoKf�����T����=�=,rԕ�M�;�|��UX�eٴ�a4λ�Z���٥��S���9���G�8�CYt�����6������9O��ȕ��odI�KB��^��eJ�2�r�@�-7���_4)�d�ƃ����*Y䭰 �|6����_oc��W� DH�z5}���!�OQ��:}W�!:�b9��j�RXw\&{�8"s4�I�ǍU@֓�xP�l*�&��ehg��D�ר���C��~m��X��J�P��*����8 c��m�j�#vU��47�1�/�a%^֨ā;�rw���W<ޫ��b+oʉ%� L
Ku<#d9/<�.�SP�Nͅ�)���5xY�Q��E�$y�0��Q��a��#�2&������C��s�c
E�@�I!����堍y�Y7�b��)�]�O�bN��Rձ&��h7�j�x;��E��D�-ڷ�ص��Z�[ca�U.#���Y�'�.���N�f�rN�4ZQ.��NA�c:ƌ�G�}����+Z������,l�\��2���Hn��:͗��)�_X-]��[��s�I"�?�bI����5_n�Xf���TanU�F���ش�E��N��@�!>���9�s-�l���5�� ���"�A�j�����W�1X���y��]좻j�������?)�2����	��"��)�O,b�%�!Oy���%����~]���7���n5�4�K���7�~#X	�)��(�����O� �2�RW�mg�����Vt����O^���L+�
�44�����p�V����ta'�5������/�P�I�wE�ɢ�W�V��� �&�K	\se���P����S]���ܘ�yi��[�\yڷ���T�Cu3#U=�,��U�\�ƌ�K_'�{u�or�E�̎zp 
c��e~�R.�0HvhM-�9�v	@��M]YY`Yq ��C!|�J*���OW٢���,fw�D#E_NCM<����j.a�Yo~}��ݰ��ϟ�(g�td5kR��j:wQö
���g�Ci-��U�2G�1@��K�7>'��Ej�������}u��	�P[[b|��3np���4dy}r�d~	�w��_r3}�fK��H��%n�U�~�
��91��l[#�|w
 !�,�f��e:�u�SCA']���nF���(5��v�E����� ��,�")��M��ø��}�ʀ�A�KԦ�(��Q��e[�"~ �]�^j6�>�}z��t	x�M{!���JzG�(3�5'�$��J%�WfW�@o�l��:�����H#A|A|��o����{s���(+�n�	u��F�P��s8_*j���8�}q3� P3���mY4[����>f6m�_��vG��O��n�3�/�yW'�6�yj�Q9���[V�����Ҁ�ܶ$PR�Cl��b���,��|��Va��] ��kJ2�ܑ��Q�Ʋ��,��+�:��^2��JH��:[�3��-����4[˫�2g�a����{;��.S�٢�:_��*(��W|hP��ni&��ܵ	dQ�b�ڳÅ��I󣂗�����dmLq��`�eK彍��A����n�_e_��E����b���潮����Dg�[1Q�h�;���W����+J��0��"��G�b��g9�i9c���/\��rq�������c��G�S����{h�r��#��YV�
����6tm��4��alWy��Ex�#�0������/б���]��ZHa��th�o����d�s�weZ�t��ᬬ��P8�F-5x��a��A��O����_��bF|?+�ڍGw/5Dk� ȟ6C��!O(BUȲx���Qʡ�3�[g����U� 7	c<����Ì<�	�<-�I	ٲc���t{��R&���fp�ws�˘<H�Q��9��aU��N�Y0�j��m��y�q~/b���Q�:�V۴��j��2fB���$e�:�bf��!O��j�W��I�L���_��������X0}����L�1���ۍct��M�e�^)j�
����ױ��6^48b��=��0��i�BV�v���Q�2a*Q����$J���	�7M�<MgY���U\'���`I �-�Ud���7�qW��Z&�Ǿ���/��E�s1
xi�Y��9�:N�Őcj�.AH�n��X��k_>M]��}����w�c��ӧ����%~����=��|�z��Gu���tIƦ�R
�
�.�Ӝ+/�pb�j��
��2T�$�&�Q���h:
mMBC��Ղ��[�����	\��+g�?�O�}�ژ}@OK�)�%�6Aq�4Ũx?�s�ȼ(��3��\��b�����X"��%aF�e=�h�"�'�ޚ:�������,�㳶��0�a�g� *ǹ�[tw\�|�TB��[�
��cK_�(M��~��i�_�Wx|jz�&
����5}!FIV `��z��s��ǣ~�2��Q�Q�k͜��Y�|t��B����3��%���6l��^k������f/�5CP%� ���m�ÚBj�UXZVa}en6��vPZ�f�F����5��P��#�	�Ń�P����m����Vl3R�Զ�0�e� ��T��D������;���$i���ׇs���{)��8��5����@<{��%���\��1kf�y��?Q��H��|��v7)�����܋�� E����_piE>�?�{RCud��FE.)ȸLʩ�r%�K�G�]p����\�A��0�����JP��{~Ɗ���f�w(0�2����cj�k��4��me*���j��=����h+ g����m��ؼ��k��phw;µ��L��A�}�8T��"*NZ0�x�J.:���Ѱh�
�p��=B��7j!��L�.���}����DG��	O��7ƪ`��R����X*3����^->n����w�(˓�Ǥ+���̈́g�`0�)�b
.�̄����� �	.���s@���8T{��.V
��?J4rP=*��U�~�1�'�����F����5�Ԕ�@�5�Pi��H�`u�:���8��4�]
ޓ��<��vZ�>d!%� vK�Z�l�B�Pq�	X5+/���䉕��^^G��!1}��J��d��wL�j<�	ڛ���Tl�[�9񄃽1k�Ϳ��1NB>�W=[�{0o�R��^���X�R(8��
���%S�ZW���e�������'Q"p� �"`�+�?���B�2'��SJ[����W�s�@)m[z�ӔF��#��>B�1'�+�fUdyޔ�O��F�OȦ�"F�=�F?a����m���ҳ��x�Y�8Q�Cŀ�	��+ߔA��qn߇%�����<�N�>��)�6^����F�=s�S]J��:�p�en2�0
��j�ٯa%҈k�n���.�8-u�.u˫��:箚B��h� k�n ^���.�4����]⤝Q�p�3M�-�.��o���4N�d� ��~��AK�;@���[qf>��X[�.���t�O�;�����x������ >H�� �
=Ă�
e	��p��:�@M֒�4�u�~szS�D�Z+���U��z@H�J��aGQ7�`D0��\��Y�g�����V��A�ZN�vױ�_|����P�J�>��a��Y�G�x��kExEB�gj\F����fU�$�J�N|TQ�?�Q.��X�j�ȝ����?�-�o�N���Q�����0D�F�Z>�Y&
�?4F�IH��i��Nڈ���w*��[���u�zU��c%0v�����Jo����!L�W�ء	��HZ�i�7��a��,l]�<O����ePk�O���p<���D�
`�Y�ɜ�v}R&K3�����E\k}jH��?U7�N� ��e4�tĪ"��nc�T�C��,�A`@h	�y��1��ʣŋ�����b`N���.��'�{�b!�3śW�73O1UՔ[ ~�޻����5)��i��DJ������uo,�)B��"w"��2�=�'}��R&Y���M�U���٠�$�I���P���uUj�G$���Y�[����'a�.��O����e걂�~�dͿ/�v	�ʁ�=X�����#��J+������bB]�^�y7:�D?5��'B�������7�o��̼� �W?+}�d�� $H��N���q�:�2��E�����!�t����}a�`#��ߋR��jIUP3����O�96^O�M�,���ɝ�S(D��g+����Ѯ�����#���&7A��9вEwrLV��j�3PD��Y!B�C�C������������w��{��G�Ϙ"�('���hs�}��w�w����i|��x
eb�B�7�R`MnP�@}O�7F��OG����S�De�q$d�4^<��ێu�ُ
R�O�0��ׁi?j�ⱃ��X��g�AE�;���Ϛe#�o�לJ5�=�a���s���z��:U+�p����p�-P�-T|�ȑ6��o� �Ѕ8�'3���o}M�W��l���VO9�M}�Lq��A5�h��d�}~d��L,�1V�'張�cp�x���a �ݛZf �60����n�I���b�!��7�y�R�^�D�V���F/�m�zz����/���L��yhlnq]l���vd�0�x�.��be�~U��[��X��x���$�eI��6W�T�zQՠ��q�eW��	B�b6d��}�-da7�q>���G�U`���&��L�mM�1����q����0�J�&)����%�_[�"�M��_����mOV���m0{�
X=9F�k�Cj��l��1<���[���}^�����W��W�hb�:�F�D~���S��XE>wj����3����"�C�Svr�-��&܁К�m��j��h�P"�y���P���3� �����Yr&0��<�)�շ�9�PJA".W�e��p��?���m�\�ޖH��	��\�g�.��lX2���HcS�vE@�
��g�-DkHu��e�!��͕ZF\����P�ʰy9tF��E�p�t�Ҧt���<��v����k��QN��ò�6̽�绣�I��А�=()3��BX��RP�G�F�����L�"HS.z�u~k��: ��X8̥<g�f=���t���ٻ��ǎ�/?�]����#G��,I��a�'@ʡ�ja夬3�,=��<�P��^k�d����w����{CU�%�NJ�F��Wr�"fj��6k�\|!�H�������Ā��4�h��İ8�*h��ٴ>�)�V^�!Yt4_�7�H�bӯ��w+���:9���%��Z��]^�-��"noB�l:X�$C�`�џ�T�7�V�=,�G��~�_%�����T�#�%��ĕXx�#�~��ۆp���Z�햿 �'ăm��B3I1��#�IKex��_��zw\��g6�A#�ڠ��,�ob4V�T5G���3C�^�Pİo2���>�[�Fr�����íJ�����N N%����t��y�2���)$lu�	N�5�_�'r@�e%j�����3=�Mٗ�z�S���n{��Ћ�-�<X�����!�p���v	[o	���n�m����� dz.�~�d�B���n�A�n���b!����Fd��s4�r��D�a�`mL���R�m�+�������~����}���n��=_���Loz3����	�l�>F
��NO��	%1�@Lj}�j�2�x�&L?��;�Wp��	,���Ky����ظ[9'Y�v�37&�Q�vI�����bg���uJU�؎���r�Hj땮+%����ߘ͗�UK
!嚬��		-��OL�+����R�9^	1ӿ���Uz�YWK�s�H�%+	&P��h��tk��N#�9�ր*�]���0��I�Ax:s���)M� 8<")>fy���J*s~�P�U�f0(��.F��e3�~��H�(�;#� �����r��K#��w���6�1�t5$�4bS�����&{�dq_{��;Կ:�P#�3�����D}�6�!����k��ti�l'M^Ȫ�d	zѥ����L;�^K�vB4�$��3�
��E��Os�����fJ[����	Xu��S*	Y-v��]C�vȤ���i �f���S0�o�S�pyA��e͹��wu�m�9|�QW�p��N����g�٢���!��<�����}�#$2R�.����B�
�-�C��C��`_�R���C������H�2I��n�;2�?��sr�0��0��	Q֧�)x���Z��H�4�v񦮆@��ď-�X>�:R88����5N�b�4�BE?�CI�t<��Ի�����=
L�U�ޏTԹwd����H��G�#k��B����/� j�+H�Z��V��6G��xu��5�:�o��*�ّ��"�*.(�Ԃޏ�6+��T-�	B`y�RG��d�|�O��~��~�<�C��I���к��l�*U�R��6��J�q�D���Q�)�]�����<�~%	���y��#XL���p��`]g�͖g2Zv!�l��w���]C^7���b|z+�j}qg�r>-iP���l�F$U����h�wʼ$*3O�e���7�Cx�70_�B�R@����_�ĪAP�$5�u�q�_n�d^Q�+���.YA�7\�'�U�	Y���v�c�Z�K���ݩZE�#�P)�ු42��������,#�]��*ޥ���7 .Q��PG��w�r�h�hT�j1�aTN�5آ.�^��	��m2%2q*ow:`���Εޑf�j���!��"�U;��T��G����1p����^�G9�5�����'��eUQ�[����Ң2�>�,����<j'!��5�	��<��:$��2}�=:��Z�[�Y�N���\/��x�1�M>N�U�ϩ4��]�2�]�w|o�L�"Ȱ�+s�7�_��^)X��C�� �o����`s������k��]�M�����/Htt(Dy�8�{T��
`k���0,H��SJ�s.��)�o�A�7N�;�{��Z�-� IO#���b��(waM�92̳b�a��D�߻��xW*����C���$ہ�R��.C�-������1q�d�k~}U�h!���+��0w��AV"�~q¼����� 4��<pmPA�U�����K=�ef(�L.:������� hu;$��b�=�q���	T�>�T���<��@H+�=E3�x��'�$�$Wc*�N0�ي2���)�K,&.�;�ZWf���$wl35��ۈ��i�$J��8z%q d����j���Z��$�7V~5�M��]�s�:���Iْ�%0(�U9�p���
i����Ɩ��9����'���d�t�X��~8���=H��9?���e�>*%�$w6qN�W��$�>ps�>e�ȵ��W�	�,��>�]�_HT���8�ka����g1�ս�2Q�H�"�n;3�73��]qj�u��0���	�>�\o%��:�=3Q�!�q���
c��
���(����5*TD����k�x�2}b�D����i��o������]O��:��Vjo����~+Ne��՗�8��c����XPQ{�ѡy$�ӣ�������n)��u� �%I��]�����)�!������Z,��_����υY��]�H� .�z@�79 )qԚ�b�m�RK
�[Bs������߃~���<�A�#�^`;?���[WO(.������.�/�@OH��Z�7�b��8E�����Pq���G8����7�{�|	�[=_�81�s�aμ�HL�@��$^���Ͷ-����X\�p#�-\EO��3��2�I]E���7�V��o�s}�4ʧH�MJ�^П��Yk�0��5mNǺѪ��}���_Y3�''�LK�LvA"8A�Z/�\F�7��Hz���	�F0~3�q�B��Z�L�J��� 4g���?����*]��h�x��V�^�8SP�F�9�"�u�U\)� �`=���~��J4Ȧ�N8s��Hx ����Qw�k�j=��Z)����Yē�V��ܩ�:~��vN���RT�K��C]�8�]�*��H>�tu��2j^Û��IN���D8[щÚ��^��27u�Q�k@�]Ͽ[$LhLK�)�T�,���^��� W	�B���q�)nD�&�ך�:sE3�*@969-��=Z0�v��� ��~�7�l���׻�u;��48㶶"S�-�+�����|����ۖ,�hk�����t]���~��nv@y"W��I��N��o���s3����F��W]`(}N��c����O��G|Iv�z�yM"T���橢?Gfk���xV\_�1g-�P�pز��O�\�[�N�憦��}�-������~��{'�쳋��;$	�s�E�r�2�����I�s���({3��Q��iD�0���,(qqV����N�k�����'�ѬK�%;�^�*uD��HM���g���u@��5���b�Ph�^L��Ş,˲Gϵ�-�D���ί��/����)1�����H�ƶZw��V���\�hn��R��ms˜����c�U)F'��1� �q;F�r,�'�z��u��1R?I���V�C_9�Y�/��8Ex������
��t�L*v��GIg@I:J�+a�yd�y���U�l��ݵ6"�\^��i՘�;[���l2cU�=��S�΋FX|#N3�]Bv И�^�sYv��Q����ͽ��U��l�2;�}w|�b`��3!ĵ#H�M����͟����2��Q>�l����#�T��[5pp�=+$��f���p�fAC�����HWf/����7��ڥt��E�\'!�n�[��;S�۳L7�0b�f:�wQ���-ZI�/��_t{"���w��P��#;��Vk����"���a~�|A�7�d����=�� =�ο����;j�L%pS������A�֑[~���3U�ض����M�@H�~HRq�=/�V2*Mc�'j����炚�!#s������.][��gm��WME?N�-U0.�M�ɲ�5�6��"E&��nΙ�|�N*�2��8��R3�c���cK�t)پ�ce��p]��]�;$����&aY��`�]>���Y�\�����:�m�A$�SI
�6I���d����rsY�$�.#|�Ʉ��x!��lF����W�m��c���l[>��x;{Т���Y�4|k��
����~��o�&�h�n�xz�k_�O �'��AwN�Re��.k��8-/A�c1�����>o=�K�_r�W���wH�vJ��
�U8����$������S�)��r#�E}�5��5�~^�l�td����n�B�|�KO�	��[��%�53�u������6کcsr�&v�G�~�UhX�����yu���H�����1������y^�w�5����*�D=B,�0�����'>��jy��CV��9���l��1��ZQ�أlӟ���ۯv���7�4�7q۹l�V����P~X�6�-����V�x�'��&�����:*��rY��Y�czZ��H�w�:�t�Jo�3 躇�(�%;@>�p��:�%�BM�ۨ�m�;(�vԨ`%�c`�����B�ͦ1��MK�cQ��q{��?��m-�������M)�	B�_���D�З�vmz�B�u@=�}�6A��>t�m�m�Y� �\\3��p�Z�KjQ����gJ�K\Cnǔx
��"/Mj������˔����>x:誏�(DxUW�/�b�1p�,|W��Q�BYWw�x1��&�iR'�\�"*�����U�j8
�w�rF�$'CH7�b�ɖ���Rê�&C{b/�`��N�RV�,��\Iח8JMS˚}L<dm�����y�+X��~+0"x��廱��j�|�-�3��s���?����6t�h�ĸ��FӴu�s�o�>,ܒ�'�6��ӊ�$�d���7̺'�c��@�1�E��P����i��M�Y )�z�A�|�,�r�cT&����sPI"K��R���Zԅ#�(��R�q�PJ=����[_Sc�+	D�j��xx�=cZд��#ZK@�%�V<��J�b����!�����xe��
���ǧx�MF��Ñ1r�iuhѮi�[f{T���PO�VGqԌi��8!t�i�;۳�$-a%�c��WgAfn֩ՄB�H��:N���g�x�A�P'#a8�_��g��W;�����"�S�~x���}�-'�o���v�~��gsM�AI��
��/�sr<���i��8��׸�V�B 0������}��O��Z�Q�:X�:S뫳�� 7͟G���6���ލ#�ۢ^���2?uד }�+�n��S�iL��x�d��Ү�n�U}�,��ߥI]&�Ş�XF9+Ps]k���Y?#��a�(��ҋZZj��凩Μ��j̊�/8�绁�'���px��g��$�����p?2P�/^�d�-�!���]��"E5�-La���*|�4ن��O6���q5�W#���>�6%uC�іV�h�׷�u�O����c3�w����t;��[����o��Td�s���C���b���pv�ۛ_�;Q�㋄i%�ȳ`�Y,a.�51;Vn� ��2.	��� �E�ǂ��S'!�u�V^6j�8���?o�����%�.�t�T��A)2����YE��x�7���L�1�8�	������wm����g0�>�1����X�#�^�S�"N��m�T;&��ϕ�5�R��-�Um����4�Q�%�\��e�,!L�! � �n�Y �K�Bԋr�Y�f������_`T��9�
��=�}Vu�JU4�l�-�$�L��F� �Au�y�bD���qJ�FF]a��I�c��ط�`���<�'��i��=��<Ŷ���E"��Ѿ�R7��O�e���ށYכ>��U%��p|����U~��a���@R��LY��CHO��+���p�Z���qq�H�}6cw
�Jbd��˶RPO�iD���g�����V���Y)J�|�5l�+��+�X;s=m��K3�-~�~�D�f˵D4��3H</L���l���U�ڦ����`��)ud��@���STJ���YWj;���^��C�lȁm;8�6���\fyߥkp���l*>9�c��e�h��_ �+����d�(h�����%Q}L�E����}�A�],]de.ƌt�"�͛QD\ĽЁ\
ּ��*���)��_�;MA��:H�g���h�����@򯏄@Ix|]�K�Rһ���Fɇ����TB�@N��P�\+09��-��<]�j(Md��=ci��8�d�L ;oh�#�J�6ۧ&��ʆ��9^9)Λ �֍�]T��NqXyG���#;�R��5��:aL��~-|%?d�u)D��ȭ�76|�>dA��PD���aEʤ���eJrªY�C# A˙�4J�lm���y�ey�T`a�A��<������R�;��.c��&~�ChzF����x{xȩl<��nk\�}"o�`�5�(.稈�bg`��et�{-����+�o��Eh���~���)w�L��)�yj�G������ 3��ʨ(�#L0�B�A����S�4�v �c�Z�E�#ρ?�3�XI˹N�pi�����e��=`�����2!�V:�#�g�/�r����}���X�8x�xK����~ �!��*�E�trx��d�l�
Aۨ\[�/����O��D6����1*̦�_%���
ڍ�}>R�:D�<yY�k�,�ĸI����~�ɏn!��7��%P�2�_��	��Y���~����;8CU4��`��\s�*]���>;��XZ���\���*�+"�}�Oe,��K�R�^�����������������;8 :#�Y�tsi���hN�r|�� ������^a��qX���t��[�6f9jGF�{W;�C�Mti���}B�n��.m���z���ʼ���Z\�m��ۦ��
���ժO9�f�y�]�ri��KraBy �$_Ij|�=�)�;�i
M��
P4��t.�A!j���;�Ss�`��1����1X%j|�������ȼ������Q�~��1݌�ӕX���+�"T�����i���P���ʠ�����~
j�.�T�m������і��n�.���ۓ���������V��2y]U�k�e�3Q&���=���U{��ߝ6	�߰��aJD\d�&�m]�c����4(��ڤR���ӧ�/�g�Z��c3�ߤr3�uh���#��'�A��)`���~+����m|��ӔF�C��k��J0���X��l�x!�'& s�d�إ�8)�z[!ŵ��^P��
�~is�J�O�R�4��5��n/�����_��C��7K�`5��O��Y�_���%+#�ng��b�֟-�QQ�J�,�\E������Y?��-�'���[&,�So$�ذ��C�A��J��]�a"r�>zB�r��S�/ԍN9Ӯ��p�5��J�w��fG��&�|�̌�����$�>�<O���~��o{���1�|�h�_~�)*��I�<�iM�%�E�F�����ջa�^}E�-;:��R%'�>A�ɟe�|Y��z�P��n�܌�6���*m�sn{����\6:�V�B˻�f�nRr����ŝ�(=�9�(Y(Ǡ��$���RT���2�������tb�4�c��$zb�])x�<=.� 2GP�'#^4�DOU����l�����,,G׽��Jc�A���y���и$�l���R�0�ZK'�>���&��O���[&�]��POo8������N�+�}�ɝ�S�C<w��Yo�Z��s�-s�z��m�H�з�7����Q�7�B�iSl���byg���k�׆zB�rv�5�^*	��E�e/�?�)ܠ+���Rw�O���}r�9Kaµ��TU.��$\��#�L�D.�����K�\�#*���Δ��,�';.�3���q�ۃeG�2���vh�"/�~�dXCLX��,2��fb'c�W�Wy���j��G���v"���fa�b��PZ���d!oW���?�b)��I��H]��r�*'�>�bޥ��8J��jO�CHATQ}+|7�8bٗ��˻�T�oΘ�O�F��8���)��h@3�B]�{d7��ɼ���$� ���)e�
���$kL^�Ք��#�I��v �Fӆ�<����ݮB6�x�P�}�3o>�8��1�ō���V�_��;�r�Q�I�BZ�]{_�J�V �rK�Ҕ?����N���-�\�QT>>=���B;�eQF��X00J��6(����z|�o��g���i�'qDu\%�J<ٍ�Qp���)��.����h��5|[��y3aw����ʚG�`b�6&U�B,�{���_�R��'ŭ���Mƀ{5��0t��D3c�5�씢���r�:_v)i��)��>�m���`ㇸh~�G�������:�~��G�X�O.��4Du_sc�Z��P:T���Vz6C�;6����7�ގ��ꉺ��[��l۠x]Z1�p˵�1���y�*;�Svf,��57�@H	��g_JAp}PI7G��k��=ם8�U�a���ɹ%9�N(E��	�,~/&O���505��m��2�*�O��2a
1�&��rW�veI��
3��AJ����S��0E����+�C�^����~<<�5s�&�\D�A���w֐��d��o�	�K.�H}+�O�ʂo�j6�¨i�����w�k-�nl�u�A�|�C�g�R�[>���<����0��q�M��vƭpno�}Lbl�mUT<�%���uߜ�Eυ� ���0��9��4-�ɿ�-L팩0=����ݝ���0.w��#���ˠ�J�!��$�{�pIX7�r�˔�/�;�Z)�������H��`{ g��A�o����sS;Q�D���P�@[�(ٝʬ�ō����mØ�3��l̓���B���AH�lB������>��"!&j"��PO�Y��wj���f�12T�<L�~	�x=���h����^K�+=G�����H����A/W�P�sof�_��ӻ� ��.Z\I����	M��e��He�iQ]'�En�_}����M����i\��=�p�}�b�xy�}f��6�Ʈ0��+\�G�%�� ��E��h��_����o,�@kQJ�B�&�x�+���b���gs�N��2�+u�ࠌNv�շ�H��\֖�N�M!|d��Y��u�̊�qQ�M�y�e���d�}�r���m�]?ۋ�sq�z�*��V�Y�D��
e6������e[C\���M�V���덭���N�R�`X>�Sf��>��jN�^t�Ҙ��WaB��3۩��aAR2���t���{l���T�wۧ��b`Zs�~4��̤�`�]�����e��i��U���[1&嗶o��DR�-�%�E��cgx�7
T�.BsW�+�k`S0U!�l*qդR����o3|!��/��(��*��J�1D�Қ�Ж{��[��-��>�o8��v+��ÏY6�.\���A[]�7[�`�j���g�kd��p(r��
��ئ_���K�#�qU���=l�!�����4�[��n�С�Q0!˳�+	xIE���R�E�>��n�+wnQ[���A�ݓ5Q�K���Ă�-�? ��K���Va�ȇ"V������Wt� J]n1����(��CL�Ɩ|�Έ?�37Af��YE�~�d�l�>�;ǀ>#^��uY�����V�`D��P.	D5�h,`�z'�Ӥ��O����Z� ;�>���2���p����>��Da0��/99t`ں2v"�[w���|�y�I��$aE�a�m�ӂ�^�ŉ��3�{���(�O��?���~�B��.�+'��m�˓g���~��N�鍩���U�.����TA���j"�Ӧ;������O��u�*��\�W}SC��F2n�N����Tr��K{2�(��߹Z{!ƭ���h�|���������%u�3�V��S�H���������H�G�Yl-Rӡ��1g���s쌤b�`����ۺ�Ԡ�'�����]��oE�\׶�ֵ�M,_����c�Tyŝ���V����gT�{<q���N���A�'U���ā����Y���Be���ؠ۪ �L��c�*�)��i�M=���G�w).�j��!kfK|2a(pk�gEe?�!�d��\:@U�P2A3W2i	�w����g�Μ�Xow���fKu0��n	��W+M�(	20�#Oܽ{0�"���6F��h�1�e�<2�mj��Tkܹ� <]�^�m1�gPڥh&�$�qOhxk���#Ȉ��in���4�X֎��?GT�s�몔�KN�L�)��,������b^�~ZÔ?�^h�G�)�;hD�[�Qe�m�?���(�λ�ar��)@=���]�s��^a�U��6I|��y��ne��<��]�N䲵�!�
}�X�-0�ɚ-"��{\�.
N!ܚJG��p�S6�B�{��WOMo��k��XX|r��ɡb�z	��zc2��0@�QR�;h���įQZ�M�[��o����j��,��з����+���ڤq�ZR��������3��+�`Z�����lr���`w>�S�q ��4l���Rb�r	�΅�r~3>sU��ja������^kd�[��E}�+*�͖���c[!l<�j�{G���r�!�֚�/�9��J�_Ϣ6X ��R`�N~<�=j����w`��~�S
_�[��w��R�o�G�ڜ�lPx��>A�q�@��=�4e��w�F��̀x��������\ �2���%*��<�$�no�x&A��ak������D����w�(��ʀ�	�A��w�SHV�������^˲ύm-�O��\���Ơ��V��P��di���,j�մ�(e��gC�z���T�5�2�4�*N`�1���'W����jz�%=8�2<I���E�r�!O[�0n��6�J{ש͐�)	��Z:�e�]ǆ+�0a������P���3|I��a��'�-��U��g��l#�Q�	_�~j�&?��{n���0��F��CW���F��Q�@S'�o��=�:�S�롨�cJ#@�p�fY(����E�x��U"ꢫ�ķd�������m�wa�Y�u y+�Q�$�[�	����M'�q�F_����B�Iˤ�(En?�C�{1zl&��3N_�V@���jk�����QZ
�zLŎ�h<��1�����F��h�~����ou�g�����э�H�>���/�?:�6�
�;�{��æ�!���<)�U�����Y򕂰����1�^;�~��on@��i�Z�ڔ)K�)��* ���.�D�.�<)�a(]��NT� ?��ڃ��e�y����P�y����s�`�����8%�R�A�0�>�*� �,E.}3�������ڒ�i�fj�_�cX�o%z:�G�ox���=�������V��o_c�m�E���	{��,}�������2}p�jҵ'�·�{GT�_��Bx���-��6���t�[�Ȧ��⌐�u�]�)���
v&�5�S���Y��J޻��kq7lvO��Î�����mli ������0#��b�km����3ܚ�ChuTB~�	;�~p���B��/���ᙢ~~�ZJ2�ⷉ��_(��/�.�_ܱ�4���Cq�a��;MМ��c�5g�!���f<��;�t�=��Ԭb%>5����ZM�<(��W���"���&�6���*LC��'>����������	��SE��4������θ�1���׽����IY���覰\C�O�!�K���_� �u���ՂZP3z-x�N[��-�_÷�U-Aab����p���{O���4�~g����/>?�k��^��@��~��w��6�P���@,t):'�a��2��[=��/�<,��ҏ�Nr�OPMe�m��e���OBZ�4xpg�(r����E3kXi�'���O
b �ƻ3��5u�ߝ�	AGUL[2�ￒ�1��3����鈮d�!�Ȉ�P>i{1ZxűG?�+ۙ�_[l\b���R���5�%ft��Kɚ�M�i�\KtIQw�6~	9a#`q
�$
7�~�8������c_B��Le+����v(��4=4]S���N\Bx:�]h��D#]f�%��T�5g�Y�t>ߣ�ZJ�F�i����}=�O��؞����c:�p�Xb�x
\�wR��N���1.
.���+Y_9FgK���Ƶ_��|�WfH	�V�Cn�ωn
'��~��B0�6�y�E#�����l���8Vҟ�1ws�7����/)��x~"�<�]��rҜ��ZAvg\z�o���LuBEI'�3c�#���3Jd���Om�0�ik��$W�7'9~
���f��{(#���t�	���Dk�1D�*M�=|�n�O��9W��|$p�ηSS���]��
EM�� �c�C�!%�O��������w*l�J|V��"�KR�`�;b8�Bc{g�z�CM�U�/�y5�Ef
�=<	G�n�h��Aǅ{!=h�]��8��10&z�^�+�T�Tv�Q��^�"�Q��D����K2�2<n��"B�=��y%���6G�����_v8�i3�?�Q6=�I�]]����{w��%e����+�h�ʗ���71��]E��������E�<��)��n�=�P�A׉��I�Y6�2}+���ǢD�*&t�yR�A�b`��O��.>�8�O�"
������G��;���V����q+�9��&����*�&X�,�(A�N��[�J@��4�x�����s`u�>BQJ�
�u/�$?�>��9��]7c�"^��Z[Z.�%p�a�h=���Z^��jG�q�t:��pUf4�,>�.E�ᬫ9�ym��z(V�?7�S�p�y�^��cl�Pl�к�Fa�ґ�������A�0��W�0e���V����}aiO���J8:��n"I�kK
��������C��@`��e��7[��Q���y��Z�&T�x'��=�$�,��Fò�7�j���ʐ��}�;yVΡ'�9�,����8����֑$������;�mx��W�Tf<�Jӯ�Z�M�>u���#[brVS��,֨f�A�� #��>�g���=4��.Q�"���j��JUߙjy���;���FK� �D��C�n�v <�G�tf{"z����㘓%e��+�=��8-�������&�U5A�e�^��_���\���Vø�)�?���gRՎ~����)c�(��j���|;���w1C1D�\�,�\
��� E�c�j�%��_��߶9�����}�J&R�C��&�Y|�5d8`Q�zX9�n����I2�۪G)~��]�n�8�dɋ�s�R�ɔ��Q��[+/ai�T��e���%�r���U�S��@|L�#�w?����b Cx�Brݪ`'����?;������]zpO>���@��BPn����aÇ� F-/�l�.#:��ϸ2��z
�u-��_aj�+;�3=��#[�.�IB��t���T��{��_ʩ����[����.����@���)A���;�o�r�!
�l�ɛi�Ku
P�Ȧ	k���]zw�fo�<��.܈~��r��tq��ܙ�����c�ñ=�Lq6�ac���<���a3K�<�������F��e�	����_�u0?O���~ ��w�$'��*���l�H!Y2�}^�2K���%��BBȏ߶�J�~.V���v;b!�c�=%DT4S�OD���)P q��1a\�G� {��*=/Jë5�Q�X�^Ԭ{����)r�R����d]�$V7}�@�"���<�n���>����뒎���@�U��t�q�~a*01�=@N,�IH+���]Y��8�����E�e��뺞s'�U��d��.j~������:bh (�?��4��8�OR�Zmj��=��<9J�fݔ��T���XN��� 2�|&7.�-�ܮWɛV
�)Sj�C=�����	��f&���+(�����<(e�Mң�n�p��V���EgBYcW��?�N�h����>�q-�t4��c�#�������;D�1��/�/䶶|Z@�StU��p�'Q��Kx=�<�&�����I��ΔNk��32��b��糭��rx4�`{�g���A�*he���ݟ#����~�v��~ƭ��(�`lp��S9�ӧœ�Y��#���SL�z�?#����M�c����▁8N�#��g��v�����_0؄�`0u��$t���L���n�6��WTD�t=�~��L����
I��u�b�<�燮`�"�����!���)(��'�hVkU����X��w���9ˏ���$mf[��۸�!�-"�^-[-CTl�4s��U>��GȉL��(g�EAy<����~ڱ��5�	6�f�/?_Pؽ�����dٸ��Ãx��l�G�g@�GS�o��*c2Ͻ���o-�i�Mk�-�&�H����7w��g9M�S¨k f�(�\ȸ���>	��f��=Fi������c��m�m"Ɖ�8��76E��1�'=&a}��j���\�%ޫ��L>�aq�V+�&�*/��ۚu,���R�����QNz���m-�C�,���͘�gt�KW&&[7X�*(���`��g�H�`/Y��4��e0О>��K�����ټ��n��J'1!56E L���=��u0�SqϽ�
��@�o�4I0t͏�m����	���e���5Pϗ�\�<@�W���}Sy�sFp,�i�g��$�1.�t������} ]dm�1�~
�wuo�[6/)�<m������ƃ5�Z6��\�Ε�;.�7먨^���Kچ
�Q�o\@�D[J0��"*���"[|�^V؎�@�1_��'��f�ʙ]��l^dA+LHk��E8x;�>D���׃����
y=Hos�s��ˬ�X֎g�D=7̪�v�ø�P��O5�;�U���p�;A���ɏ�)^@�ᓗ1�u�^P������$��~p�x��K�:^�2���������s,��[�%s/x�NZg�QE�.��U2D�m�Qp{ '+{����۴4���®R��+ �*��*$��v��A%B�Yz���_c2Vx�9�3Y�8�P��~х'��B��m��PZ$�����<p��CH���c�[���y ��h����'2,��\z�!��S-M��H���n4�%�M���+��$�������AGD5��K���KN,}�*�&��_l�,v����Z���?�l��I-^E�`W�xd&��{��l�+z��uГ�GA�
��X��@�7-��42�8����6h`LV��m@��6���r�� G�:���萭7*��J4��|@��;B2��n�[2�X�8���#J��F-F���dQ�@$QLo�WY�ɹ��d@|��������� �,U�����D�gib)��J?+°�b�^s@lq���Ii� �@�h.�3��KE댯�O�Y�1����|��ȏ�b�]��̓'�G���5XU��.���$ƆQ��)�F̤��s�6c�� �rn!.��[�`��a�VS}�Gy�IW�d?��YD�Wu�:���J���0�#n��K���ʮ1��uP��_N�buK��sD�̭.Wn��G�����2�))���N��\�/`-�_W�n&�]��_,��3��궅��u�����Rt�iu��\b&/�g���E��ɂ�IM���Q������s Fݟ�d�h��J�\4{^�@G:G�1� ?m���㰊�"�~����.<��^�=L��r��-|�G���-(yt��p'���3VulD����Y��U3T�z�ZG�Bdd��)�N]
���h�^�13yH@=�TPk�7ً�m0�tY�tGTٜ8�C�?ܶ�����`v[��!�+�IV�si!��䪩� �D5��^ �S,�Y��zC����(�a�bW���,ن�Q�AT�������]f-1�]�1!5���%,���8�z�p �ۘ�<Z������QN���������o����``Uv��$wR�-�:Q���P������[OI��3WU���%V�J���O���yO�����y�^�ۑa�%�;@o>X�໳[��z�+���2[�""S�8Dw�F��΄P�+�LEg����ţ
Vr��4ӓ �8����T�<mp}c�[�ۋ��0$���i4�bf��~���Y@�6����Y�T9������pwf���B��Z�s�,�
��b� Ơy}0i<VE��x|W�`C��0�k��\$5M��k����")�9���R�K�f�<��I�VY�C�P��]��*#/���PI=c]�
�����Q�d�����m��h��0X�I�c��Kګ#��xDO�wz�9�EĢvNe�'?���	�o�2�V����\
�4힇\����K��e��I�_�M�j��� 9��z��w�++�8�����W��z+,�X;�rV�����F�C�eX�{�3`$Nb�N�-6����~�KӄDbW�4��ui��TGu��e�F�,�s�2 �ܼ��g�a.\`q%R�[��õ�S��x� ��=�����=l���t�m��琑q�믜�!o���XS;Oz:R?
@�v1���q��*��[jՈ`��;On�gl�n�w[{%s�ް4����y�0i�	��>�r�.�t�@x+��ߧ�ӏY.�FB�Î�n�O
�9��D�f�QP�u^p|D��|#���­��kj��<4�9�NX5hU8��Dq�[2ݠ���~�#���~H���@߁m'긌��<"҉ ��UɄ/�Sɠ)��W�(sg��3�Eh���/`=�uG8ǭ��qw�] 8`� 4��;S��)��\)+J���:�ƛ�i��Lc�51�x�x���k�Hr���FS T�6�I��I�FOR�6�%i�u㨋��B�0�-����Yi0��c�Hy��/��3N|;Dv?���B J"�o�CسCX%Ԅ	����v�s��Y�����i�0wN��A��������?��b�h�i�+�3��QH�z
@�](�9��[����}�8��꾉3�b8^?ygzy������6�>�Y�P~����&��@W�����+E���4r�+��Km�Q�HJ�����~Zv���r(�.TH���@$+w����aI�3)��9;A�㯧'j���B��j��<Y|W��\��]:9��I��!��(Y	��G�&��/ڹ�I�if��6RQ�%�	r��ъ�=
Z�ہ)1�hx��䴧�t&�c��F{z(�n�h-k���hR	V�7ԯR!�u\�z�08O��V���T�*}�.!��	DFe�hd��9�v��}/�}�y�E@��r�V�KZ3N/����EI���~pT�>q=�m�j���Jj���X>��X�T�I��5}w��J�Qع�4cDW�'��`Z���bF��,T�4׼���h�1��`�L\#����A˽U��3.�&�Ʃ���t�h=R曬�������]��t{��M����l2���ܬ���+&h�b��C�H4�E�4.��c*-���Dt�$�2�?��N!��iT-I)���:Zeܦ����W��Q�.�඲, Tb��بs	���.�D�A���cv�M��� J�����Ǌ]�F���)���É&~�ؚ�x��
�Y�T
�����uX���=N vC� ����0�-Y����ۍ���bo(mğ]>�������'�F�s8�6:HG�\V�+1b�F�߳�K:��T:�?��vY/�DܾW��bv⧇%�>�1:>8#�?"�z�f�)��[>��|�qKL�&3�g�Կ� �˓T.��!��h��M��s~��soq_$~*�s������*/:*˛HS��+�!\�L�Q��I���ͼZ-��E��4 ��EP�d����A���">	#6�i�ܥ�A61��Ż*Ϟ�P{]+��R$��{�mÜn���E$���vA�Y"Wٱ��g�S{��n���
xU2Ru��˽�˭��Z��0G�L��,f3;l$�V)n�>�>�F����̥������l#�JW���XIS�"�Q50�@w����Qo�]�pFU�مsb���� "�,��<�L�����YK�k�u���K��F ��k��~]��E>D䀃$�YRÒ��M�5jG\��_-�<��5|n�/�:cl҆�.sk2Av��p�A%�[�jX�EY/c������t��]�s�@70���A{�(�#��N:+.ܐVZ�Bi��jd�����K���E����m��[��@��$�'q��id�o�f?$�x��a��#~�nH��w��s��h�Zi�d�A �O��L�����/G��xr��b��T�����^������i�GY�k� ���s�.Δ9M�r}�a��U����8-�Shϻ����n_̹�c�a+�5U�˝Q6o<��CƛB2�<l�Y,��Nj�r(#Or��7,+��xm�~W�c��=U7EqE'���!D��4�=��+��|���'�ש�B���a�V/2�Rg���F,���ת~u �+w#3�$|�Y"v��ݐ�.�Dư�����w
��"ks.��~���s�-�=���za����+�V@�������m@�&��dYJ��J��<i3=�qf�[wШ��������g��辠4�g���NVț*l�b�����6bc��8=��3u��a��ċ('k���K�]I^N��f6��`�M���?Q�i���ԙA��0��]Ok�
�飂�lkû�}��^�@��/�ΐ<���'1)���	��g����-?+��+�)�A�G*RDJG*��Q�"	o�'n��2Lm�ʰ��W��{���^=����\����'��&Jh��U��EjR�nڅxiT������5���Dն�a�`$Oc%2�K�*4N=+�f���L�����,v����7��s>L�9.@U���B���RM�,���T��I���8�uu��
b�34Lc�&�֢�R��ex�/�.S����6; �L`��u�
�J��<��Hkv2O���ң�ZX�C���� f��X�lo�D�����`A���`��s�4��|����AIY��_�W�ojg\"E�g�lO'�o�=��)q���/�2�5:�fv��_~��h2j�M��=L�7����뱍�����"��K둌c\�Bʼ�{�t
{��djZ8G̤��.�Ψnm��_�������Æ����&@��q��,$���㹭�N5(��(J��OZ�\��`9g������܃�؊$�-o$N�f9���[�z��,�zNb��ɻ��q�{ �C�
/�@��׷�(~�.�A�������XU	@��	PDIp����}�@��Z�w�
����<J{k�� �����2udA�M{>�ߚsP�.����*b�/fEuW��1xs�I�7?+��y�>[���hq���Q"�l�����&��`���})>l����EG���
q�sL��\��)�q4�
Ğ���-Vy���)������^��Y���`��C��,\+��������'�d�D����X���(AB��~;�b�M ��M }.�79쑩��L[�}��l�VZ|��?���wEA,��n�wx.��ﭥa��p�m(������ {��͍e�j�;n����<�Q�G8�s���NpCOv-�D�.�̩? �v�.���.�=7@LDX6�&��n��<�~��[%M����+�?C�����#D,KSP�p�l�C�T��?��ſ�Hm'�e����{C�緳����3�I�ir��@���gn�3��l���B�4:h-���t��Ӆ��b>�KŮoX@.�],��c�V"M�Py\�Oh'>Vb�/Ih��a\6qCeп�����_�So&2��r_�}w|�N�bs��ފ�i�ßOu�z!�i�!�Ju����"cpB�&v���^�c�nAx0�$�+E�e��^�P1���e������Mo���1�Q0�a��^�}�88H8am�܆�P����ZQ�˃b4��I��g�֥B�T��u+"v��eL)���ч
)H�%}�Pr=���k@S|Ѽ�=�r`D��fD�A]@1���z����o[�i�(o�my��i��>����L�>RF�7Z�HYc9��Q� �]>@@�"����Z����F���2)��:A߿wѱ��h%굤�{����B��,a�e/D 0	u�G!���o	�B�O��g�$�Qr�z��tYcUށ��P�âEپCs�B{��x@h.���P�:���Ѫ�2Ӌ����^���;Y�����Zc�<sT{n������
�w�A�բZT����SO���\��Qw^J������s��+5S��ͽn�����6�c!��<��dB� z�������K���2�z�#��-F�����?�RQ��j�W`���| h<� h��o��9SKE�������Keg�_lVh�*v�tQĴ"/F��6ޔ���G� ?��v^�q?U�ڊ�y%ME�ߪ�4�_~�	��@p%`ܸ��,�:$��c�x�ۑp��c�d~"�i��x��*T|�����m]��L��˕*Qɳ�m�E��NVq׷�vԇ������Yz*	L���\�%����?�Z���*z���vY����ޘ���5���_ ������xK�����_�0��:}"�I��Z�l�v?Ðw�5�Mw��V����CML�T-���!jb  QW�3��9��Ռ�Z���������	^C#6��l�!�㧯��r�	f�� Cb��B�6�=L��g'�sh��e�FA]?�4vNt\�M
�:��E��h��������!\�䅀I�#��x�� |�gB��r��+Cs��@h�f_����D�k4��w�j�B6+�*�e�O���}
i�(k�1L�__����cx�b���!�G��8��_�!���V��Y�fo� \�ͥ&;�9�"H"�Ms� ���+�M��ⲉf��I�o {�{u���9#�@�~�O,�(����BX?�/�o)~ڬI���;��-�s���ޙ�=y�7|�0�oƯ4��\y�Y{~Q��9���G Nozx��:s�S2�xY�,�|M;�B�<�k���c�e��K��N�lm����*�[@��K�GF�`���e/��)^�٪�c��������~踎��E���L�H�Z1o& lI�������W��7�n���w��/�!�{i�� yo�}m��]�5��}9�	�6͞\�n>SQ����6H���=g*�M!a4z>��"���Mh��-���3�MF�	�S�躔@�"�!Gdsv�"=",�8��.�����G����,Ux@��T7��/�R�La����nl�k��Ƴ����M�������I�>(�JF?Lef��y��M��s�h��">`��7<�ֳn�_��D҉)�hukQrnK�"`���ŅJ?7ق����E�#�A�����Xj�J9q/8�?x6�g�c�\M�Cao����}$�����g�q�{���`��[��� G�(#@&���u'6{��?Nҹՠ���Х��02��l�6��v�t��gh���2��8��M�\�����3�E�3�l^YÚ�?�Q�5BL��O�\��lH�l���9=D6|�r���O$�&Ku��)˒n������6�����n�j�fTWj
���	�LpX��NR`�.�`u:|g�����,9B�(�>��a�ZM ��O�ܳdn�����ō��9p~V�NQ�� ��������3�������Gd���"��Q�O�P��OPt����+��}��%�̓s?����<��om�x�|Rl���e����Ua�c�AmC�U����N��ŤR�ʷ8� `u��pYE>3n���ODS0��n�U�b���L���A�O��l��l��7�h����"�[L*	��H�^#Uh&j�}�����m�j�ͳj��+����?�N�[�v�����ek|p��}�����[66�XQ��ĞYc�d1�!�9�Yd�ֶ3�$�|S��iXM��Tz��<�3�q���M�����j(W��
e����X<������!�����{P
b�t��tNIJH�D�:O6�R�Ph!7�ԤGW��Y�GF��5W����~V��'So5/u�"(�&Z	!f��7�ƒ����.��b��M̂�����P��&�Z(И3�GJb
��H����&�X�����.>�؂ś~��"9�բ_ ��$୏�5|��-/}���Ȇ���<��õ�T�^G�A7��_ٖ͵/;�2E��m��X������݄�@¢�ݹ�TЕ�����Kes,WJko����	W��T���m��S���L��?��Z�6�{˸#�E��t�*�Ť��Nf�e0a깵�G'и��ނ�@��^��|���u.���A�AX9��iE����ˁV3}��Q�9�%@p���M�S��&�W�Y�-3 ��G�N]��wk��M������c%�fzAr�t� 7�� ��@�y(���q[g��w>�x��!� �u�u��T����q쑆�����2vH.	��|��`e^�!P����z-��en�j�"d#��P$D��̨ lpD�5 ]$��| �o�hxe��X����P�Q5]bH�`�9��c�x���v�D�@��BMb!C7*Uo)����֖H;v�����g��P�Є@㊸�(�W7���P�����0�8�\d�����9b�sW�&�q5=���6��Y��� ����ٵxv��%LS�%@+�:r|x�j�����E�m�\w�)l�$����Φ[���n�EO��4�»�[0C�Ѵe�`� ^��0��Y�~��\m�HY�_�~1������,@�a��D�r�F�YO��V��F�Țe�ɂ� q��/�c9 
)�����O.}��4K��&��E�S�Y�4Գ��RS�v�]Pg�aP '�F���Ѥ9�����=�}�ͿJ7��H�&�ƕ(K��ߢ@��-��3�8X�iHֵ���"�����8+�2|��݈��忘���@������TZ�S��:�7W�|����p�
ȹѾ��1����#����=�!�KF�(1�)vѽN}�K��s�å����4�1�%\l���f��ln��)q������l����e�x3��%�e��켉�f��Ps�|�w�Y��6i��p��s`'d��c� $��:��kk�D>*l,$�&v �Ad��P��ɶ�?ئ�re�v�\��[�@���N�Ջfo�G`m TIT�to��<:
� Ý/�_$o�.9�D`8��`�gL�4���%mmQIq�)����YŪ��H	'��P#n̰�N�@?h�-3��ƺ�|��e��9I��5K#��^��҉l�����>f6V�C<+�{:��]��j����/��/W�.�M�|}JCu4�S�C��UtB4���W��=�<���� �(O���Wʜ>�h'�U��=�M<D�8�ҟ�Y֬�a�`��p�;��/�.��r`۝���F�~�ۨ���i�:�	�z%b�lNy�������rw�$=iw0���FU�^�pu�����3 ��ΐU���#5���Dt��E�KW��tD��y�0: q%��I��XK����,&��եr)&-�
�%��tB��9�3�vZ�z���_�~By�=��>-��r����k�)w�ǋ�����	�c�:T�S;'�;DnN�%*����8;�"1���:(�
"�P�,�`��0�,�q��Z�)V����k��M��YQ<�0�����-�gՅ�:+�D�����!��@��m
K�fU�j[7�e��2�q`��Z�.YzH'�Yyo��.��)�S�{�)<>��j�rG�N���E��
7��<���0��#�/gn#��t�<_yNKB�7+���/�$������ߦ[%�aHE���4X\(����b�*��O�>H�O6�0!]$���,F��P"��I�z4�ct��Z�t�P=�mL�ȓ}�χ�
 u��o>0x�Ǎ�cY����Z�"�;`�]4�
(�6q5���g�M����Ȃ�"栿�З���R�1�!��u�ߠ�AL�(z~���mQ��o� ��2R�\*���29%@�Δ�W���xՌ����r���So�K(u����R�&��b�6���5����1*�S������"��8F��j�9�c��J_sC?��m�	Z�����	}�s�6<��m���N?��ٵ�X����%#`�e����9Emq<��욦V�]��Ko�B��\v��OP��-�i|s ��%<>�5<Q�8UC3��x�92?n�q�>mz�oKA7XjWZ�@ѭQ��y^+F�P���I�I����[@����{s0�r`%� x�[���B��� �I��@P'R�V���`;i,��=0����SrB����3��T��xU\�UJG73��>��W�zϸ�u�tR�1�ę��g�he�����Bp׆�-��Ǻm͉2I�$�Z���as,(�T��X`q>T<s����rYK����g@~Ԩ��o�I��NF-�b?�z7N���b�����v����w�{��`@Pj��pA^��	B�57XQ��c-N��ulɉ@�ߞ��zR�}����:��j��=OK��V+�kt�Ԟ��_!Zv%� F�������zX�������EP�q�P����Z_)<N�ľ ��"-ѐg�:���*@PG0uD����k��5 �{�٬8�~�	xi>׍��Y���%����<�u�J: )��1[��?�MB��:��]M��řd���N#�$Oi'�;
��*�u�L�輙�١�d�:��^�M||�W��şĚvX�=���3��|�C	iTH!$|o��ޑ$<��$�,�&E��W��-d�J��%M��k�`��)�n��o"Ç�۵��*�t%��@N�d��r��'��S�>�R��Y@��F���������CJ�����T���xa��n����G��Zh�����s1�oFo?ˋ��P�yXV�s0z�!��e��p���-�o��1C�Av_�r���y"�DPK9����Y���=i���·I�几w����G�K���{'��g$�����:�[H�f���9X� ���_�wQ�����=k1��|��!������b��Q��=�bs�{K7�_�q�mRA��TޯQ��z@ߒ	h���,�II+����=��<e����)q�/l�*����.����xu�ʐ�7k�SY�L��;���'-��p!B���pM���=uR�hpW�,�ֹW��+���2�!�Y�|n��2k$R��;V�6X�:%Z�*�N�~č���XQmo��P��%���.~��Z�xy6��E���J�wO`�l[X1<$�!3�m_�n�r+�u(^�K����ks#�;B��O�>!2kA1�	��
7F�{����K�Q��b�T]�.�Lp@+��v��r&/���cm�PF�A��'�l�h�F�Rgͫރ�)b�����Υ��l�D=�Dã�[t���c�8��H�n�_�B���`W����wN����icN��Sc�����*:-�qo�K|�D8l;������p@��'�����f�눲CB;�:(�O������8I��|rqɂk�Ǐ&H�[�H����Ğ;j�oy���~��}�����V@2G�;܂�7M?�׊��eP����uR����P���V�k�Rt052=�~R���?�S�"�I:|`E��Ru���"����A����9
�9�����W����@B$��,����Oq��M!����h�Pl�c����!�I���='Y1�w/�^��/��r9��a�Kmq���ʯ�.��x�[#��[=�)3Z0�	pm:�5b�8(
�Y2����'�`S���D�6V/�7��I��O��}[�$�2�&�))SY����=s��x�L٩�- >_��wr���*���.ѵ������/�>�/.1vz�N'��w�u���v�<nѾ�I|6��㣁<U�B��/+2~�)��
�%J�P�{_��TT|�r�n�`,1�#�qBʤ� �s��д�b�]��%�L��d��f���I������=�g��VM�����hʙ�; �Ppf�kw�.��F%��0G���aЎ��0;X�Y��Y�d8Oe��?m�УW�?�� ��q��ƣW��V��AM���Dd]@PO(#��������;:�_g���-�����5��75��Cv.�
�;������%b'��T޲��&zwMB�-俀���Wg�Ξ+/���M|�F�%1��Lq&�e|���&_��w���Mf��B�`V��q��9q�.�r~oxH����R��:_�h3�P�n��V|c�I���K�ADCa�J��`�X��z Y��*�%�]|sJ�p� X������q*"��;Z�ݵ��������ˤV��\�d��+.`�13a̩��0��Rd��>����i�3�F�/,��:� Ko��	 E�P�7�{�c�^���� ��֪��%&�aQ󃫀G�vv}��$g!!O�s�� Đ����|�aJ*(��~n��oV��I�W$(O��YzFx���e���Eq��K��+1G��qcJT}��׿��7x# ��$̛py��'�}_����WqF�&�[�?��v��9p�aR �S��؈�e��K�>�� ���j�֫F�Vd��b�>��o�?��BR#�h�I��J	��r+C��B\<�ӿ�F�gH�TG,�#�l�"�w�U�Mغh/�ɜ�>]�I8�����d&JX�I7��/k*J}N�g����� I�`���À9�L�5ϑ�Y�����p�dP%s^��Z2`k9�^ЌH�(T~�&c�P�.�BL6@D}��~�p`��R�7?��_F�t�6�o$�MK������-����Xv[���L�ؐ�+��$O�D+�����2HM�"W8����"����ӛ���E���f����(��5����w_��N��~PG��HƿN���14K�q�b^�>S�!�>��_�٪����v̠hي�t��܇�<�j�/������e���]lα���)�����/Ѷp="�j�z�	�u�LǄ����6C
��V7�g��c�ꧾ~��ݾ������)w�$gj��|��3;��qj����nUFΆ��&��Y�s��_+mM8��(1}{�w��#	�A�a����C��٭;u��.A�y̤��9���4�-��F����?�V@��~���ֱ���W'�r��џO�\�ߓ�h��5u�qF	�!����1�Fc���gMwj��b{��UW�P,�T��"�`�U]-�<Xn�!���ۥY��(��<C��H��΍��S����\oێm��FE�T��T�ɋ��)Q���;Ad�<�#��#���T����}�pgɅ�4�p�=_�Ǻ�{K,^*_3z�g��)�1�dk��U��}K~J��ύ6�!&��$Ѧ�B���f�&�B4��.��`��������m�#�Ə��M����,ÏX�i�]i��ҷ�����`+����r�[,@��ط�X��E���"��V�����n.���Y��N�#M��V#��n�S�7�+��g4<��?	��;��>�]�IM�*�#����jK-�p��`�J��:��;}�*��9� �P��<�E_�a@�F4����7IL�k���9�ͬGMe!Q��Ϡ7��k���ㅳ��)Dvr^�?��CQI9��I6��$o��W�NL'Q�ip �/�<�q�_�c4��N�����_�4�u��mc,��rV��D�[U'���hב����Q�[³���N>��]��-��>D=o��3{��Z�Ӓ�kt�G�[�ecO�	pG�ݼ�s,�YZ�ȧM�WZ8(�M��]Fr��5yn�>U�&!n�(fD�����[kP��w����b�w_L����:T�Ɔ��ߺ�L�w#[�9��
����� #�)�$��N��cb��#�	gɰ�E���za8K��
��y{`n&ν�ld��&b�¡�1F���b�'E?PٽąO�՛v���8��(��f���� ���[�'�P\����>�.c����V�P�7�Z�?q�#&��a���B!�ϯ%cy�=p�~�8��g�\b�Q�sۢ�krL��;*��9�!���Y�Ls�?=�@��oA�C^d��C^��Ӈ��*4��u���hG^Iߴ��'.D����h�uFȞ��RΉgF�?i���kVtP�����9���j����y�_�pR���I����a� P��5�U6,�Cq���T �̺�9Zꧡrǲ?���������2u`���%#.������obp[1��}u�G��ۛ�0]��Sj���׻�P}�
��2:�q��?�b'����G�OW§�]E�$�ȋ��jM}gN�o�#0����9��7��_��[h�`��dF5:��RQ�.��������rpNC�I�-��܄����!b���X��H��n��+Hx&>K^���-��-�.���V�r0�;���à�91 N��H^raxs���@����\V�~��S�~�p�q�Q���l��B�6`�<���z+��tYG�G fI���Х��ր�0c��cr�b�7����(4�*E��"��4�^����ה.��{�R\#�6?2��>���m��|�$�����y�i����:r�1���&�v�z�^���;}��©�\r�iF]���y]p�ba�����o��a"�� �A}maW�@x���k��� �wq����K�^�J,a��I[���F�j�� 0����|�ʇ����~�$h�w��SԨ�p�I�H�;�C��Hyaː����RTV/o���>c�r�@�OG��c���u 5k�[ߩA��7�M���y�q��e�
F��>��O^�r7��1Y�/yϋeE]�kbO��Z��&������I��Ѹп0�-����&ԟ�j���u���J�װ3}6�-�t8��կ,�I���d9��0��4	k�^}�~��U��_?~��#BÞ��$Vz����){��x��8@X��13�glMD_��mȦB�֡u�Xl>X�݆��o�h}G�A����L�Z)��x�n���"`�>讂f�2��t�o���G��f8�궟 72{��O���|SJ�Y�����HO�ab�O��2;�`On��{�˥�)��4+"����y��q�.̿��@؂���t�]�Pf��i)d" �:>D�W�<����62�[��0�9y���S0x q�5��6�&qx�� ��7>#�(p�ڥNOx����^��U��bXIa��i7w.���Wi��X��?҇c^6q�F\�~R�Z�m4[1q���(�p���/�&��wJ��wǳix%��4;Հ���� 3��Ω+Dn��J�r��G���yV������a�,����s�L+&:@ND.�sB�5�b�㶱6�uA(�`2�t6ǘ4����jհd$�{?t�YY��i��S���3�&�U�Qd�j�\���CA���G��xc����>&6NTW�Ii���4�J�,��Z�8ky~}p&�C���y�FQ��j�n�A��|��ˍ�3��S�O�xULoRD]��G�q:�7�]�nx�ow���|�;�B҃y��?����0f��5�!d��u��F��c�c�{����E�*څ���}ư��i{L3��,<��7g�$�l���>�+:i�m
��nl�����K�� S��򱈸;ʊ1���OC��!Zmkv�f]�0�?IO�f�Py�5uB��y1�����[�_�6�� �f�K�%�$�;)?�����$R1R�M�ϗ�E����n�d��N�C�9���.ބd�S�1�2j��jgzM�ȭ._���ix��wOy��e�mj!abA��;9��-�utIoz���e8��#��*uѠ'r�^�����M�nK) ZÊ:��i)���H d�(D	�� �R6�>��U�p�\˾�[s6��!KXba;��{�^Gl���Mn��d��s�q�\�����U�5�,��A9�(g�� 0�]��1��B�5��8]N���G���g��3�ߙa�	Zq�q&_�� �F�"���o=�X��#�oؚ�B�q� LR������h�>�$�x�~A�N1��[�4|�r�io�J;x�u,<>���Z�����xS���������pO�V��|n;���y�a= �4R�*�z�s���$%����o��������m0� QSk�D��#nρ��$�.�Ƽw�QZ7gl^�����2���ѐ!S���b(I8�e�wQ������6�*xߣ�Pu�:}W@�|�%������ٲ�y�)�OS����?��K����Jue��]�	9�-#�4�qjy�T�;E(b:4���"�&$��ì	�<������;�����0�R �J��4ѝH�����c!�D\�������|��5�	�*�f����`_��.P��!���9��Kʖk�ZUetjRo��|̜Ȫ�P i ���dKJ�D�=|:����
�[�*S����X�/�Vx4
2S�(	�����)2"]���jK98�l6������C.PL_F9G߃��g���d��8��l�ˎ�V,Z�r��1�Ĳ�~=�K�@���֥�A�v�(2��S�N�_�֊?X��)�����MC�#�X�ܟ8�D�7S�F���2�h<���.����I�0�r}�M��*�ǩ^�S�xfS�E�:��J������,�k$�^]Ⅴ�=A�N�c�Z~�h���S�x���/��\,;�P����+(=/L�.�.��īU��
�e&�]��! %��S![_H��.���N���l;F��ä:��:}����� t}"/V�o�oR'�S�;���]7���l�åM�6��v��Rci��4������:�֍@	�P"��p�
�.��I,S�ˑ�9��+�cL�r��^+0��H�bu�+�7�jdbR��&�ź9�w����bk�Ȳɪ�c���SX�TZ$�*,8������ll���e@Z�*eTo�[�UW��oW����g��3��(,M7�W�w�B/��rs���0�ǥz���P؆��NP>�42���u���8��S���梸ݍ(9^�XT�s} 3`���9���9��x�W�R��{�2�b.@�r�T��������o�Զ�:w�F�E�e	��H�m���o2�Ԑ��qd3�6��20��SE���\?�yحF?��yo�z�����sv�U2y5v��ڮ�N����t0�4��+˲����'?���w�x�t�)�?���m�Rxr5�Jk�˰��/�`|���������t$0�N���p	Xp6��~�P��9�FH(�J�!~5�֐Ӄ]�喆\�l�c��� �<�~8NOJ-�9�U�"��
�n+���M�UDu"�r ]Y��p��%�o�����z3w���
�cj�V��H�}^td�{�Zn4��?X�e�x�xG�ףvX� ��O�4�]b���D�LƟ��=�k)����<��k���Eu��X��,yIx>(c*�¸0��ڨ����q�b�����ho�d �t��^4@'2��2�;��rO���Bhfe�Ǧ3A��%�=�)ن�Ÿe����Ո��,Vn5Q������<;��:*ćʵ3�+��}���p���H�H@|ʫiܝ�]Z�d;��Q��r�Y���o�g���@_��Z��O�剙�C2w:�xrW�{�T.�N��vp˜�?��C/y�[ښ#a\%CD��ȷe%I�{���=�2±U�>�-~��0<g�8_�d���U�8�\;�Q��<�B���~N�R��q�U��������`���7��W <#XtiF^Փr�Ȝ
��֠Ǧى�������N9C鈫k�u�(�0[g�'o�;�/_�,V��<�k`�
Z%y/rT��`	fM��@���Y��*{��lXd<���su�>��d��-.���{i�Q\9�jMC4���:�k�w�=�8,Ѕf���FO��-Iʣ |�v���o|э��,�Gk���u@�]̃�>4>&u	��]��dqM��6�8��5Rx����;0��'D����*�`"��2 w�� �V;��+*E��b��5�9P��G��|�g��,�SJ<��Wm(��zףSd'2��Jt7۸i ?��`��D���F�M�����0~Y<�ٖ���勤��6V����4�D����v��込�
+�Ј��R�׹�F��6���?�������:~�=;�8��6���*$��i�$�?"0�`��S�ߢ��dWp0[�W�:hC���_�f�?�%��X���iWҖ10��hW��&�o+9�+�r���l���V�
��[�t̙�L�ؾI��HD&NU����o����]��s7�5P;*\!i	ܻ����
S�����Jd�EM��hX�o�#�x�G�y[T�w�����d�{��i�Πm��In�Q�S�V<F��)���� В��}��긳�4Hu'U'�=S#Ź������C�_v`�^����Z?m*��db��	b��Uʽ_D�
*r��P�,,�n
�ÑS4���6�q�p�⫸�	I~��E���O��)[ʲ%]ф���L���$�x�y�U�Id͝?�Z%�LBa+?�T]2�u/���w
2v�1"5��,d�4ZU$�!�����Mg���,K��`혤�ؽ�rJ\�i����r�3#[?�����/c��t6�RW�ϲ1������%�� �5�nc��I1����Á/Ը�Wtdn]�1"��2 v��J���U�Q������[��#�	�;P���e���І@ːS�a �nA�z�w��tU!]a_ǚ׋�Y�;�$���6���	#K�s��eO�0C��n��"_�f���s���y%X����Yx��4J�~�Y�C}�\��<�O�4J���&���K��!�b5ݳVHGc��*iɈ�̄I�6����������5�_;��
#�a֨�@����nw,��ӈ�ǇtX��8���0�[pg�T�7��\�rj��	q�F������{�0^TK.�4S�1� ;���z(<��y��/��V6C�k�Z�����i)b�A[Y���w�rJ-�z[)��F����՘R���1�~ 	�	~�i�j�����KV`*�P^��E����&m��$�s�{5�?���&3$IDE�m�μ���f�pM$��|�{S
܃7�u6�L�������b/��j����"��-4QH)b@F�����`���*��+E��wI��m��Z[��F1���5-T�����D�G�L�� _
�Q���e�]��;���^���>��I������'��o~jz��Ӷ�v�� �]�q���UD5q��%�����Ln��5�|`��TsMgA;�,��c���X0D���ZX�J��������ֹY=f�S��5>TW���AB���=�s>O�����9�n��D��.�P�۩#6U������w�I:|T�J�+v���e�����`9�c�G%{���P��{.[�#��m�_cS��>���r�רeȨ+�a	}�/w
.�C>O{A�5�� Q�
����^�X� ��`�vd��П-����l�o��s��y0�4{(���Oڜ>50Kr�þ�R'�F}�,�;:c��E���b���`jB������R��ˋZ����'���^d�ܕ �yh��r�s	��C8_m��A�����^�T�^��Ya"tχM��[��ֹ\�K�XGM!t2�Ұ��7M�`}�ڭ|�.�=N��D ́�<ㅬ�k���Ӊ�]Tfe�0������oM$��L@���}'w�&�U��4�WP��5�7m
�cq�F���%\ڸ����Ia�_[R��Qg��n�ɘ�Jx��n^=�yB��7�z0L��Խ��(r���w�8X��}�k*1=1��z{"�7�b�("a��uH���<|�~���"~ļ�:���)2r#�B��ZeJ��i�����h
������k~E���Rk�_�B��ybGq��k�a3�$������V�}�-�#ơ���s�t�kv̉��Jک=����c������~��_3���e=���֞U��-x�����A��1��DŎrk����k����c5�Kj%��� ~�ڹ[�P��1�V�����a��-�e^��X)��h�n���5��t�ϰܞF` �����ڬ�p�e7���}�dl�����d�(�S�'���:�ҵjc�u|�k�y��q�Y�_M*苷4	�&��ʝ�S�1��g���Aw��l1p��m�*���ˇ�2'��Sc���#%�gL����PC��<���{�c����[�!�w����~���§WV���G I�ڝҥӕ-���"���z{��IRRS�Į�A�މ��Q����h�l:��E��D��!�6um�P�,L���^�l�`�N�������u:7�4j���Ǟ����j�x��!^a�a��Ä���;� �*�"@�C:�}����ܑ��V�F�
=���J�6�_��XREVa������)Ip�Hjk��;0�	ĂK<�L͞I���RFD��P���]'��z��Aw��h�~��T���y����Q%�$��x��������H� B�/��.X76 ��;cZ����>��jm͂aD������	Z��.�z",��Y���"ɜ���3r��3�q*R~r����\�Z^��)��c�D@]+R�&�b��[6�U��L���N�r�����{��ɴ&�'Wה�A�e��Ӿ��0Un؆�1횅�c�����f�m�6�,#"Ss����v�NX�_Vhx�s��bgImў�:V�{R��
"�����0���ܰ���0���)CY������T8Te3|�.Vֿy���)R�����G*#�#i6�=!cn�`��XVu�ե=驈�Y��a�������`�,�x(�t�b���'�l)NO����4eP���ނ�aM��갲����]�Y;�����]�ݩ�x���;�ۍ���eL �C�	$�z�D�$zaB*l���v\��uӨt������@Ԁ#Ǡݜ���Jd<�z$#	�ԩ:�,�!�9���jIϓ|3Bo�آ��6�z��>%��J�.����N��H�����揈� �2��xU��>��­����[��c�;�ٔ�Q�L��&<������'��T]�O��a�&S�hVm�q8��^"��P�@}Ց�&��(�R�7�8���,b��i9T��z�	�x��xr���hr�ە#�[�H�쭑4xؚ�����Z1$̭��r^�#�|ڍ��S�j,���gy?�o�g�D�84_��RѹAݱ�~���V�#��ٹ�ٓ޳ed|E���(7�#���p�c�Q����/9%FZ&��z
F��G�Y�4�r�����n��S�V�����DR3H�����3L\�tde�i$����-���,&?���"������!f��"C�~��,��ª������.�1���#�zNF���B��1v4�p�7W���NQ�!�D�\���)O�>�0���Y�n�]q�wh�>j%�w�v���G��k	�],xD3j5�21no~�����I��� W4��ΰ�%�����7>L�8�h�-�H�������Pq*\g6Ӟ����-y���3�:8<�޳h�͡���u����d[f��B#��Á��4$P�K [,m�{ۆ<��Jex05�������� <�tJ۵1nQ��������������.���t�Cx����[V���o�������b�F�5�8x����.h��yRV�n����a��j1�[h�R)Hc]�o���⫫K�u�hlrM��@�
�,���;�7�E�j�t�e�!�޼�5wT�ƹ{�Ɇ�4�X�
��3!�Yg��q�p�숅#��2����b�ǳ�;Ͽ H���ȢW�p�P���p��7����#u\>v�;;��<l�)��u��s����Ql�z�]�âQ]PC6�fsR���͹���x���2`�*��P2s/��#Kd�X��Q��=ʹ���.��������������(*x��*�ZD�R~unr��-g	���D-޲v�jB�:E�Oe�+���w���M�����߹Xk�;L��p�Z���sHf�,2�c�
5f{��E�o=��!��4��� dtF�Q>m`-�xx�<�ށ�4�����QzS�?�"��M����f�twBpX��N)���)�F�|&/Ha;1�ɲ������a[���]c6�k����bazvl`�ek�cF�ɜ:��U��Bm�v�&����?�>MY��!23,���<����
�O��j�h��}�2�5�J�F�8`�B��x�J���
$Dٗ#�t9w�)�q�*��+��N|������b
��u	jU=D�G�؃s|���N�_s�([#[�`����M=��[��l����;Q�n��/�L�i���uJx�XH�l3��b����1��vu4��U#L�Ks1=Q�3J,W�T�23�!}��T�r�3���>�JQP��/Wa-K�
t`��ɓ1_�!�}qc e�e������f���\��v���"�9~��p7]�����������}V����U:'�<<
G71��YN���jG��»�*�$�[�q=�$Ue�����ȩ�����X��kt�����Ug��/T��h�fU��!���4׏]B�����^��ڀI����et���f��rb~�A�軡i8#ܪ�$F�X/���^@-�2�_,�`���ts#hϽh�Z���TZC��ݛZ{���e�a�������8ف���A<��(d�(D���Z����o���eM�ñsf��J����T����d���;`�u����)��7&�p�"0!9@��I�K7a���إᑰT���:Н��,�x���#�oH=���..WE��r�H�cWV��Omk�/�[��l�b8�0;)R���:F�@�7PxhC(�&��� �������j��#�KT��$�(���
-DE����Q�E>�6����e�YՁ~,|,�Odp�'�����5��4۬���
F&�=��%�$W����������f�$��9ÿ�����)/�->�/��f�Ф7��;t!���i�?_�'!A��{Gj[9�p�6����$���`7:𡺀̴P�������{k��l]O��_�tbN���K#6�v�P�w�C��7����4F�O��g�w]�L���p�znS)��5��\�T�t�K�ą�Le���M�`�n���S8k��%�u2E���ž�s���S4�����'�V��sJ��4�b��yd�4߿U�M�7�<k���p���[f�7��I���E4*v���8H^�{�Y~eWn:b3��*"�#�꾹� V�s�w�!1vL�q(d�C��+��h�����_bo� | �v@���w<�F� ���n!�6+#K���{�+�����N��\?۷͟���]�AGx��#��ׄ�L��r@��͋���50:�t!�Zj詔i�T���{���Ep�،����J����d��bG�k�j8	�謴AxHL�.��#b2=��By��Icoħ��e�g�&����[���Ė���9�/O�z�d�r�n�� |{�y�9��1��Qc�]�����,���2�?jF6>���~uX�`&�%�+�?��a�Z�O��<w/A�X�Ux�3����3�p�|_�����t�ώ�"���3��M������]K_�z��r�`pK���w�6FQv� ���E2 �Q�"1f�K��L�a^B�R1��f�V�b��7va�YA���4�ԍM"L}��7��q$y>�zt
�����vJұq���9i���u\R���LĈ�w�_��j�f�yU4n�t��\�:�_A`̡&��:����u!蚈�p�v3�n�3�]�?����+?��,�m���i2wx�*����I�~��+ �n�+�j��
�vơ�uX�@@B���Ü7�!O���A9�7=���Y���6뉳���wN ��,�b��i��s%�����n�2؇
��e�)�;Ki�ЌЪÄ��)��k��J:1gm�m��(�K�0�Y��^]+2XzRZ��OĢ�SX�d7�XsgiZ���ɶ\�xsҐ��� B�)[2މ�3��3���q$���Y[e��g��1�q�j�.t��5��D��P��G��><	��'��Z���腦g"�UN�T�,��0W`���]GZh��B)#��F�ьJ �"�:kz�Nr@T���ӗ�cC����u<��OT�T��5[Nԇҷ��'f���9HԠ���9&=��5&��ذ�J=���)��������'݆�
ةfoxP�����T��ǂpC�^M����ݎ�N��8<�vO�r��S.�u�4������CχU�\��3�X�c%�u�uH�sH�~H��:G��0�U�C��f�Fdx-�} 2VD���(xX�L���M�a�I
��~�ד�V�ߩ�9Ҋp�o?���&-7'p�[��qe������y=����#N��K��D�GYق�`��R�����P�r��6g������ţ������:�8�ت-��߿�9���/���vfD��Li8�Z���n��Bp�̌�IS�z�T?kM�|%(�ݽ�-]��`�2�:Ǽ67��9�J)��>�*!ƃ�U��\?m�k���~$��s�^>_����X%��8�i�m��M�W�;U�S������7���t"�c�f�=[��!�9&Ӑ�ϓb��ٌW����LcϽ��[�����fL�!OY��mo�wT�c$3�%؏�g��4]��է�&_rY5������떿4��#�?}|Im~�+��.�	�]*��Q�4��$:>��$Ǌ�+R��1�"P�ֳ֋:��^��d�ۘ��T���T�<�čl1!����$�/��>{�S+Q�o5*�'�r�����V�nZ�mLvW�Q���8ć(���p���%e�~h��#�%���
ܣ��=Mڼ{�A�.
�c�64���8�T�kɺ�>ϵ���/\i���8;��> �u�b� 1��<K���:3[\#��j`�s�n.���"O/���ޫ�+��ʹ9����.P�a�+��Y���L`�*���_���xE��O~�Ք�N"!|M�/�Ð��j	��*Tn��( @�GwD��>M"u�5N6�I�VfQb�k$�3�:�>��/9SF�<�o��gλ�8*������������!Y̵�bC�wp.�$q<�7�_���	<PX�7�qædE`��4����2{�&�T�6�Qy��T�vi�:���-p�`5G�%��=Y���Z�������:y�K�ܪ������u����-�˺���2��;�*��/.�/��-����9����C%e*xJ_x�T�5=����r1PBpY�����i��75�a���m5�9)�1��'�}-�6_&��܊Ϲ�%���8
3���gGczF�.C�x�S����j��n
L���}i��b$��u L��?彑�4�6rq|��{;��ߧ�eJ���U���T�l'!/�Um/co�����źa��N��̚�D 7B��Kl�t���-=���_9�f1�'�n���8�A����c88��؋T0x|����m%�b����Eew7U泩�kI �N~�F��
@��\A^}�������ȁ6<��t_,�,VtTv�ª�4�]�&�Y܂�+Hi]}Z7��$�Pk=ɡ�wc��J��=2㺩�C��^8�k�ǔ`�l�P�H����7:	�.��e���I�`��|�^1��"~:e��s�x����4s��+r����~��x?����AsKT]��ad�I��X����?ۻx���0�r�e�g��bVc`m�~uo��[����PX�l��TL���8��6Ic1s�Y"�v)��٠��歆u�ۀ{�<$��s0AEO��ɵċ_:��M���p���,�K�ZR�?���a�Ί��Z_�+�1�]<g�>bb���:�|!�};��c�����ȨLh�a�7�ii�B`��J�aRͫh�̅'R�u�*�1M2Z ��B	���K�z)�Pm8��%c��Ǿ�&ň�Z�Z��x�y��O�S�\-���B,� &���l$������v���j1z_�DFj�
k���5L��Oi%V\"�׏䡷`��*=��IM��.���'�#zH�}�U� $��U��zTh������xMYRD�yۀ��Ń�=ԇZ/�gkU���p�Z�M�����_a�� �(���4᫈$�V��ĽA�¯��̞	��Y����`�u��:ȭ̫-�V��T���8����V�_O=�	_�p�չ�����z �4)'�޷�Y�hk���rq��@���.�Lq>����r�"����N6�r�Ͷԫ����\�N�s�贅�%Q��t�O�.	W���]��`�[�u^P~^��Q)�RSJ7�M%�X=���_��Հv���V���0��fE7�J5�53l�B���"�߾�{(L�b?1iģ�YD�l���&6�a���R�w�\�a��	I �퉟\����q��!�8�S�ۈQ���}�?��7ꌑh�^}��C��"�ᯊM��u�⤝w��1�6��R���-�?��d�-�/��d=>
>l�ݮt��۠���E%�-o�w$�$���g����Y�f�S<����L���c��g��g��� �&#�>6��[�H��(¡x�(��n[���7�k���Y�T�ͱ� d�M��/E��Zy�f��+6�^H�"���d�[-�WFM�����C���Y�����4[]��u�g!!L'��f�����:f��?$�J�B�b�<ýN����ˤ�>�����	.��*����X��.�(Nas�ԇwv��Vk��3�2#;�="^VV�C;����F��A$2��-�y_2���7�������,Y��T�Mw�ZP�����w�;Y�h��G
;`��н��Z�/��~;[r��9N������T���8޽�(k;y�-%5���hG��Z��a,�7���ؠH�n���M /��`�J�?�tkJ��ok��~��T��=M�Z)�t��j
��l�`%Q�ҩr��):���'�̕+�
hz�Rl"[��ˣw�k�t�O�I�Z��J$���A��2w�ҿI哐�r�2�x5W�K_�e�O��}&�Z,��mY��}F��^���%-���
��8����99i��;��PԮ�Nz�yٜ=�Ho�R��d� �#ܶ���f{�*,Ʉx����E�'���y�.Į��PM�P��Ϯ���A����7�[�s8#��.�Q�*Y8zR��
;}��>${�6�ݪ�q�`Tf�'Tb������k��*�'V�N����k �������+�0�B��EY��Y�:���I}��Jf����鵼W'�fg9z8y��a����?L���I�|�
4�Q"6"	�w�\E-?��� ���f P���؈��c�do;�c��B	��K4R]-��ix+[�h��r{cx�ҹ����ц���(Fc�5�S�6�֓\"��IP��/�7�RT�W!�X �DvW]��Hӑ�3�yv�("��:p����n	Γ%��̹ �6cוn�[��D5���lT�D��@U��/G��j�앉s�#ƶc�,Ҵ����U��o����>�V'�Ru���R*[B5��~Tf@��Buc�>^���S>̶�z�)�d�7X�%+�n��1[�]��.�mH�T��׏PT�f�F��,Kń�|�����o\B�:��ƥ�F�gc03�{D�h�Mb�<��:��?����3�]��h���Ӌ��O��1�WIF�_�~Iɺ��&�Ѷ�v�<�/����,�&g�]�d������j�Q:b��)M�U�2�p��ɓO������T9e�Ĭ���S$a������a�����'&'�*!��5�oB��3咞0���?�E�p[�x�7�Z�P���k% <N�x�"�n�G�
d�p�0���W_��*ljIJ��@yol��>�+7h�X��5����/����Ray�F�0��3��8������w|�}�)L��e'(z\FX�v	�:�4��]��`�Z�6���S���'�>CW��?�)	�y�`Ď�H5.�fi1v�!ۚ~�6ZS�޼;4�	�)au�T��Mi��{���1��ܟ�~�네�Ȑ�ZE*{�����ar=K�Pa��#� :+���	�NYИrlk��N�Oo���J&j�\�יt��r��wx�2z�dS��[Y0@D�>��P�+-z4����p�?)d���RY�.�z�ud�-7?X���3�;��%bݍ/����z
�8��G4hT�̿L�7�	]�8�[à1/1_3RCKu�H���U�h��O&U�4*B��Az)��Ss`�ϓ2v��ǉ���gs�H���_
�^�J�Ф���[b��J�㠞��V�${�X�K�dR<�`"��i/!�#�\�|뎹(��c#qĕ�3��\&iʵCg�� a�w�)�׻�������|2p���t��Hb�i1�Nrd)�2-��Mzxo�!�4o�0��-�T�VX7V�*U��?]㖼������I�#yl~w96�3ʸ2�Poq�(�������y�0�{�G6(h�Iz�{"NW�yC5���w�K��&�)q���c���0����"�z�6-��b`p&Y���W�=�c����*UF�q�W��� ���[�,��%�&Z��D�=0�z�)��XWn��"zs�Z��#}�e$�s�R8x���c����Kl������Q��=0\|�!4���O���LP�	dX�w1pA�N����6�G� �U/�7/��x�����[�v�2u�_�X��5����sh`�Z¸�8ֲ��r;�ڔˑ�*��Z�_sՑ���@�Ϫ`�V]Y�$��I@������(Ut+>x��s54R6���W�(=�y[�Wo�$�կӛ�����ՠ��^����bSC��e�#pE8(�m6�@����~qw�EG~~�����ź��@�ͮ�*�{|,�R����kF��2�ni���ԏJ�bX	4.��xԲ�8�LU[�V��!����a�,���t��UY%'�P�3�rս3���A%�cK(mᲿ�\�A�>�O�禪	�n��W9�c=r�:��7BP
�:3��*���~�\�x�B���x�|gp��d$!>O�%Y{��^m(�4���bEJ�h�Ԏdr��L�_m�p#"���g^�H}
b��&�j��Z��(��SV���Q����e�㦙!�P�l��ό5�9��\�&�&@�U*M��
ɹγ0T��<�\P�A���%h�V�Q*zB��08����9�)��x��3��Sd�g����b��V�["�(�z��"�繹�Ut����[�\����oW�w"�E��@�o�@R1�7y,X�֫l@���䃎��Z�e��s��R[ܔ,{c�y^VؙO�:�Um��}4�}I)ٛ�5�����M	e�Q�5.f���)P��Wk%������>�39�YGbd�u�k�t��$5���Hr���Y�4��Dn��o�(L�Yj���d�5�7J��y�a�Mν(�!�A�7_��Z��Z� bd���6��Z͠z���)tE�����AT�/�@��Z�	��$���@���m�������LH�o1o���9T>9K0�~e+�������'S:Ή�KfB�S*�S,�UH0gILF|ĉ�j	n�G���j'�2��'�!�d��n��$F��N4���)�;+,��R�C]�a�>���~I4qѶ`����h�D��0Z�,<'����	*���L��akY�d�??�X�TK��أ���x�P�{`W�����3<���y���x��04M�}O����$s�Z��n�E��a��@��`��Uα����S�ͤ	�=J���{['v%+�Y�!��b�m"G�Wp�y��==��6��Y���ӏ�����z��]ذ�:UF�S$ ÇLb[�k!R���?�1��Εz�B���W��\K�yҊt*����a!@�k�{�u��&�L��g���B\�%2Xԑڣ̛m����$ͷ�)���0���d��td��26���±Э��`�� �E�/��;ɿNFF���_��f��`9��BFu�Q�+y��7�~�wJ���B>ğ��x%c��NGTw5H���+[{�Cq/6BA���r����;MmrPFJ���kcA��ׇx�*�K����)���Ɏ��|:��z8��Bׯ�F�L�
E���~ځ`�B(e]��?\��U^K�sYLk��ع'V�ě��o˄�"����aE���s>]�4*ȵ'!qx�$�?��"m@�����^ER}?��HG����,��3�Q����"aʶ�=�t�&�F�w�����j����E.����Oo�PK!Ա�ە��F[�����@�\P|�8�E9��NÁ�#��K��.Q�@�|���zr�wB:��]�x�8��0F��'�*�/;2�~.++�O�Y��o�f?A��6��m���y��0۳^J�Ef���%'}���ޢW�@��*�L���|�R0HҰ�����-�]�슏y�>[�5�Z2���M~��=��DdRT�pՍ����0��)�>��Uح��^��!p�:B9��ЛA��O�t 2�7j�3�a�	udZ�U���E�K�����NYi>�U��nԛ���vo���K��,��rFe�O9򬡠!%@/ص��o٠��6��e������l���8얠��1?�K��'iv��Blfs��x�@�Ƀ��FF$/[s]9����l4���?cQHe�CYm��&�T6�|։��7�B�PBD�&�@
�ނ&���Si4��N�uc��`��&,�,:� &�G�Y���+��tr
6�v�Z��q �ԭ!A;��QKp���4�F��ק�?W��7��c���&p �Wp�&��"�!ݐ�O5{J�-�P�ߵq+E�֚K���:"����Do����0��U[�J��A�� �_G�uJ�w�x�b�"���Tl�t���`����<^4G�g�d���0I����r%�Is�������3�T�(_d��x���M�����~u"O3i������<�.�W0��UQ��ωLpf�6J��Dpg�������2{@�'w�6�c��S�dus�����9qF-6tD�]��
�� �N�����ɝHΟ�eM-��bDW$-�L_�gR@	��I�(X�윌�[F��G]b���%V�s}�h���
e�*o��S1����wt�i�?h�K9Z����yЅ��'cY�'���H
�V��u\'�����b��
��'@gMpF��q�͡��lt�����/?T_W��#�����$��}�
&������3�Z1/hә�-��W��S��MXw�����cQ<0Y>��3�h�E�.|��-��oW���D��,�+l�=u��Q��%�}J�@c)jAic���d�k���J��H�bʰa���s���v��V�⭊gD�=����*�����;�1`�!��9^~���$e@��&(dL��ɪ_W���Ygp�ź(z��������d����ԕ*�6�3��5�Y�O��|\2`\�lv�9�K�RC��]��{�l�\\�Ց�40A��,@��g����0����p���"6����S�9|�'E8x98��E�7��׿c��{@5@W,3 d���~7K����6�P�è��$ټ����y���m��o�A��s%������췅�G����$�t���X�����{@��^HvK�,/L�Q22��G�!J�{�R���r��gq�_8�}]�����M�/�,�Y��l��' S������4΋���y����p� mΖ��	�]m4M�)��Op�_��>ճ�l�/�ee�K��J�;$H�u����]�;��#~r��99ѷ��)iu����n��������JK`T.'�$~P�C�H�Z���qHʬň�A�l�zyr���z���e|���� /�ӴJ^O�z�}� �I���"��>�e����/Lևn����cQB�U{���}z���j���*���%�j�z;������w��D���C5���?�+�0Xٹ�-Z<D�(P�,κ�S�D���(�?�>��D�����plaQ��u�A����[�d�.����zf�.w�<A�%�s��]e|�.	��ֻ��if{v�ԅ���]����7(sE4��ZXt�Q���%����0tv�������AS���1C�~V�1� ��<Nq�d�P�:��x�81MS�/�$�D �=/�
\�|W7+�V�-�H��T�9�Y8ċ5��:�2��Ȩ(=�Z�G���"�e�J ��q�+L!� �v��i.\J ��V��iC������p��NM����8c~nð鈹�2y-�(�܁��vk:מ;�	X�WT�3o�L�gԆ� u��U����l��V8 ���m{=��RU��n؇N����w��[Sb�����E�߁8m�9E������'F!c��"z�.���*_������*ōqEȚz�0/��Y��#��iX.�X=��z���ݬ`�v����(y�v�2ø�n�a�P~?���w���n!:�>應�[��kws�:�⇋��� �%� T�9y�FJɨ ����Z���� �v%��9_Ob�Zi����@'��/�ɠsPn:�R%���ZM.Z�qjp����T12�c����P���)�f��:8���l4��.k�q�m�u����K�q��f��l���R8��2B�`]cD�揃�1N�,�@n��3�]�2���-4�����h�!;ċ�����s���;�)=��i�8�ej>���������}w����j����|�/��4��b~�/�����ߖ�e@�5����@1�7�s.���~���uv8���P+f����[u��v4-�W�����e�?�P�)�	)Q���4@7���# �]�e�U2��ȯV=��E�T_)��n��e}(3�=C+S2	u%�H��R�keK�c��
#�bm�@bh��l�R�[�%�Z�s������x�GHIt�����
4S�S��3�r�(Ն<�ʝ����_	�8'!��o�x>�u��}ƞF\*�Z�TED�`Jpo���|S+���9g[WdZ*�=�̚%�7�WPē/pO���N���B����
�5����������B�3���e���6���Ss�-9O|��f�H��A�}ơ��W�d�O��j�Ǥ�È��%��3:��Em�c9I�W�+�@�YN�RM/7;c���a�ӠwV����ڨ�{���$#���n�%/��.\�7 ȹ�47L'8�1�.RmUgKf�ρ�,��)���8�m�1"�B��?�EV�KI�"� )YxZ�;u��U|���c���8�8h����>/�9־���"K��7w�P���w	�xM����Ko��>ȢӨ��a9��H��oA?���^�ZmA"���Qݎ㞝v�O̹տ��]`ߧv�,�ΈMmy�����;�
�
�kW!��>�%$a�q�n��)�ul�����K�i�ZJک'��_B�@������?���s�X�DN��V�`FB@��9��N����$gD����6������4��5�;ͯ|��[�*�`J�
�m�R��?�V����a��1�0���.����>�� s�4��r���Wj�Yк�XX���u�i���!�ӭ:eI���42�/��Fm#���<��v�v��{�pF���P-��W��՛yVBj��e6�B�g�<F��}q��.���]7K-{E1[��7l����׵R�Cgn����r�O)V%��D�b�a� �b`�����Am��Q#e�