��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Z�xX�GPW��si���骿5�շ��3��\o����u�.n�Cez!�������8�s���&Ĳ��<A3����֛W1�<m�7�p��ۛi��*7q+�/	�:q�F=�@�_ڟ�]%�.���]A��>�-�X��;�W)"�"�����y7�m�u�m�ٰ+�Z�&>�7���N]��uѤ��a�m��&��􍴐ϫ[�/�{b0��Go�{�7��jc�K5|X{άԝ�Μ-�e��j4]���J��D��s�;��c C���:�1��w1�C*}8~?��r� $��'���,rO
f���m�]���[Q; ��Y��Z.����K�����7��qD��a��7)T��8�#B��	��>/�"�O��i�B�H8��G���L���\s ��$��#m	�|MiJ^�&s����A��qęY�O�U�U�2�l!C�7
�N�茽�/l��#�������V�< ����c��u�'�q< ��J�)�ĺ�i�����l����?��ǃ�’8ؖұE��"�[����-d�K&gu.�� ػ�[�~�r�=�����s������&�a�i�%�����r<V�ym�1.�m��f�5R	D	��a�ǶW��N����Q��|(�h�E���v��M�������bt4K�j'^}-�������e�O���׎D�����d�{Z�j�U���*<�w/t�>�K�Pw���B�")�1�ƇL��ej�wmN��ݜ�����Bk���vi"X����u�	7�4T��n}�hE3��$��]g�b�0{��/Y|x>M;Tz{`�U�.?�0[�!y��& ��b��D�6-Q(;��N�ަ��8��G�����]>)F7�m����[��:��"D��@0�3K�RN�c���x�X�yey�T�����a�'ZA�
�R�{���� ŭ��}�_�'ҋ���RS��v�:O��KM�1�~ۮ����v��q`4�'<��a��o.��^�몡]��͐�%���\e�B��b�m��_�xe�{˂�q����{?��
���̻oCuΟ	�z�G��n`ʔ�$<׼�@�ZT��*0�%��W�AH���~�q:�]��L�#c�6�=���2�g[��֝�~j����M�y%�UґޠH��Қ�>q��P�WNN���_�i���m�z�o�@��)>�6;���}���o�2��*p���cA�c�����v�Xe��<1� � Qz2ۿ�~Vn�{8-�!ǵ{�S���*��.PR`��ÑN���y{� gS"�?#P�ƫWJ���Mq�]��Kn<#s��ڐ��]�����Cz���C�z��3���_�p�ۆ�&_!Y�Nȏ�sm��_�N&�>ǰ67�����B���S�S\����s�,f�~p~�e0JבP���D�g��W9.��L.g�����w�����Slؚ�S���@O&��hѧI'��#�,��xo�{mD�n���((��G.1�avԛ�ƴC���B�O�����{^�q9Q��V"RE��|u2E��B׋�'�sd�~|RO�"a �rq�;J�h���4V���2��"��@8�t��!�M�q�Q^N��M�y!B%����W�o��D�}�X!&gү�y,�6���!Gk=춆�2�Jy��ojMk;��.�e'����WO�'[LӀ�*S�oP}�;���3d<2U�T��Qb�T6���X�kr���̷=�(͒�b	� ����G��Z!H��Ip��j�����q�jx\k���`���y�G�u�t�/����R�o���z���J6s��q�n����*!��c�EÎ�?�8�l7�mOF�6W���#�ƾ���I���\C��{xش�K�N��_�Z�n6Ǻo����
?;�y[�E;��)����9��?�S���T��Iw=��:�	�eSY,@�+��@��s`������/�y*\�_L�N��l�~��z$z)$_�72t�*6?^��fuˢ���������&��	;]V-W���_�ށ�;�i+	htQH�
�I�e��� ٻ�0�3{�O������ W^����6��ժ���/a��!U���\��(JX��x��DF��q�!��V��m�`(#:6?��X.f�RUC�o����t(,��;��"F�ٍV	*���E �C$��7A�,5C�M�&�KhdD���7�x��k��މC���S�h�+��V���-5�U_�DM��N�~拎En����9a{�	�OX\t�n3���=�oxc'O����p=w��LBM�'��>�e�3+���fj�2q�ө��H'u1�R�e����������4�����[�Y�be���o�h�m��0*H��Qd�&��B�K��9����G����e�̓�#��xή]�n����F�� ����΃u��Ɖ�Vh�࢘��۟�� �4��ymB(��Co���T�1yM����\��NM�~�J*�b_i�t��P1FJ�����6Ƨ,%�pP��4_��ğ2зex�U�\m9�✍�8��{���py�04MFD�J�5"��U�r�+^�s(����_h)���C��}�����)�Y�EBD��a��:Є��	�\�jG#�32�%.o:֦;����.G��#���L�%��πw�|�9�ٱX�#�g�g��H\�z�c�? :�S-���]P���ߊ�h�gqW3�z'�/P�g�G���$�U���a3,�$�(�hz����e���cc�*�F���� ;�Q��X��ຐ�w>���$��\"����*l�E$%��D���F"��2���:�{%^���ԇS��a��)i|��Zx��L��gA!t�\�Oz-^�)6�D~���1\���0ġAٱ
3�c�Ċ}du ��mU(�cո�{cn�n���̦|p�����z��@�D_l2�������ˇ�a�,�1�����<.<�W����3�_u�j�M��u�Lv~d���%�1r&�eqU_L�M}O��Lu��`�rE�/��#��׋!�/NXC)�.�o����T����������O�[�yz.	�Hh�M��G^Y"kOz`�E�k	SL�52m"z�ڙ&����AX�8��=�LN��ǟҢj.,�HU�`l�ϩj�z����m�J��N��?1P٫ �d�z�9"�b��>�l�2�_{.�6����
�>wz�r���9�%��l����j�y"xك<r>��7m��\ZGF��P������+��̆����m�Ǐ`=��2F��
�33��~�(g'X<��F�H�}�w����L�ڈv��ϗ��/s�=���ͬ��f�]Q�����瑖���.՞����OI��kI�6m�#Ĝ���o���x�Аb�P2�˵hΤ��9L��t�[ Ɇ(�PR�ja	��X�0C��0�)��
}�T���S_7�Eύ�B�#̌��-�����D�Bm$R}�}�������V��s�cpP��7XYZ�Ne�%�s����I<M	���B�0��t�-����I��iSc4~�z��*���ot盰W�c�X��C/.*�a`�=1�5���nƳ�'�Tz�l+:���w8؆�ѯi�i��j��R;�f@�!GR�c�;O"_���Ѷ�m?1���SbP�G��ƥ�%Ot<��f�	�oP��Z&�w���O�px��5�`�77�"k��L�>F��|��W}�u��M�{�*��^ ��4��G�π�	m����'���-)��q�Ȩ����iƍ�����~ց6;,R�Ը>��3kSd���ږB+m�a9�7�#�L�	B�cދz��ж!z������2ݔJ�A�e�Z�=쿖�K�s�	�/g�ft'��܌M1��p�<bNB�Z@����9;�r���2Fx	��m�c��B搆 uцmJ��O��`�����[��#�*�S,x�ٙ�f��̣��DE���(S�ȿp�����x_x1�oP��d���8Q��r]����D��
�?�f�|�&��%f���r{�,tj/��dU@�IHJh[��]>�|�zuh�?��@������hEg�w.���R�݋��J�6�������PF�}��aou��?̃Yn8jyUT�QB�6���0��5��\�%A�����?r���l�+�O��aJ�c�@���Qwg��/|tn�ܗ�EqAi�Ȓ\8��>7��vq ��; ><�Gߏ�LJ:$KjA���Q�r%���sn�N�X��������I�*�N�qq�^�R��گWa|v����XHM��#����m�^�v|�������W�̛��IW�\u��c[<]�qB�h PXu�U(Z"��&c�F�����A�DW��K�^� f}�"�0�l��dRUY�����J?xN��H<���{O+��;�\��"��Q�����z�o�A�a��jt7lj=��#��|��Mw)Nh�o�ض�"MTBY="1������	>:Ze�@�Jh\�����Kn�*��YY�j�U6�i�Y
��g/7��-5�<<rܑ|�?T���!���ju)�/��Z;燭V�e���iv��e��z$�7^#%�Y�3� �*�4SLr�L�Ճ
Q��!���w�m)�F�75I��"�T�w��Ƃ��LZt�@^ �q�����q'a%�h��#�%�ް��s�a�^S3Fǖe����D˧5?1J�K�vO���kT��>��۷W�����X�P�i���m����������#V�b�3�r�3��w6}�Yz,N�9=�ef�V�/Zt��x�|�GŠ��X�8cr�y�'���р�	��@�M�FL�!��:=i!���g�`P�s��!�~6�<�R�
NF����� r����9d$�����d um]�5k�Ȃ��|��\,bں������|�B�ѕQ@aQO5�y��*��rK�i�g-:�� ��ꊫD�L�djGB��<�v�u����.G�;�i"?JB�d��*���>���_J��S"���&O���/��D��v8�E�e��?̤l�UQv�/#�
�2g�i�IZM�o��5&-�_/(.���lYo��tq:����q�����?/<i>X�Y���O���)�h����2^n�����w��Җy�$/V�Bƅ�(%{Ki��<�O�T"�g��4��MjRt|#E���4��t�V�T9�k����L �� ���G}�>I�u�p�������u�r��Z�f�[�BW����D��L�?1>�~/F94^N�!V�t3�[�Wݭ���Z8����>)�Ԍ�����GU�R��0^*Ɇ�� ���ͮ���F��ف|�ؤ_�^��8N�@v*hN��A��I�H�wZO��c�ۘT
����pu�"E��MT��ՠ~,����_���4RQ��L��ߦ89g?hr~ܗz�4+��i�:u�:�rE�-Q��Ի/�I{����)cwfhVDZm�S�w�h丟]ָ����B3}AZ��~�ƪ���}�0`����<�����5��?�l�eHc��bm�K��v�$��#���2�� �� ,5y5H��u�0nN)�>Il���Hr��Ĺf�9��dH#��{`~�+���8��c%�4(�/��ok�$:�j7
`������(L�$�CkƖ��G�ׅM��w�ū�R���̴�7�o���FN[X�3m��;�wS�B���P���W�bЦy�z�m�pӞIo(�=YkMi �Ls�P>�]ڼ�<Zn;�J��&�2���Ҵ�6 �n�1�Q	�G�Vԧ�5�֍G�
���Q�zn�M�1����L���bدq��`�m���G�ˠ[ ůP��GVvB�~��������zo�i�V�#���	�1sQZ��o-.�Q��N ��rw9
��d KҠ��eRk�J����>�< 0$͠�AT����=<�P ��_� 	�����s�4Jy�����1����b�ҽŕ���
�h�|-"�2i�޺�>�pwz�%Ϟ��ԀO�xf���]0��xH���_J��CwAm��ɾ�n�<wӃ��}�
c��еH�=��^�C�C���~{hH⧚!R:q)�AS��(�S'h;E1L6<j���� t�ϲ��zp��|��4(O=͏�9�����YC�;���&�ɑ\�+�#Fq����~��A8�j+$����=�2[]B�����7Mv�z杻��VA�(��&9귄�k���Y�y�h�L�\8ڌ�8sDQ����������D���Ðz魳��{�:��.�Ӳ���@��<��m���x�op�H�J�W&b��g�W|�ٗo��ԅSp�?��n�o(���6�� ]x�~Te�I������tR���P=�������3�n���k��^
` A�65ԛ�njQ�W���)5_V�IV�v*�V_�{Ng�6DXG���@��MI�:!I>��qd���L�҅\��2�(�A�So뻱s��{m��D��
z�Ċr�Kg��f��f����i���AZ�ZN�"��U�@�>w֨`{�w����]}���| ���K`t�O�l�,Z��c;���g<:	�&{�Bɻ�f���5���G����7fk�~-�O�y�:Wў��軚t��w��Չ�z���	6{�	�k�s�Z>����[�[��Cqы]���7���C�al���4Ĝ|n�^��òB�q���_�DĲ�g�(EqK/%��f�"����l7���b|*�g�%����P�QR���)�Y<<S&�
�i)@�v�td�<�1�5�?�uv?I䷛me�M9<���=5_̾�*�B �W^����| ����V�n�l��[��a�N��Q������<34H8��5N�gs����D�w��a�z��|�A�D�/o"F��4yg`PX�F蔗d�h�+sz�3�Y�d̘�8�+!?I՗�F^őV1j"���N/�7��\���Y����k+����>t�f-���D��X��+�āpQʒ5�
�r�5�*R�d�6uh�-m����9ܭ&Kl�w1��L��Axcg(�es/��Z\��)I����«*.�LYK��R���7m����f���U��^�7N����Gu�׿��oʾ��Ca�s�� L|�dzg6��I����Jj��^�@����cp��6�r#���ֽC[~��#����S����r,����yEudH��KY����J���L��	d�������TH}��<��T��%�|�?P���`�?d�m�N++����Z�G8����]�SP��p�V�ɇ�ڜ�k�?��gZʸ�ݒߺY��߽X�g�a!�^AY}`jg�����w���j�#��@�yќ�'ZH�mI�]n�3����Y��q94֎�Ȧ�.��h-�8)��b�>?Вi�^r����+��81������wѶ\��^��Ro\�^��1v4;:���[�s���Њ��?`[�,d�;&:&��r^��Ƞ����4���x�8��;�_b��J������b)A�6��:��6l��WVJ���j���+�����o�oy����j�����8)L��q �%`��vf�Z]�&}���_ڒ�p�&(Z� Qݭ�-m�J: �8<1/��i�!.	�wE�T��#�kK��@ݱ�(U˟6��Q�X�h���(��a8#�n