��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� f
���O�Q��Y.#�d'���J�"����4���d�"�Ŝ9͜����
�~�a�rN�����o]y����1���nJ�]s 3L!��,���zَaw�{,���{�b�[;ҙ�u�\��������.7���}����H��ΰ�&���ے9��y��y����͍2��ё(��7q|U9��1���i��$>�[�G���^#fU����S�"_a[7B��7~ez�#�5��-������>[{Љ�v��G]��Ew4��5`�|x}��4�y�z�f�|#�դ�e��5p���1��L��d=�㺔��y���h����V���Q���t�̿�rբ��6�j�mcP�iT
���c�j��5�j�KL��tlV��d��x�Z��"ks�kCK�|�i(�;�����6��12�XTeP��[��'�0u ����r/X�<��/�]Gȥ���%N��]84����Uwp)
���un(c�Åf��J��f`9Fqv]���+�<�w �N��fѧ�h ˞�C;4��#�i��T6n�Q�T�����ڸ}�rS3�*�x�٨�j���y�~E�s�~+s�G��'��%`+�w+.}��(Jľ�$SL�2-�M�M�W5~���/%��t%���0;��3��G�rq�Ħ@];
!}ˬ � C_3ZjT5�ъ���29L��>ԡ��I�#iDn=*oB'R�؍����v��< 2<���oc�M Yx�R5��ܡ�����2=ړU��oLW9oq��4S�um줂f�X+��t)�a��� R��M�Ć8��,=���LIQ��[��Z���9y�ڜ�|�a#��C)*�uL;櫲Q������:�4�t����I�i��w�k��Î}���ѣ�\��{Zin^[?�����B�!a�hF�`7~��$�M��]�'�]��1%6�̬����|O%�l8�$&��l�إ��VI�0{ʳ�NvFɹ\�c6
��q��Y��a̷,��g�>ވ��k"R[�o���=Az��p������SԈ#��e�O~7z#{{&&^��E�?	���-S��hU���ܮ�tDy�>�a�����\�4�҇8:��Pxp���@�t�
�|�P�����A�Ev6`F�^t��������Y��Lu���(o^u����6��t(Y:�&w��'���11O|F��-W�A��}��O?�+D=�h�D��[t��_S�R։f!����@!�?jNM������O��L�W`,��t��ׅ\HT��h�N��t�JG{��ӆ�|z���^��+�H<���dˠ�R�|��3�/�j�bN
&�5���{CS��1e�G�p
���A���ǌv�����˺ޚ݅��������7�\�ǿ�Ӏ!��rɎ�D]��-��C��K��䓶��D5���乃S`�zx��W_���p��ݠg�Z������+�&�Z��/~�&j�Z���(j�#�WaD!��r[�j�9{���.uq���ؘ��sU$���K�D��
��r0U�"��S����c���<��1��	/��v�穩n��.���<�	�����%ހI<ǭ��������Ne:�Q+��j��g��3�$W��G�.vPt�s���(�������ѵ�lfB8�N:_LS��/�֐�����iM�s��*l�z�"�#:��m����&��cFή���iVQG�*e�*v�&vx����}�v*p;A��{CJ.e����L��PG�a�D�d�������6���2"�W����a�� 6�Z�	\}���K�;��|��b��&6T�[�_2�d����s?*�?��3{TA�|�ȣ�R�Ǧ���Q'_����bV?!���	��z�`�t<F���t�f�? �P��P�Ey�4�Ǌs^
~K�Z�n����`|o��3G���1��9�{���1#������"��
�����͝<W�ۑVI��m�L5��{+ݐ �S�anUNkU���Ę�����G��%rH��/Ȭ
侨2���� ��C�T���tl�qؗ��Gkn���k�b�A<$NT�yk1���ݜTq��l�-e�[��}�d�xC�7��PMQ���]�$�:N�OcPWNK���	�P�o��H�t���c�sΠjTq�)�<I�HG��f���0��?��-&�4�s'Į��x<Y�F��yfi���'?JNwJst��I�o��fI�~Ra~�k���:�N�X\=��e��_��&.�v-0(��]��/r�ly���+�����c�G������wۂ �*������:%����O:Wɵ���Mvuf��q޳����������2��9��	��٭ ��0������T��4���d�N����|�ZP/�=ǉį9�ĕZW�$���mM�7�H����L6^~)V(?���*<�Z�&\HI�@v�"���c�XG'��֟{�0���']�	42�=y�@���gJ�p1���ǃࠣ���nF�t� ���;�޵8��;�[4	m�G�M���P��L�2������A��:EO����^(�v(��Pa����8��_S��M>��L(`�	2����\{����MMp<}Q�8,�����`���c��̅���w~r�h�ο�V���aTQf)xT��rc��/��Bf�Tô�RXPWt8<� �N�wY�W�����a��Limj�K��n �[�U��	�_���D8{�#��q�����S�� �&5?��t�R��j����*�o�wc��w���+%�@�"�;\%�Ϲ��-{��x�8z@�����l�nn�:ǎ�bؓ�I���w	��;2�[�D���2ż���?�yaZZƌ<Y����������ڏ$�Eg7e�t~Ax���@�x�%��(b*��`�:�>k2��̾1p����|�5O����Λw��I�ٺ�q��ƪq�jB4 .fQ��0{�^�s�pjGW*��qۇ�c[����B��1Sw!:!�Я'.�b�/o,l��v s�E�����g]���BG��l-&����j��S5�*@[���g'b	����P���{hw�m, L�Q����z��-�,HB�?���Mzߗ����d���BL�yi�N