��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K��mo�G�
����c�LI$��#��%n*�D������2
�<_&A=/ĩ�vT`%�2�@�Ӯ���bR�)��(.C�>�M_؍2,��EA+(����H_(�Jn:2��f�1êPb5��[B��������ʠ}iƭ�Z�k̤p�<�7b��F���� �[��GG62�&�=A�ъ�0����+�5���_��#k�s�������ю��pD�*g������Z�w�D=��p�7�X* �K(�M��<��lB`	��z�`?%Z���X��_櫿}�{y�0�Zi��k �25%o)��e��VI�� �͙���sY	�x ��!2T�4�`.Ӝ����d�X�(_� ���z�-wK�il�|�B�©n���A���0�X�>{��c�������J�7{�A��P��^�3��P(�hƵy�Y�v���Ⱥs���\(��xi_���Nt^9�=��Ҭ�I����8����Ԃ�H[����`@��kK=^���88�*;���t���`|�ؒn\[ϴ,=�F� v����D96f��N��PO����9�$�v�k"J����M� �du-�sm�z�hR�\���䖥���zßw�=�HUK����	�{��سDa.��_'�Y$��	�>v?gي2�:A�x�Q�OC\6��E�M��wӏ�6 vF�`V��A@˭��H�U���[8�^�s:�@�F:�?K�c��V�%�*͞k{p�j�`Ѭ��yA1�/^*�O&Cwt�^*"Vu����D].@b�7�ʅ�yR;��*P:^�(D�I 6��=����]q��?��w�j���e#߿�R�v����}Iʻ�K��@vM}����g��ž`��8���"e�X�F6�ۓ�3�5���5��T��+��x�s&�&�Qf>B �y��f]�5fs�
}�ʋfV�iF�F擴}U2 ��ْ��{���\X]9F7�F�k��&įE0r�
���6�s�*-Y�ٻV^-"aYdb�ZQQo]x	L��K׋���j��ox�^�fK���4S�?��~6vy���s�[I=���Nl�!�r\�tU�s l�n�#��i��q���	�W_ͧWJ�5���zG���8�����"D�<|��3-����
t�e��7�Ei�l��T .r%a!*��������J��r�����_��ݹz�V_>���&������A��4��������Yٷ��~/?O��2!y�h���+R�ڌ��UZQEA:��l�zE���� }6v�L9J�J@����8#�k�A��`�k�Sy��_xU���A+��b~~$����My̅{�I���LXg����<�X�u��o	��|{%}����OT�T��A����'�'�\L�br {�d����\�?ƃ�-��}�w���!s� ���㪋L/�55��{z2z�*��y��٤������\_�x�e�!��W��>�ڶ�g-}���
�,]G[=�	�l��7���7PI�l�����HN+r�����W��� R��tɎ@_`}�&\��GPb1�:yõю�UZ4��5h�h�yl�S���ff���(�<�J���z\w�ۨ�� X(�F��Ǫ��Oj~]n$,<X5z$OM��q��%���k쵸]>'3����W������������iD��$}Rwjn�����'Z�39�M�}M�X�l��;�^AD(O���W��֚��>ܼ�5��o����`?Ī�/J���r%R�?RI6�T#րa��g�Å�j((fjy�~:��im2P��-b���4@�8L��<�{������9�[f��_E�T $�`���u���7��Y�Bl�;f_�f	J���k�6�y��U������f��qRl�z����@����O���	���� t�b����/Q_�v���^>1�E��9��4{����N@�P[�7���Qp���6�&2E<ݫ������`���6�yg ���VY�U���?Q�I�&xr�W&���	�������l����'Qvm�DT<eJ��xNV���S]Hf��5m��,N�4�2Nt�UF��Q�����8��^HZ�v�+ �i=ԍR�Oʉ�YU�+�t��������!����%<�P���1���ni���3�R��Q�[ �r�h@��1��6(� �?z��ځk2
�L��*����oo4�qj��v�Hf�!�ŌE޲���ے�f���e���W�w�t�ط�e�Nx�ǰ>= `ܾ!�"�P��a�3�~�}��-SU�fN�8X���?%��u��q7�,��E��ֺl|t�q��5H�14��"����ZV��O���2��d��"tL�QZ��F����'��"v��!�sM;̭-��h����1��&0���2Y�v0.R�8�U�J9���G�3;(���f�A��1����I�t�T߿�Ԁ������<����^iqtm*K�B����I���]1-��!�u����*�?���y������[�o'}Yn�{9Ϥs(��@y�TjZ׈WNy���~�.'}Y=�bfs/P��0(�^b@����vB��@�h-�gd\���Ѣ��JU��Z�X�L���7��4б$A��)h����M��J�
�����7��;�ѷ�2c�Q��X;��s��⇜T�&X�A�T����9��'��M]բ�H#=)>�ʤ���Ћ2
v�rO�{�Fa����NŭC�>�%��<�w۰Y��n_�5�E��'[�?�T�_,��GV���4J���=%o!=���$�QAؼ�>�CΝ����ʵRf���k�z_7��ZW_��0��ƿ �`B;�P����D�@hY�x��� �/Z'���Oe���NA��E'�Ѳ��5~xaK������N�SnP�7`�P�!�O��F��|BcsNLa_3�}����1�i}��ާu�ߺ�6 ��P�Q�C���χ���x� �z�F٦>���%�owZ�	�IJ�5�Nk��7�F��LE����MA�k��v�Z���^WᡣAR�X 	S5���"�&25
;�uęf�?n���%&.���tm/ 3X.Ec����G/�� �t���%���dt$�ฒ{',)��b�X�0��3�3����Yy?�xw�-�P,��U�������c.k=���zͬA�oh�;�y�9	\��F�����@G��s������4�������N}Hi-�f��e�Ɲ4�xZ��:��z~O�T�>��������R��-`�ѴA��@[��� �k�r�)�@.T�&�� �ޕ��Z"�rq��Q8b�1�Q����ъU�o���V]�ջ<�ڙ�QY�<�6Yqq�C��f��
l��S�/�+�&��F[��*���v�Ñ��fy�)�jk�E��I�#��(