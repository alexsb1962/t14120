��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+�7;���I8������b�bM�D�czC%3��B{;�德(�����z1V�`Z(�+� ]�{9�+�:p(Ve�B.vvO�*���ߒF�q�I+a2�jV{�*�����V�T3|4p��,�&�Y[3���;�)�m���){=7Z��/��,u؄Z��Ǟ1���|(U��m�+ޏ��K��h��d[��s�"k#���mvТf��I�#�(_dS\��x�`a�>=LjJ���z
�eÕ�id�6"h2�Z\�	�+;A-Vy$�V�9�z:� �y��"����@C��Ӣ����:�^�"���
�'j�q���O]D.�}���(�~��t�vI3�KG/�2��t�Ƹ�-Y���! ��B>aM� ��q��kПS.F%��8����~��ϲ�QSP�kU���V@7|����+�~!�Z*�K�5�6�Ϥ�g����q��ȳa�=̶�&�`�+#�ʐ}D7HB�_k�zȩ�g�L�@&��"N�'5-��k�v�M��S��
;Q+<�r�"tS����ک>>�1(��������Ur�4KG�^�V��[t�@�{
��gh��s_g<:3��� })�2�¨M����/uYF�=�O��#���vx�p@,�|I���k�����x]¤3�*p�.�+�*��5]�;I�����*�#�Y�LY��o�ͽ�Y�m0�v�Ȃ�����ށ�
�[	�=iz��6�+<�h���-;�X6�b	��z�8��6��������F��:�9=�0���=�,�L(�~��,����h�e�*ӏ�� �ƓL� �{�l�3�.�Z��]���Q��H�-��+P��d�����CT���h��5�Y�`X�.����J1vg����G���_0yӬ���xC�{���F��!T���UF�<2�t/� ���?�,�
L�y/��#x��pe��J�y@�~b��S��"�0BU��,(,f#h�pnH>8�\�$t6�k�J�8��	s�i����Q�X�& ����Z[nr{ݜD�T�8�
�<��?�E�����7��*������1�!����!��
:-�Y���`xO���GNƪHe����\�� }E��*�l�/�r��q�bi�/���	p�O�� �G��/.K{e���O�H)�к�W"z��6j2��W��L��pɋS\(L���rV�~��`�l�%tzԥ�>o��
�t>�nsH�=�lx�#������?"H�i�a|c7G�d�ҴեU5�U�^����YC{��������tE�4��� ���d6�t���U!�8���-e5����9H��NC�@\������B]��G�E}�A2�����ޯh� �N�ぐ}Z�b3��[)��s�B�7���g�����ݜ|'��Z�b����9H_c��J�
LP���(H
ow�!Ȋ�)2��@�����-��`��of������F�kɴro�X|���Lw�G�Yjs�h"ο2�{3�S�ϵ��T
7�"j�4ĄMFKI�<��� �����D�ru�m6�z�Σ"�:AR����E�9�9?��=w�����4��������8?�<��/y:Dnrt���mB�� T�J�ʀ��O^"UȬ��
� ���U$�B�Մݍ{>�R��qgr�1,B ���D��5��rip����Ä=��}H��������/Xd$�<��{�`2<G&�Q��4����âą��x�V�>ҏ�3�5A���i��?��y��I[��"w4�^�+�&����c5�����A�0�[�����J2S�1�B���|�$p��	S�ͥ G�N}��1�����m�EnK�
���N`1��zlU��0W��*O�U��po�^/����9�7�����?�/o�0ڒ�3�g�N7߆�	<������b��SG��0���)۞�\��as'�e�7ɢ�\�J��J�>����'�}���
�V��r�ɂ�M%|��$���q��0�i�r�czP>,mI�:S^#��꺊�lΰ1�m&�Ђ��"y:#$�����ǠÙ��u�R%[ƫ:Zf�avIҩ�f�xa&�	3�$AOl�Cz�:��&FO���Y��M�IM�`o*xx�E2�5<bލ|o
�����X7�ڮ