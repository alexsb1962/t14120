��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`p�l�z�����k������2w�%��G����cׂE�D��dF�����/p��g^���҃\��%�KҰ�}o�AҍXGܕ�_Ɨ32��ٟ�l�d��'���甹q�����pⰈ<�Ӟ\����c��ML[�A/Ĭ33}����m:�!zu� �B�2�z�V�B}]g�5��2x��~�ڢ���/�'H=�D'�K�O�x�i���B�+�o��qU-��N��T?�r��P�����u=u��/"9�*�W#2b�0�[� 3#�:ye4����m�Ko������<c�H�����H>�
�ֵ���9C��~����6�P�z���4���7�����t��� Ć��d쨯����o�7�ݍFEgO^5�Xz�f��S=���RC �=�\��z��H�K�T�f��b�T��Q�s!�����d�J׬�uSfݴ6�<~�!��՝�`|��"vj���N��%�X���p�;Y>a\)uC�L�+�vV*"Ϧ�]d���س��I��E�T��Z�]���B�����2x5[�k+�'?|�~d@�~�*�g�O�4���#^�t�m�xoF��-���� _]w���R�_�CJ󙻥�̨դ��7cs/D���$������ƃ��Y����!���)f���c�1x\���&� R��꽞�j�G5�w�F�Y
�;��g|�]��w�!�%U��g�y7���!�Ի���J�4#߫��ZU��5��E���7dy�ޣ\ �xW���-��{C_�>G����]�Q��4���Mg]�tZr
&�iaz�syUm�:.<����]6�<�R�BGZ��+�+��71���2�`/2���&F/�S�66���*.���)������X�)S@��:�C&��5shT��Ճ߃,��6��v���Ԝ��wҍp��6�{���E�`2ŧ�� ]��ڼ�f�+�St�TYղ�0����X�}�b���#����m�;����z˚�W�dayV����Es+]��S�W��!���;B������{J;�����mԔѻ��3�.�3��G,�|s�����&Dz6q�v��O�YR�L������;�L]����ߩ��#�?���Q��brMq�O?�g(�^Gp`�P�0(�U��-���ЇЅP0_�m�.�ص���BOV/�i�)>Cۮ2q��E��:��T�,#.$�V���n�Ae��*����X�V�x,����ᖘ��&�{����-
*���4:N�ꐶ:��Q ֨h2�W���cW�	�Q\y޺,�����2����X�}�9��BM?�����Ƹ�׹.��E�J҂�7��>���VPJ�R�Z�[�MJ�3.�-�iʚ5�����[�zI;r��^3bs�ZVF��"�+ө�\�W`�j�U'Jwz1�}~��K}L�!���"�S%�K �L��Ş?~G{�M(�g�-�y��,l����肛�]�%�eg-΍�\�6b�M;�9Tڬ)��f�V�g�%�|���k�m?�wߕKΒe�'�-辪�Tb�)��
��ք��zռ���JH��3��eaǠ�����C6���	Ƭ�s��OR�~PLz`���n�8��D�џA��l}��}TU���S%�1u{)� S/�i�I3�.՝O�X�v
L*��3X_�F)����j`薩'qH�6`-l�ٻ�*dm�м���n͒��4�
o�#�h�a�N�N�4�U�#�Y��ƶ�����6���Xz-��K@�$&��X�1M���-���uG��-��'/߅=��RB���6b�t�C����݉�c�M~�s �8�d-w�@d�4WV�ʆk<˾�������.4�ۤojF���j	�Yͤ:�Z;C�Uϵ�}�Ʒ�VZ!� �j�;j���K���G��:KQ�޽ו/e��S��}�g��.j�Ӡ�N�p!�4G��zw�@��I��PN�6�G�+��ʪ��M���c@�+�"�����z�4O!x{�[ƔG��׋����&ldV�"�F-�HW�Ȗ���_ۏw�:E�{I�1+��P��I�m�1L��	����Y٭��x��q�Ǭa�WH�v��eH*���P�pQY�Tm�э���#��TZ����k���	[i(d,�H�L�P�̥�s��=���i=��
Lܽ�� �l�f!p�6p�����J���%�������{�%��EB+������W�a�s�xz�t,Z�wx!"t$OV9��8�H�xvA���iQ����U�9��CF�� �fUܽVQ.��V���{_��f ���lkiemUs{�k(⥭����i�[�ǵ�N��kۏ�}�y��j�jq��ު3�wY�\47��<~��<Y6��+G����M�N�-�}^&��q��4I���W�t�־�힑�|���##��k|��-���vR,�ȍ��*�Q�dW_V��� K�Ll,v%B��t��/�*
n?���* ���*��jqrt���JUg(Z�S�fD��+��MG�Z���ُrN�%���S0�jU5m���!i�⥱e-�!����3�.�-���.��{���o��|��R]��KKz-"���i��JK�)��3�)��ޥ\�v�����ʨ4����0_'�h��
�u� ������?�8���+�@yO=����QY:wI����:)��!� v�#}�+0/��}ڡ�ͮ��ð�+4p%<B�9��'��>�,�~���x��?�/� G3���ῼ�Q���G����/���l(B�M�����O��������Z�sH��%	�@.V�j�v|`s_�����W������ ���{��J9O�����_^�u�N��h������Tx�s�+\)˞P�w�X*-#� o�I��c6��8����j�s���s���鎁Π��EJ׀)� ^��GTLVÔa������0%�P唇���r�W �"5ku�Oې�P�����O���|�%R�V,y��4�KƧ��K]�9�le����"�I����1V��\��hZ��o;y!�����4�	w������	8hD�صo�����N{�>=611�)���d$@�U���T��ט���y��!�vM�4;�NpP���J�U�-OK��xFX'4_�}ٙ'%(SL�M#����zo`8�
.�og �O`)�3�q���a`�c��l>B�'��+��=�QDBu�w�h�!Z�4�ֽ#.!���k�
ޅz�A��
��V�1��ԫ�1*{����������6v��o	�3�5@��b+��ꍐ;�����?�Q��4������|-kr��i�V�C\��`���f(ZtaVP��R��u�)U�ܝ;���"U���l��I�t��M{ԫ�B�x��u�ta�K����"W��`��b�m�N
sxS��h��!�lP����<�h&���ү�-;G��z��*i�P��˻�jmۈCJ�Fo����h�㖩�����v�T��Sr��7��[f��*�M��"��6�h���ޠPGV����xcK�c��O�[�q_f�)�����'����\����`�.�R�g)x�4��R�Ϳ߰�.U��!��YM.w��ci�$oxf��u_��c�И����7�9>��!M��z7e��^�����E�s��o�E]$y�P�ʯ'����ѿ�����6��̣>d���.��]�~��v�:�14�0�_�_�\H)WB1�2B��ӗS��ׄz�Un���n��̯�*��Iw�*o�8�1�B�
8[)��i����(|&�D�w��c��b��R�0[����r�x�3��Q�t(\k��;�ia:	����I�����\��`��-G���ވ���ɑN�Ok� �ׄ;�W/=��$b~>Wy*;�Uu��y���4��	�e����Y(�[6>�Tn����6��+�ڛ�Xr�����!�툦@q!�w;]M�X�ᱛi��ZH����.��S�#?�y698��&�����Vwۓv�E�I�qkKô"1�j�`�H�N��M3b�)��Y�_2���~˪k�րI��� �����N�t�|�I�1�tɄ�S29TÀT�J�R�ÔI�Yk�aZ�|P�5V;�8����eP�^b��%�\���F*��Y�ǗpDk% �Ό7��/ˊ؟{6L�4�,��WϪuy���l �X2DdA�Ot����d,~IL�<jMG��4�S�9�����#ՉfgG��L��F=)�L{ڴ1K�n�����1�&*�d\���)?�#PS^~��_��*/���y[/z�!��-��"�P}n�O�e�� �9W���3}D�0x��Ӆ�f�V?G}��aԺI-)�;b\�� ّiڡ+�z8�a�@�Ź�]A�qh6�0c[�ܡ��ƫ��|+|MX�8a �9��mws���P�7~>��`˻�E�G�s�N�����M�8����l����5�6�G/c��s��ca�bB)�e����8�|�oc~��56U�4I�Wep�0�Z"�fW7�Α׷��Oa<��Ҿ���p��0�?w=L����v5)�2���[�tKa(aZ�eZ���V���:����n��o^�� �@)N��I�Ԅ0,D[( bjX"D�P�6LN�pu��*o��f�Tj�$�w|�^��z��{���hI!C�g��K仳5o�d�W\?X����V�R8�R?�/�Ffa�kE4ڱN��fj&�UM2�%�������^���Z_|�^=���W�j1�
xSr�������9bk�]��^TY��m� ��L�񚺂烈�
a.?H�0� u:1�*���h�T�mX���K\6Ԛ�[EE	��N���\l)٢Y�M��a���l���1{q<H���/�l��<��_��Qn�U����F�`�z~
}~�>h����O���K�O7��w����#�i�#�g��L4#ņ�du�����Եپ��N���Y{�����`^��#�1I�9O	��������C��d;M2�b������$��Q�� B����%"����M�b}� &��x��4�T�6�qR��	Ţ�\t�;��M�Th�!���
^���!���A�~ؓ������q�/ �Ԙ�M����-
; z)f�wY]�GQsc���4ӳvj1ñ�����`�(f݁��'�?vC�4��.���AνU�p�9O�N��8ƀ9�`WG0��pH�������"�{V@�`�{�|��{�
�M���s��:=f�j����7�7�6��X��XfpS�?w����q5�$��0K���F$_쵮�]�i����P��\H��Ā���D���u>l��f͞���C�kJ�n���b�̳tG":���i)�Jo�t%v7~f#�_�$�>�C�d��G��b;53p�^&�{}ݏ�DM_�U���y�� v����5���&�h;N���l�� ��ɴ=����b�|:�֘ي�J�?T;�ϿT9�0�ZR\������Z\ƍ;�=	\g�3���D���E)w�Z���_��V�z���Q_+C�~MT�_�"�3�wF;��P�P�K1��U2�arx*�jp�4����ά�eZb�i���6�/zC+e{������_�8^�vD�S�D�e�������)*�oV�oH[P���P��N>�@���lU�'zN�a`L|+�������S���^�����<A��L#�t�G��j0�g1����f�B���2iJl^��#>���{�mB�5�b߃��t�0�Z�p�i��6\�j6�K
��Gr��K�E�Zڌk�hN~1\��2nY��������X�Tu?���,�G�$��h����N�5Ap�S�Y.�3�QR��_]�'z�f���RB~CX��G}��^�w��KH3����a�t�S��-�0�_(vI
ǯ���A����&����߸�W�*��	N�k9�+�R�`�`>��<(�8���S`��ʞ7�6'[!�P\�s��ְ)_��������d��IafN��� �S�s49ZW�Z-�W�E������"}`iT���������"�m�_tS�C���?�fng�AGyh8;��ܸ����[g]T�΍,�Ye�ou�(:N��}��	��s}P�ie�΂ؖ�k�o|~"����B�HJv��}�q�k��H�&Q�a�JL�����N���!c���Af����ҍO�Bi���,f��P�"�izSaA@��eu����_(�:�E���Q��q��y��β��a����@�G\�o�W�����$M��x(ƃE��8�>?�|aFO����<�
��%qx�<bn�m�ZJ_T�w`�����9�u��@���+,�*]y�ٹf��$oc��.j��n���O2�g��M�!IuH|�W[�;��rq�����ϫ�!?�z��9Bb�<�kC���])��C �~	���OP'��%�Q�:^���u��x$��.��P�����lQ�)���o�?����ɸ6��Ķ���`q����u�bcuRI`��cM*���_ ,/Hti֪���? �x�8�+X�UܾAU����o�?�t4R6?��`�9�|�v�?���LZ\ʗ�$P��
ק�~��ܵ�@��wy��F��2_���J#��[)K�v�:��B���j������s&?YWˈܓ��O�i�� �@�_}�����;(S+�z^�/��f�џ�O�݀hc�-�]63R�ATw
d�e�xݪ�w<#�]#� ..K�8�Mޛ��ћr�:.�;<m1�L���;�I�2D
 ޹n��|��j2	�G:T��@�o�l�ཹ]��FS:��Q���61%���S��KG�iM�!U� �6MB�:�I~�s���jO����-N�/���x�q�Y:���ܤ`i��7gX�K��E��Z����Z~�ځ�cD����*���顨D=���H�5�A5�	fMH�t6���(��khF����6hք��ʂ��פgh?� 2���|�͚�t'�%�k���� 	�΄�B���	�ݣ�R/�mULehԂ����!k�C�d}�#~���OxtGi�j���"�\:�gid�߷&]����5
�����!!f�ʜ�g�~���Y�$�f��K �(��(��@S\�S���(4+ש�i��%nh�Oɞ�C�&U�
���l�5Ty��,zb|��0��ic�-Y%QB�<�����?�v�R9������l�]��Tpf��X?�^6}�\��GOvN�	$-kt+���՘�K��C͠���_��BTL�Cu�G��e��2C�a-����J%�~��D�d�d����"n"OuOvb�)ie6��&Yʪg�Q,�-������['4��MGF��V~De-�������M��1��El���h���7]���/�Ց�� ���ke��@�l���r�"��}�r>DG��F�l96k��Ԏ��b���DP�9���!��5��:j#*W��|�^Kߋ��	�_7�K�̞X����Fw�+��/Yc��g`
�`'����2�Z̪�!Z�N�3\|%��h$ե��<B�AQ���8��X�X��1;����� �@���Sô~���#|В��g��Hk���E��[���!:Id�hv�$��&�a?B�(�����Ȝ�4Z96�	�{0� )�r�@��'��*l�_�a0O��9	�޼�mq�Nb���dݤ~��(���u�pcW�r���凊fE>�y��,jf��<-{�{v��Q�b�����@4�u����^��j����WfEfm����bq+�Ɵ)'{����S��8R�#yی@�6�7*�_�df�p������`,����wE�K��R�Dӻ��/%³�ď����Y�*0d퍖r���)���vP�K���C��XuKe���!v��,�+�w�8�þG�ʠW��v��@��dP�!��q����#	�V'̋5%ϩk{$3z�#L��R�i�fUGC�?N�`{!I��h抅C0+�10JW�	��F�-��<����_*E�B ��+�gO�Lnj�S�@�3�tV������V�^�	uSw�v�/ǹ_��G�%���O_�q��X]3�L�)�(6�*���s�]�q@� ��#���H������Ź�H��U,���1�����%.���p��,F�r��}b_�G�Ph���7��Y =��l����*m��;�kW>l-<�4��Mg���7��峑А�{�u�/��U�i�]8��6ޥM�b�����	����{,^ˉ�G��n��`�,<�oyR:\Yݽe���}����趔�Q&�����`x�T�Ӱ��NScUj}����v�=*7����5���H�I��C����3c�M�7/̤.¼��f՛eI- 1v�i�'0q��1<���>�*���;"�4 Hv47������g��E*a�B/kr���D�8y���Otv����Ҟ��z�Nu���A�L��'��<" ���|�����.���/�Ky�9�p��h��<I�Ŷ"�IPr��Y�B�c O��K��;��aiHrrC[� ���h�0z)h�6�<�^k�G5�m��;��K	7X�>r�ؾ��Y%B87���:��ۏ�2mYs5����w�z^��F&��������K�j�S�����*�Uj�P��[��Bh�՞�W��`��ӹ9N)3�~!w��f\F�ہ.F�qS��4�-���Xi"�L?���~P8=8���#W:xZtz%Ҷ�3��?����`t�҆���kR£��}��嚗v�R��XeL6�X�c�軵qVR`�{&����P�Wt�q���?�I?jJK���Ҽ���@�q���.�f����t>Y��)��>H�ޤ&s$H�Ow!TZ�1p͖��
��fMc���x���/���c<��� :�mEP���ѭ��t:M���ő��������Teԍ�����C5�9t_��͌e#>p<4G�\��/$��=��7⾗�I���O&�*� ����sp䰯E��d��)ũ�1�U$f�!:=��P��~!���/I%�
f>o��P�d�c�3���d>��I�b�Qh����b�	
q� �)�:yY�{s�E�?�e᭤O���`<rJZ��OlՉE�y��/�]g��t��<�m�r}�:/��p�<��R�'��mUD��)�ݩ�s8,��ۧsJW����蒐�f#��T'���Ki�
 �}m~�7v�(?���$�:9�=H��/K��O?vKd�&�Q/�����,�K�U���N�pJo�4���^D���P/�3~w�愸�!TSOǄ:��<�� Z+x��������ۅ	���APy�in�� ?�?�_��a��=���tlq�ZQ�p�$���=�챧�@ذ�j�ЉQ�����ի�ƥ����n�Ye;@���!�9��>e
�H����`�l5���tȬ�2<޳39�(�����甠���h~����E�c�g��\>��d �x���x0P�.�%X
���⤸>qφ��ݴU�1���i竀1��-w
Jcf��XL�'4//�=ܮ�����c$#>_���7�e�i����^��뾾�����U����G	x*�� ��:臽��y��\pj�%�-Ƙ������_�W1���E�R�Yq��^�8�#j�.9����RW�9T�j����IӨz{#°��}v-�1���̥\�����T4�0�%�q���=�M$x�2��KeZ�<(��,�Gr�']:ӊg���j�?zV3��g�S4"�Z������ |�u��/`"�-h�7��,���;��z���b~�I��@����GU�w��}����F#�� 	!6^R�� iF��v�	$xP�vՆ��[�áˋ�ZͅR-74��A6KԬ�%Q2�岲��eKpg<4��q��͗��?�R�j�~8r�%bg�������NiGQ�`�ı���f��	~S�������D=�3��Ef0���Wk�����W58��Ū7��HwM�ǈ+* ߖOO ���o�3�ub����!�N͆@EGZ���s��F�'7d<u#�r��;����ǟ�2�a�"mۘA�<s&mN��:�DP�穔G$l��ʻ�s��)9��<����i�G��
_����9jgr*�K�֭w	�.�Ո�#.kՆ\'���rS������g�Ēӕ»P�m�b3�%^���ƛ�6{i�,1�#��T[�s[X�B�%װS0�!P{rtZ�F�� ��G3x�`V��>���]�$�u�|&f`�J�����(�,��@\��qR�1ޑ�:V��n�׶q���y��2o�)�4M�-�I-]{�l��=���V��g�І�vzXwUZ���$x�}�*^}Udϓ���=�}~2~{�x+̮�(7E<u��ĩOf��;mHF��#4wO���l������}�qS�#���M�^�T�D�"� �敥�+PEOE�/!��1p�95���i�����
�W�8�=��el�dO�;�'?#��S� ���6�����m�Wc+kI�C �HX�f�FR@�9�ڛ���>���:���d��xb�6���bok�m��l��C���*�9�nn��C-iЦ��.ҵ{i�X�83(Ku�i�^���e���Ѡ#?���a+C�X������Us�HE�\)��gXr.�Í����R;zl{��;�JbCZ�����E�Z��[<�._x��e�F�t9�SJ��gU�����ȑ�ӓ4��)�Wʇ��U
˥hѰ_�sx���F�NY���27�����覣Y��+���f�$��C���U�)*�h����/��a�2!�����T.T����c�)me�5��;�8��׹Hg��nCU}F�a�7��)"*������=���Ku6ؖ�t���k��s�ӧe����%`�iq2y��[AO��T'�E��l�+�=����K�R��+Bz 0�����5�X8�%�v&xTO�r�<7��7�uţ�j�Ҏ�\���A���5�O�#��::�q9�U��ۓnC���k\��KxJ���ґ�ޚt�2ʰ>�'~��j2.�1_�a����0�+�>+��n<,�\A蕌԰�"jv�Y������ƪ��x��P� )���(!u��KKB�<�	ˋڱ���gи���|���D���hg������a�q ad҃f:��#>Q;�8�+��?'��L"���D�
+硆�G����C{Y\YJtˈw��4d4��Lo�+�5�#&nBh�~[l���O㫝A7�5���@���1�=��=���
If����QTr���@	P'�ܙ����]�w	�J��P�xP��U�zC9�^R͍H�����ط�w�J�y4龔Uh�(�eI]� ,�z�9�k�07�5.6a
)���c��xG�R����Ӎ�2��2+S�D�V�b�՛F�� �j�luZy燰5��_��٭9���Vf��n>�@�g5A�?��#�~���xF(I�3��p�%�O��}�(��h�׆h ���������?2��;�Rên�7;k�h��i���4bg����u\��uōH����&|N���Z* ��"�٨�ᷕJ�)>�l_Q���}h��PBW��$_tI���{���u������w���t��LXƿ�H�0-]���]e,�&�j��0���|��d_���6U+�����q"7g��v^>qx�[� ���-��	����W�B�[K�ȿ|�<�'�%��� ��"�&�u<;��v�����x�r��Aɧ�34F ��/�Tx�O��2���Z���t����G��g��rF�c�BV�s��glDV�F=�ܙ9T�z��W��7o�t@�&
տ��:�0�~l�p����D��3:[+�4�S��U
m^�}򌅷��.-W���fG�3� `�Pk0��"ڶx���H5�x;�OU���uz�����ë�~JJ�8�t22HSaE{���!M�]�a�T򆖳���t��a��I�»�2]K��~R��u��:�W�PR����w�b6�\2q\˼��R���9yj-;,R�"S�c�~�h1r�����`�����-M�ze��T��`���K�a~[�Ȅ�嚑�u�H^�Et���>�&,x+�q|u'�#8�m5�V��Y&O�)MBΆ�T�i�cn��V2�u��mr]3
2wc+�6ΐw�.Υ�R��)SY[榉�zX䮣�'��Ԏ��l�( \��[�[��m;�]�^��]>HE~eg��p�C�8:�<�(���5
H�SrAh����� hVDo/�1|�y�>'�)�A�Q4���:W׏�m3hF�˒��Q�J��:j2�xan�%���t��D�,>�+��I�P������>�G��-���� �v�Ç�AE�U)�{R�+�r0�!���)��ܒ����˟������ŀ,�<��3�6z캅�'�$Wt��1�6�V������]Cw&$0��.~n4��7G `F:�o͕A5��i���ޡ!���p�A��u�ۆWj^ǖ������/��
v���]�����ߣٳ��F��h�jE�:�®' �^�&n�o(8�4�ݳ-[�	�o�[��(�U����X"Q���^ �Z����h�PN,����/Ȩ���'�/; �sf���¢0A
 ?$����mJ�jN�mt��ﯤ��V�+�=;P�X/�EEW�Öbg�e� ��_z�ج����}��aa�X��]TM�c�S-���=ns��ؓ
m�TG��,\�%�F+S�~� 4tXe���
��*o�dt<;Y<)����V�+`{���[�C7�g*ae�����ஊ�����.���$�Fh��,r{�N2|{S|�Pd��[�D%�d�zu9�!�j�}��K��絛�D�o[x���^�u<����w�û�^��FD�l�R!E�d%&���i}��}T�I߸s&�������n^h�T,MHB0+�RF���qg��|� `i�=��V�iy���`ٴ������Tw3 3�V��2�"��<.\m?SMI��`��t�[��c�9��܍����~`W����P�ޑi�9Nn#��|��(�ʔ�߷/�ĝ,k=އ�o�Bp���ȋY-�Jh*wp<H'���X��i wKcP���<	(l
a���N: [�_n�V�'>�JL�6A����޸���w�%P�V�RAu�z�(_r��'�T>��+F��z���4]ᜏӋl���o���#.��Hs1g�略1nn�p�T��x���2/ :ج��"����"�]D��Ja��W��ͥ���v����Ώ��1�љ#��n����j�B8�c��.~�M�i��2�$a��BGN��S�Ր7,f����S�NKw�1 �c�s!I�����!a ��:����z���Ox���[B����5/�D��*]�6�A=�Бk?���3��#ǳϚ&P��v|s�UV=����oZq�����pJ������.��ʄ,V�]p?_*E��B��)��,	#��X!��}9n�=��J�elx��,��Y4s��CY�)UK����JՄe��ʔ��b!�	��s��U��r&�!w�d3,�=�q���5!U7�S����a�y4��O����q%����U-��­���&�����wvm?��S����\^������D���+#�\��'n�!3oG}�k-ܘ�;D	��=lY.�o��mWإ��|��Th��D��|����@����d9��@�N����|TR$h�y(��QJ(|���J�קS�tJ��^���=�[}�+ӫ+>�q�c�Q[�>Y�j�_����ZN�Η�m����,��i�lq�l��qE���7��1�%Y��N#�<^k��� ��%P�]�?��9ZP=-5�zH8܄�)8��B���	~ �=ü�4w�P9�n�G1��z�Ot0���!NT�6t$���H�.C!��F�u�/Ju�>ɏ�.���fQo�a���m��!� RB1t�a�-�q|۽��n�t��s�<�M����lPĶڒW��hs��:ݭB����V�t �|��q�7�ް���u1!�����_��l5�˴��0&��>N�v�$�W���o�,ٮ����`7@0
�����z��� �+�t�ݠ���*l�!m	����\Y_y�WW,����ȫMJfo��e&��T��Zj��i6���F���s�->�me���?��~�#f�3����_���,@�%�~A�M�rv�ջ���yR�}��OBS���K����EI��P�/�Iϱ��-����\�2)8gc!��F��k�oD0�g�b;VQ-2I	��*���0�8�w��{N®ӧ���%c�i"l����(tLm-Z��e{�Ͼb���2�v-A�!��U�v"�V�K���fq�h��1��HRBX"�J���f��m�g���e���*�u)z�Z��0$"T5��yBY-�W�նw��-����o��zw	�w�V��$�`VY+d�'��Ʊv��f*�B���_Ʉ&�e^�vѺ.�\�]�9�k��\�Xz]�,b!��f�[xw��@2�{M�[���hc�֭��ݴ?ձ'�|j��F��)P�FU�H����6�ӷ�ܦOA$���-� .��~���ͤ�/î��J~��Ő�OJj۞@b�Ba�w�u�6e�]Ѩ�)q��X�R�Ilm��=�6��/a[]th^�F�f����3D��;+d����(1Muجx�پ�[Z"���{�E�q��?��R
hC?�Ia�.�5h}�E~L!�ef��� ����$+\�bB-?Q�Ր��]����2_7��Z,���AW;�7��͑�؎c;�RB�GU8^N:
�_�Nq?��Uҏ8���-q� ŵ-nWF�[�iF&b�B���9zm ��J,�:�Prl�+�ˉ&�ޤ�{h{����EaO����Mn�%�_v�sOnB6�<az�N	P� �̹�]�	zK嬟��$2��܁��mb=4&��kx�پ/M��X�����xE\��+	K��`餮��De�P�g�ǡF�UݒeI�IY�@s�R����zz�lɏ��&����I�,�K[���}?.0{l�{��9�>h��Z�L�����;)�<,�ᥤ�J�+���ex�:��i��@�p�t�]w��܁[q�*�)�JE����
Գ�RA�\��Vo\gR��^�J�L���ӗ��'��#�̑<��Il#&=��� �I{���AZ�Y�J�FH��˔�)w�h���v y�ؓڋ�����P��5F0��l�c���'�؃�~�(;d�h)� |��mTԩ?��?�!��=�ύ�"�[X����
��PCU���َO�e:kn��Ds��TyS�D`�N�P�q�v3��]@ܾ.k�R�JM���l�-n�,M#R��!��u���8����_~�d����*��\�^^|��LMYQ����r�7�.]�Dg�����T�����-҅z(�î��Q��X��[��Xs�>�ZS쭐��ZE���	=l�,m�9�s��|rѤ�R^�m���N�Kcm�t�[������(r�
�$ڶ��X�[�I2�K�THg=Pr�fl�P�� 6���6�ɐͶ�H�B��=��6�7���)�Ѓ��p�7�w�D�L@�	P�{$X+�c%O3���.I���o�pf�i�dF��{SYKEK�фh!ܘ�ޏ���ΐ�'�)��J_D|�d�ԁ��`������ƴ�<Ebl��˼ț��JK�U�r��W�����I��.�x]ק�Vb�N���4,8{����LH�S�����qI1΋{���Z[�.d��i�S��$���=���H��x�t9�
o� U��g��K���N�Y���P<ޱ-l�@�ǁ��ޱ<��&w DI�������c��._�e���L/q�����L�'e�g|,�UGK)�\�#Ԧ+F�ym�M������B�ץ�ЂI0Xۏ���hI鱩@P�E��קcfB�,�0(�8N�5g�Dև"����oqZ��u�������s �>�Mdm�n%�gT�x�~��d���<Z���(1/������ǌ
O	sB���x��\8�j������t���@^�;�q� �����П�Ϭ�O�#ӏa	4$~��A��@�W��i���u��Y��'dל�Q�f�CF�%S�?�lgz��˗.w9��k��������%�=���I�bpL�9&�����;�D쪨D�h?]���8����(�uq,J���PLL�iv)^rҨ�5BS$my��U���lr���RJ{�1���ʷ�H��A@���!�?!R��Y_B�����""��:���X�읅DCH'�
 $N��Y^�V��*�}������lo~�RZ/���aL�h��W1�0���Y;[���>�����eZ�`�����<��_d���]u𳷅�� _����nrl�H)3��h+���fz�0�q�k-�٦0{�����A�f�Œ0�G���KƳ����&rh��� �OZްf���@Y+��{��5�HZ����_���J���d�4���E ��=ׂ�B��*
H�ħ�Ͳ��Ή�N_{kz�V���b�-���]�[_�@�3�j��>=t'�Ю{���2����Ѐ�=�5j�ƉrMq[~�nt�Ӈ���Ꮷ�@�)��������UR�jC6���q���%m��A��Oc(تp}�]x>�o}�������bx�a@2���$�\�xQ~��fZ_N��n�S0��%�T�&;#@)9d�v~;�l
N�Eg�s���3�v�q%j�\�!,.�g��!��)"I�,� ���jS�����U	���8��Y8�����RB�,;�I����gfjOX��Zy���J�]8��kЇ��SKܲ',�.W ���� �r�"2�A|b��^���(���P;����;��¾�k����������$����Z�Q����������������\fӂԋ�1)�[y�?��:��=����|2|�a9�=��,`������V�6۷�b+A�tԂ=�B_�D����N�����v��7L/"�"7/2Pb�����U~!�\s&�AE�-�>�P"�طP��cP�3�{��'�)%D��N��.,�~�@!�������GA朝R����{�/��~(�k���F9�,7�^!��7c�����'�2�@�����:��w.�c��-�~�7M��$��'���Jv����3�T��>�bZ�w�O!z��K9+���83x'���PN�p`�Ck1�J��>/��D�<�/��]�/ݗW3�YB�y��|8��W��)�9�� �u�`l���(0�qZ��Y�1��A�+g� 9�
	����xp��)�>���r"�[E����?�Ћ�y�=�y�Y5)ԂDqX��I��EG/J�#�Fy�M��Q���	������Q|��p^7�y���<�
��~�~���k�z/��b[���m�ˑjX�S�r'�&�/2�Q�&��=��#�#�]O�E��E1B��؇gbF������X:4b��PKt�w����f<�t�p�:����ؑ�N��F�����9����C9=.l�/8\f�m&�;K!�l�Ka�����q�>����W�>X�_��Ɋ�^����Q49Ɔ3|�M�y�H�)����av��C~�)K�G���Y8��E�{�}�F���iD��V)���H��q��+E�	�զ��A�j<D�91fic����|4o4�jr|~��rR�M�x�={�/W�3�X�Ϋ���ɵX�N@��m<���.�ck�ܡf�����[�-�!3кbV��}`�J���k��*��m%c6@�i|qk�l0�Ǟ&:���]�᯷�-�cF�TΣ�=x
R���U�VF��R���<X=���<��sÖ�o���>J-C`�%�fe�:� 1e0�����XBq���t^�`�&�E˻f�ko��	6?�C���,�'��(P�Y&���\s�ғ�+Ci��_�m]�lc�M��C���j7FzV�9�v雚����g�fâ�G1v��C����9��C��rC0��BU4v�}0��E�A�En���?1�%�s=�������s�wxYd��`��\�S-�"���C33܎έ	��ڇb���A{z�ʥ_�WS�$p�Z!�D+�3� ܄Z��Qݱ��x� 4ކlgMo����]ɮ��a��������?��6�ތ�Sw�$\|zU(5gR����)F�^����d�+ly���h�ދ��u�2N�.����:1=]&�oY7��#>�Z�����^Q�Dz���Ah��),F��	3A`�.���u؀J��T�e�-�^kN���f����?��T��U˹7�.�'�m�5�g�ޓk;>K�OBa���p,dy�r�W߾�ou��3��|=����}���K�ma��ۚ��
+�.��-*pEm<�m���]�6^�3�.�}<{Apl�k"ΦH&HO��8@���Π�.u�4^Ǔ��? H�������R�"�n��ׁu���|C�
���D�=ͱ��\o�j!��>�yJ�&@w��%iVۭ}����:t�U�AǷ�h�Ӥ�������T$!��$ܭtSǋR��83(y�3\�����7�Ĵ�x���P��2$۵֠ӵD?=>�"r��`K������� ���Z��tVm�;��iQ��+�F��6C�j��ŘW�f���|�q�&�?�z��0"8(̃���U�+P#d�,Y[�G�UF��ٺK�Jc��0rt��j�����C��0�V���^�,�.$k���O �pH=剸�rF�|>�P*�-�j�){��?AM�9�]���Ne�G����AnP����� 5�D��8}8_�Z%�;5��%;9,��nq��av3���]���������I*9;}|�a9�%�g��5*�_�@�Sξ�t}�堀Qc�X�q��ԗg��k|�]*p���$�˦,�M(��0�D�c���t��g��l=�<9g�,zC�����Z/���80���r�x���}}����E��_a�i�k���kH[�f�J�:[�-�Mwu�B�� ���JA0�*[�fJ���)�m���b�)�������p_�7_�*��۲�"���*F��d�-o�ʆ�u��H˿`��1Zk����W���P�)�
1���a��[4۰�_���)��@(�S���ߵ2m��f�$h�Ώ~�������	�Z;���G�5��iSu��?�0�ꆇ�'�v������H��p4# e[�.�9�m�m���X��~�o�삹�J�G�A`�ѿC�	�Xf����S~�%��J�ʒ�Q�o�S�2m���b��C�[�;E{��m�~�9��<��r!�`H�5I�<N#|��v~Ƙ��a��^� n�m����ONR�Cg�E9�7&ؽ�03�؊cN9���u#K�CiU��|�� ĝ�޶�0ă+�:����߿Ξ4�+�{����`'N�E-d
iyz����h)�/�n�a��s�SD����lp7k�2��6��5�C�~4^�5��޵����P ��K7ۣ�#M�Q�\1�ض��5���x�s��=)�+����@q�ѯ�D-�?¾�SB�� ��+�3�Б��'Ֆ�)\(�7�)���'�<S��A
ee�L�W�'v(�QO�RaK�	wwJ+; u��A�r)ս#�q�$�E���N��3�ټ|,���ʤ1G��@֗
ȱ��c�v��]:~��@Q.=��t�+?���D$�_����*{�
]�A�E[zT�4Z��!sk�7*��(��x��畊��"�q��򜩤��M��p��xD1�߿p�]A�}8��o�ѧ�OG�U�6�����/��E]�#�	������*G_h4���0�Lw�x
pőt��;- �p�����/ej�$b�Pd��}eG´��7���R���'��FүT��5x0���<dQ��9�nxW]
����=�7��r�`�=�\����,�p|�k�>��cݥ֎�X�z1z� =Z�؀�f�~"��ڵ��ux��Ȇ�?��"e���ax�j��?��rȋ��W�L.���L�Ro��Q�?[���.�*3�A�+����.a���߫ǿ�ۈ�YZ9�j(СZ���蘜�-�Vyq�����(��8�7���p��Љ�|�k�u6h\}�/���ho���|�e|�æ�P�WSP8���dv*�U��G�H����	������h�sLA�8�P�rJ��}��l��X���=�)Ü�?��M�q����10�
�u�p^�V ��L_�X/H�Nf��ʥ�;���/�&�WD���������Td�h͟1o��pk��p�u��8�R�� ��H&^�8u��Ӝ�7% <�E�O��y��	�5�~胏�3�Lܴ���eȩ�">���'wf,&� �f�B�l&�d�zV�9
��A�o���E�M���?Ȃj��Zn����s1�m��5	���T� 4����;�_wuQS�$�g(��N7s/�(�4䀥^�d&���6�}�#X PA���ⶽ����3�1(����K��gF��e���0��rp��qE�t�3E7�-���d��v�Z}�!&����aN;3��k�\/q�IS���~��4�����J�ф4�T<�w�A�Q�+Uŧ�E_x�"w�S�#q^���[�j��>=�B��v�EVhɢ9=��HrJi�)�0���C�B8��s	-�Z��7v?��v�����92�nE��]&w��Oq�J��%5i���<Nи��8��x����d4r��#����T���ɍñ���o,��.��4|�V���"J��������k�\�_�OA�/�m�)wK��otLU����&q���">5��n�yq�v�`��Ih1�-.  �M�s`+Y�u�O�>M�'���yrj��#����W:��wb������w�}m;�>q������B�{V�Hڙ\9��P��'n�m`�l�8f���2�������nz�ө�+��T����(�NA誵Gg�n��$�9�e����o���o��"v�kɫd�r_�6v�����j���n�I��~UvN�����=,Co��wB�_r[a�Z����j��[���qH㮠���Ǝ�懃��{/�/�:�J��H/;틲��&��%yE�~L�n;��s�d['G_�E�<��:�F�l����e�6��y���a;��Y���U��\ˋ_[(�9e�ڬ��U�o^�+���C�H��_�y��M
�Z3�m���'����o=1�����A�]u��A�ʣTS��Z�����F�y橓q�,��q�k ͛|������Y$c��c1�G��yqZ�T�[n�+ �tG���L�_j�sQ\�i
���Rs�~W�G_�:�L�y���R�;���)��S�-�M����U�I����)c3���c_c�_�jz�r���9ӑֲnm2���8_G����!�3� G�a3�A�e0f�a�^�p�z��kڼ�2~ml�J�(\݅��ҍ���%=wտ��=<�%:Y������^�xJj���m]�A�>���ތMR�	�����?e����������5�s,0�4���t-
�3�_u���B�ܲ�����T�;���+�
��f�����2��M]d`��g7�*z{��z�4�+\!�K����0_�i����Hƴ�pH�3΂j�S����!D���g<���b�ɘ�4��݉H� ldl������88ҵq�]�	\A=O̓"׋��CD�֖5��t���d��*�_�r�R�K�}`�o�'+M/��w8�����l��[���nЯ96"����t^'���&<�l�CYHcwãj���*U~Py���V�Ht��h�-W��0�aS�Z��3ځ��5L�^\��NF�M�ܥzס/v8�]ؕ�t���u���?)���5|�m���:���̓� �4{�:mX�cB�����u�� �mIE��}m�m��6b��4�w��3�O�#:�{eg;�+�<9�{����U��|##��J��~��k>[�1Eb۰QC�4�;h_C�6H�9d� %�E�i��	G�C�MG
V�'���F�A���ۗ�za����й��Xuw� Wdm�)���]xe�ֆ;h|�0�a�h��D|�џչ4D�'�]�^��
)���&Gm���L�	�s� OWC�����	c�{d����V��R�Eߚk<�v����T=*L�`s�	X_�S�b��`-�ۍ׻uh��7�f��57N�j�WQ���	r�2��C��H����� X��~V
�@�N�9�)Ѩ�i���	[lX�5�P��>����XȺ���;@q�u(�7U��1'���3�,�����Ԗ-��^��ҵ�#	xŚS��"�������*�8����A�X�h+M��7$2/�.�#㻦�9����vb󰳆Yg8mq���8�c$R$����П굚�I_�vܪ�;���p��e�ږ�}� �Df�u���
�N|_�U��{8��DiPXa��fHd) ��d��a�vL/�t�m��e\�U#�s
i`"z�Q��$D��g��k�A1 n�
���|�W�T���jC�b��f~�H��_Z��6�"o�D�ڙ��^9�(� g>�����<���x}y|�xZ���+���Y�'ɂZ��#�f�����5Q��受�:H`�&��z� ��~0���t�v��Y�GW�uuYҼtG)���.S��C1�<'j��_�]B�!��Vm,C�~��T�o��b�Q�+/����7h�3��g|��)�o�#��<�¤��V�{��3�F�wQ�ʧJ%"��gA��2�ǎ��&_[�)�x�� ����E���~$\G�+|nc�NՖʴN7�CF��͔� r��YvY�)�PV�S�cE�kP=�g�$��#���k|S�P���Rk�,�A֛�J̚�F�(�����5�I��l�x��-�V��L�q��R^3�`�3��_\T-Z�vԭY�q����q1��i�|[S�ٵk��}x�#q�q'�6s�\�c-��nW�g;NW�d	:�`�;y��xRP��xH�ʌ%��/���x���}������4�	E�;V�8df�k����L�:M~e�dv"�0��$��6�.�P����� 5a�/$�}#[7�w<fqb�]��cփ�6�uP"���h�[���ٽ%x���W\������N��ޕz�Z���7}�
�����S�w�
%�䴮�S\�<~������V���;f�c����wk�s��i�#{��x�G���)�S��o6;I�/*x:f�?W�ޗ�,�����Q��[��]EL!�]��:�Ǩ�`DZI\
:��ĉ[��c��D��:�.�_ۤ`ᚴ�z!mx^���)�I ���������3�G9�Mr@]�Ũ�q!Rp�Y�������*�d�_OY�(�)&�XJDUH�DL���O���t�{cB�D��$Ry
�a�-����,:���}� gsƴ��k�+K�m���=m��m��`�%f���~��,�	bx�wyh$D���`���(_n%���Q�lG�+i�uJ.�i-�-�'���d�B�}��D���%&��##�b��~5.�$i��Sv��)B��"R��
:`�+$l|$S��M����y �y�
5��X
,Ia�|A=�M�`5ۦx��z�jM_{�0��Jy�F��b=cU���-UK�f��x�ə��/G�.�6ՎQ������4m���e��YL'�b�3�M�gk��.6��ef�){���W�@T�o�Y��f6�* Zx}
&��YfZC��-�ݖ�5O;�*�!�9�*����IY�t�\4�y�(�P��/��*&�$&��
���X� 1����$�� �A���4?j'��]V^�DZ�7��&��1���"�u�}��{8�$�4�m�"����Dʄe ���C�S+����8^����f�P��)�FU�,�-2��d�&q������>2}����:$%��d�/:{�-m`�Ղj�E0�e0���T��o^����/P����/����[2O-d<�q�b0
��&������_q�6�hO�m�����I��d ;��+��d�
�>;���A+�+�%��}�+>J2�J�NL�×V�]��+`F�����5zx���í2��Y�@�T��x�u��-�t�S�aO!�9!��;IZ��	r��D�U��>\��$�Rx��:��,�~n��?Ė	��13�Kv}����6o�K�Nv$�s�B�����E�O��G�!.}����f�57ph��Z�X�C{?*60�* w(�P��z`�����p�{����Q^'=��kF�M�d�T���1G��!�����R��~�cR��]��r����V��/ʝ�j�qfX�Բs.�c��8�)�v�9�g�>j����!~\,�u�m�u�CធQƾצzop���2M*g���5�\h�R���5�N��L��ᤤ���������+���2�����I��˓���g�9��3e��H�������e��4��F�?�$N��f����|sZZ��&�sv��U��GF#��I	�����mv�@� �9@��u �y�a�5��ߔ�� ��ѱ�&iZ��h[xد��w�����l7��r�s���e�V�����.���DD"�J�C���/%"9�P�(��7!��, 5Ka4��v^I'%��������t�77�ri��n+���?B�8�����^��g�I2꤯`�waJ��L	�."'�!����'��NHIaq%�&��z]�_��	�^��}I]��p�ik�]��Ҳ*;�zE�ߋ�PȾf�ps��J�@�o�5�f�GV���C�wjT�vY��MIl�5C��^f�:�	�rC2a��iȃ���Ƒ��}V�:����۰�Ȫw�nU�41Z��w���=М�'�\BT�.���7�u|�q��T`_����J����)!��臞f?&�F����M���Jf�δ>�]���l�%���9�&�o�е�8I2�-w���c����+CC'�'s鷮�d������>��`:������rը�I�Z.JR��P�BMJ�­3S��DE��ݝP�Y���Ⱥ�����2���4�DS�G�f��="�"6k�#���cٻ܌ͫꎄ�¬�����a;��*�e��dzA״�/r�1Ov;(���5Cl�[�s�-ǲ #�y&/�8k܉u���@W. Z�5�V�o�m���l�4�|��H���[� K@�$b|�\h�]~�G�((c�.�؇�9c:0�!���Xk�h�YL�!�Zs�o��+/�hd��Mi��&Gh)����	�kń�^�����u��$�gt��+H���jڏcj���&��Uw��)p)��ku�]�A��g�����p�#\3|Zп��q�cf�F�\L<;���+D�|�AE�d'�}��{�H�z��b��\X��K^"7�>R<�۱�q&�o@�S�eq��0�,�����3����N)�u2�UD,������;�+�Yl�W�Q�;�݄vX|�F5Z�Lyt,�NJ���u<��-�d�o��Jil�J#�'�|�׸�l�]G��}DS��+>��<�%M�J���b[O��[S7|d:p[�V�5;�����^a�7niߡs�&e��#~�0��k3��$�z.6L�a�z����eEY����v�jI�Mf%�y�4O�c�/Zj�-&������~�F_��g
�&� ��.���*�̐c[raX%U��̎���_a1�o6?9M�����	(���m�B