��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�/R�ؙ��a8E?	[��C��|_EM!���MP��� �R.Cw�j-1�,?���Mׄ��E��T��� IZ$\��h��I�d���cL�mG }������3���@T�G*C��'���"t�a�3kM�����p�s��7�Q�0�[0�yS-*e��۞�`4�,u H��{�k�p	O-O���I\��vC&�] �oV�T"f��.�=�-ԙ�v��vd��__)��#� !�z~A�]�=^�O��@�;:uu���B&uR)L'w��c�N�DC)�-�cLF��wc�k)�(�z{K�����V�N�[a�PDr��������:�v����/�3=�aF,�{�&�"�v|����g�O;���|����[2��;Rؙs�l���,��U�d:�[�W��<ߴ�<*1��/�x��Rm��/�G��&�0�337�x�L.��~n�"�kaPI��?�ɼ���a��q���9GDwG�d�V_�BB��Ì�+��wǰ!��D�K���e�A.��� ��8:�1��5`��{�At�;����^[.X��Mdύ����1�a�wk� ���oW�.a&�����3��!Ǝ�_���/j�/�.��f����f"dK^�4&�9/._��F�Zu/��ʲ����H��}������ܒ�ǆ�Q��pli��~�e}��cS��*���#�Ax�/���� ��ݔ�#�̅z�p\(�������l2�ަ�o���ǕsM��#�iR��z-��i��H�8ݥ�*#-덳��W66�3���C=�I��/柂hd�����-z���������*����?s+��{D�0X0����K���ȗ�]��|�j1>��gM���B#��$��8VY�q�?/W����ȵ��+vrn'��A���z�ϖnq���?�L�_��J��'�Z�i='POP�WК�#�"6�E��ߏ4��Kk�r[��QcR��=�z�k��ӳw���@��d��s��.�1�A�� ���|����0�a)x/Y��x�S�S��Ya/�$�T����>2@_ Eq�7y~��Cvmn�?IPǾμ���Ӿ [������rU�����m]r��a,M4Z��#m����M�1;PK��0��Q
$<A�_0�Z֕`��^�B:|cY���t[� C��ENĔ���`WB�]~���:>x��ݝ�P�Gٙ�s���/�����HәL,9��r⼲I�`���8�۬�D��%º_�����-t����d��*LQb����	K���]��f F)aAvB��M�C��I�b���!N�>"�{B��)d�ѷ�������{^K�d�ܣm�"o��yR���+8�ݪ��Ld�$!��)�8���?�^�I�q�X?a_�U.{�e����k�@�����v\q��}�N����	݊3�p7e���g���τWc��`,�v�e'���B��~���?cI>�zR���t|�j�� ��T���*-�k��k�Y)��_�� "�kc�� !������I�����E��]Z�煫��=�'��~�ۗ�3vKr}�p<����w襥��Da�%�4S�UV�W��'�e�ƎQ�$��a6� ��_��K���C٢�4�.�To ���	�f�̔�9�����Ɣ�h����F����@
����>�u!�5�>ٿ�!j������(��%�A�{��R�I����g����fņL���[�#Ǩ& ! ٯI�":~Ո]~6�=VO����Ų��2��Fz2�C�����{l\4:cߐ�ቍ�M��v����Cͯ�]D�^�=e5�<]R�K9�L�	�0P��߰]ű��T�O����r�5�B��̝L�h�jW�����*��7a�MT���قv97��+J�"�
ϕ�D������:p�AO0���� mY��A��w(,sj�*��Jh#um�}wz4�2@�|kW|��a�A~l�T��U=�j�,ݭ�Ϟ�.E��iԹ'ѣդ�?X��ЗBA�O����}UXv��J��A&o7���:L�/e?�J��Z��v�a����2i��]Jg%���u��{�E@�dJ��Aa1�eR����"P~��g��U�Nyz�t3X�Y�؆Ef̵����ǖ��Q�X�{A��:+��p��LD���i��bJ.3Չ��P�����F\V[ة����ʂż~�Im �I�@�����f%� ���7�p�	���x'��E��9���Ќ"9>J}Q���ea��C�o�̉O� �mO�<6�jy���W�����o�2T6\�0����`�i.2f�zܖ��� &l(n��I� t4�O>k�?g��[@敘Z?�v&.�)�&އ�p��O�W��Կ�W���2Wg�Ƕ׵I��,RΆ��ԞApa	8��34��'����G&���%� ��]�M�l��[��Joc�X.�f���g�d����(���~��������� �^��0$r*/�ӂ>�����c����c+��͹�k�@���[��~zL�~�����h�������
�H�ޞ��,�\p��@���~�S���IgA����0b�/Z��=�ݒ|��\x5�C���-�	GnQ��"a��2:xE����/{& H�o�;|@A��Jx��,��g��Y�0 EH�b=ƯN服����h6y:����fN�:�*��y��|F����@?��s��t�5�qV�,G*�u�%!��c�'����KYݔ�rd�2��{�Jy3Tn �G٫^ms��\�S�!�Q8P�j��UV�ZGI-�,b6�n �|miא���R:e�� �\��)�/?B�{��o�y��p�`"�&Ǵ9O<BK#5q �E?HFE{w����h�ޫS�ڻL���G.wSvh-�5�j��!�f�,N�T����*/En����@�(�4jk�Y�`��b��r�8<͂ᷕ�<޹�য়a��j�6��(q#0��	��X�63 ->(�>B�y 9�J>Q�5��s�D��>�m�{ԩҒ����$�>}=R� CP�o��(X��=�����ԗåp�4��3�Xr�d�1��- a��n��?۳�0h���9�f�-����N� ��!�UB\$���'�b9� ���3��p�Y��O��qj�QK0{�ic��L�c���`p|�4�A�
���'��bi��� a�X���\BȈ6#�[�=��y�͘ޠUͤ�t+!$bi���:
�da'�݆�k��`v
�D�!��?�d�<W��T` ]��z1,KZ?�/%�ZPOB�Ϝ��ZUX,E{�*3�V6���HM���/�M�ڍ������l�N,�OP=u�� c��̰G;hxz|��������ڻ���e�BiX�$��lI���r�2����P�\U@�u�qu��Gc:�"��ǀ�%�M��==K�����!9\�۶�@/^J$s�⪺�Č8�wP�������0�r�e�'�w��;[h�g6�����X��33�ƛ��������}���\.�i�/��.T�*�A��o)p@�y���(a���?��ό��g�O���9?M����<�k�I��Q:�щt���6}���~s����r���u����C��T����S/��n��OAˇ8��]7�w��V����ѵk\����~xW���$�!'�
l�b��TH���ͯ��Ʒ[j����w&�A7��=m�� vT���R:�z�"�C������t���:���؞�j|�8�~����FX��:nP���7^V�"�.�T�+��&y��O&1��:̜DI���	����������N�r���0���H~^4�Kg>�R$!��������'�;h�����w�P0d����Ɛ�9+(�Y7,W��yJ��-�	�U�2#5����7�:��ɸ����0�w��B�y_���[�-��d���'��Lp��8�����	�i�;>5Y�%>�k`řz#����l=Z��,��ԭAa�S�Q��`�c�d�&Kx�q�"��=V�զV��}9����$:��86�}�  �
�|U�R�uH\U7go ��]�G��]���B��j]���Xi�)����;5�7�����҄��g# b��gW�&�DM��)g���W�z�ll��"],��q��>����K$=�a<��T�-���{�xHU���pη��_
U�r�b�%�i�[?��MJ�#V�����>m���F�J�7��)�-�L�N���F$���b��8QL[#Q�7�Y,�J�ҸK����
�a�Z�W�"I�Ur:	"����u���ԥ��ID+��!�[�U��%Q�Y�؉�l�W��<�fH����z
-��)�n�NWh�ѤDc�9&�'���-f�� d(�r|j��*h�^�Eު�!���G���b�HD�h�Y(:U�`*�x�y[	���-f��=�l�������DH}���Gf���rm`����?��ó���S��^�[ߐ��5�'����G���;�j��TFIn�������Q���ٲQ"<���[h�W�u,�沜Go��r�vR@֢!V4;��/�w��� ?�2����T8a��m�Lz�	p��iX��:��K���Z	p/�Yf������DL�ww�;X|�c�$�3��aX_B9f
{!(A\K���
�d�J��Q�i�҈�Y-3ɸ<��?>�B9`}X�sP���N�q+���Nӛq�E9y:hE;R8�3Mn(m$�Q<��d��:O�D�T'�/�X.а�u 5^j���A��{���E�W�+�.�dgGB���Cw���/��`�N4
��Ϫ5J����E蜹�P�"�L���&�1�o�S�`i{R��N�A�Sb�C�Y�	���4�3�5�+��(���C���g*)"�*��Q,�X�鶲�Y���iM��@�
�Y?%�Ѷ@��+���c9!��_ ��'��u�ր��GW2�%@�D�hm|dI�E_z�?.CVγ�Yu�u�.��p[z��[��8e+:j	�^?�W^D8��T��"��Ȣ4ӯ�o܇�91��
=$��,#&�{�&�wU�а�z̜�\H�� ��b�s����|a�csDY"y����ˈ�e�m���:h�vUkE�I9ƕ:[��?7��Lt.] ��0pZV����	Կa��-��W�h(.���w�^y�4sI��P!����e�X"K��
hA{Q#�I�f��?K���5̿X|�Hu׆Es�Xk]����ӧ)V)»6�핽��PT=��tj/ë���L��@x��00����3��:}=K�?� 7R�,X���K�+3>��ؖA�u>�ǽ�M���
�C;͐���m"_��64��Gر�M��d�j�U��h�?�#���(;U��GzD[���\0��U���랥���1���e�|�&2N�U<-.�_Qq�[�o��_�lJWE����t`�Op��ta\��o���u��K�@޶_�৥�����=���%> @ĀFhie5��Ck�C��f#�m�E�=����#/(}�?�E�}�W��n$�\V'�$���$�<�4]j�:�9U�q[ȳ	5��p�*��kV�w��#�Z�=l9|:�xc%�=�	~�i&~�Qo���Pӹ��q�JeOy0��I��[ǀ�0��Ih������]}nt"h�G��|s�G�����l&�S 1�@�q�`:	4{�~�E��$l��j��Y:��7��|ch���E����˔�rx����	�6��K��|�\:|:�#e��qVb;�}�W��ɉ�=�vy��y��,����[y�*<>u�"޴&.�s�תT�NX����mc4�.��U㕤���R�#�M?{�kJ'����P0{�3��P'���8�\"^uv�b�y$�vN����*��W۶O��v���7��n����D���05���0CUǿ�k�i����q�;-9cu��]v�Om&K���&�̸�������nQ��Z,���i� ��y���3����d��&2��4bQ���_AF�0��u�B��p[=i������>fD0hڼ_�XeW��$v�}�`;�����^L�Y�<�da���Ұ���o��ˣpph�������QСo�f�u�`W�������8}�@+��	13���A�s�����k��M1����W��#N��JZ8G����(��d�
@�0���~?D�k T�U՟!P3�����1�}oJ��؈9zo��u��Э��/#��͊
�\�C�����h6� iӶ�K'E2��1�7�9(1r�eڻ-�Z���&q*�b_2���T�K9'HK����rGv�����J��7�o�N�-������W���E"�-'�:Qƍ��ꩁ_;6�t� �Q�Ylſ	tGMYK&����\�y49���4���P���d��R�a���S����Br⬵ݼ+�Jݮ~��2�_�^bi��|�e�D5���X�ʢMy`���k���[i$�a22�n�}�=/���Q$�)��e���A���Y:.�6���u�.��Ӭ�ѬU퐺�)��S4䯽 ��޴�[���z+�� ۳W9��l�eF�p+%�}�v��P=客��f&�v����g؇���MR�0�G����or�O�EB��T��ڑ�EX&O�-rs��!�"䮽!�D�+��\˚8���N�۵�=�T�����E�}]�a4m(ɩo#v�Ӎ�1%u9}s����J�uN[�$��'`��$g�D����! �k(��|�Q,A[5��0�����gg lH픵ܕ'6k� ��<��2�̣Ҹ�D=jH�>�&]X	d�j�p�6$�f^���Rk���<&H"Z}�!a|2ky�þ1���v�%\� ]��u-D.����D�%�' a�2��Vn�����Q5�u�Q�6\M����w���ET�cq�������0�]P9d3(��]7��z+U�>Jm?��8�^׳p�|s	�H/n�:��e~o��R����٥��+l��!Ob��` �٢�K/�蓫/�MN�a����J\��-��]����ox2����uZ�fM磹����m�O:�٭O�H��zn^�D�� Hw{����}p��c�����	�%ͦ�b�j/�6���0�k��|�,=rx�t����,W#�s�b�A)�+ȸ�K�JLd/<r�A5N��jV���~����E'����w�,��Si(J-��rAh��fp��Դ~SeY�7��k����-���'�nT�1��Ӻ�u2��Đ�1�FJ��ӵڗ��U������a�sy`��x�)Gu�n�#6�W�"*��5��������)dg�7S���֖�U���ý�� �Q�4�cM����{/HIo��'���i������P %��u!|	���˼Tt�GR��:s�9s	=�I�\� �^�a��ۓ�&��v8�a�4��s
��Qp3���`�3�l;���	���%6µr�l�D��&��k��q�̻�l>�ՕJ�,3�
X�u��[=��@2	{F��8�N��0�$��d1&���sT�/Y�*pdk���3ZdFI�J̑zD��}j�K`GQ]�(��2�%��y�Gc��|�hH������?n�ͩ�$�/f�Ӧqa�3Yf��x��̥�z���EP��i�����6ӕ3o6j0;lwϼ�3]��G�[�'�m��*��7�]���t�%��%�~3[�8�7uO�D��*QXAQH�!��,j����;��a��o��?����AK��f��O3��pQ<�a3A5\����x�UC�*�ҍ���5�5�j�C?�Zu���`��$�GuV�#E5�(���Er�ÄV��6�3�z��j�OQ��ω��J��]V%/�2��S��p��P���v����YN0?�4��n	���8@�eB4�<�%�y���5��M�8�bo���E�[�sx�,�pN0x�s�������Q����xR����{.l��0<(�T7�����$@�p��K��#�U6?=K���i)3m�;�:�0��W>jQԃ>��O8�p�:;�����~(Jj�p ׼)g��֒��H�T���!T�F�X�Ɇ�:4�:��;��T���֋\� w:Ir�}D�]j	?�?��Oгe�Yė�b��Ri���fM9�Áϫ����$���������]H.R�P<�z����r�u���NO�C�%�������Qb�Ei�:Z~�{;��C�����G��Iv��7�T6����d��x�7� ���%$ʉLs��0x�����HK�A��Y� t���6�]B��GUEn�e�>,�)������ip�=ᄘܼ��v�����5D����1�li�����H��4�H�UEF/(,��t�W��2��$++"����ш� ���4��ZHɡ|����^fc���kz��f����뉙Uj��"֒tN6�4g���U̘Ž�V:���}�ѽaH��0���4�%�C��(�zޠ�Ş\�}`�M�d�U�g�6	C����� ��}ϔ�����3��9�����b+�H����6\V����-��0�B��CP|^�P_܃�^��9��DY0��$�CGx]Q�V
���V��&��j^(���Sym��^ȫL:1�% J8\�5~cbs�b�������q���y���8R/�u	1C"�˵Wᶓ��BK����)(f��s�(�04�${���h"��3 �X������R�Ӧ���R�o��5���ۚ����!�W����<n�R������\�ֈGS�	�ɢZU�zu�J���@��v'���ͯ�	�����L�b�+�7?pT��&s=l�}�k���JHx������	6n�%�GQ�M&yIbf�
<��y�	*���Հ�@� �nz����ȴ��?�X��c_5R}*��w:tQ���,�2R�����u^�0&)�?�����&c�Y�K�=GM$Mh:��}���p}Aj�j\���S��g�R�=���V@ەo8�+�	���R��
3彇>�Q��� ��bt�z��T�KM�x�nm)������������)�XMI!��~NN)q,��,� ��?��D����(��[��7��pڔ����F2�mwĞ��E֚��WϚr�9�SJ��\�A�u� ]�����6�R��V�x� ��LrF�U��S�y����������9���ɗ�qvY�'-Ңu-`
�\�.B�?���qpJv��\��k�Fb����]�"��]ӷ*��������B���b'���%������^ئ�!��3���i����?���
4�5��s��j�n�� �S���ΡǊKo!��_����2�QPˑa�)�z�ñE��(�9#�MI���(E.�N�j�Q$�Y:v�mM1ȓ��VO4�kE�dd�L)�?k��D��@� �
l�Du�D]���']I��E�g��-"K��/k���4�.\O1}yR�s�;�*���u���k]�d<�_"�6*����S�ԈA�+�ҕ�QÈe��m�5=��u�/	��N�a(`�y��,����m��%�<�9&� 6�@�,���g�sx|@��� ���B��'A5NhU%k�(�����.���ĝ_�Q�dr��������(�Y�4Y��=����7} �/�i�w��J�W�A&���%A��4Y;s������ klt��e^��H�+�������\gE�~����Z�˗�5�ߛ���
ތh�9[��`׍C����w�����:�fr�g�GH�.�I��p�ф����sS2�=(���2/'*��_�H�m��X���R���J�3=�H���s���W�7���>��'���� ��鞮�f�A���:�3'�E��Y.�es@�HINf�v@<7��?�!5��.ȑDG���S#�Z�-Ym� �ٴ@�G�S�L�Xg��ķv�dq
*mr�3����!k33anB�Ƶ~��S�1��M��r���j[J� �1�b�.%�4fV�ǊYf�_���)�9���`���ꅗ����m���[����i����ט8'�e��D�)��`�_\��&91h�D�WΘoٍ���1_U���I���zI�=�2�Ѧ���8�y�`h������H"����=����YZ�GTZ�M�_V��Q�ݧ1�C7W�)���YƤnd6��>Г"2+�bSq��캾��Zs�EV���0�-@3͊��I���?��,<��x	�r����^<ڈ.��I{i�k����x���vk�+Y�xscQ�` �k��I�c�&�:AwMwf��vC5]�D����3�x�,�y;ã��K�!#8~��>�s�w�+U	=_x�rg"�L�4,��E|�Sءn
�]Ka�<�s�4v�b��X��<��L�}��$�������_�����G0*w�s5]�E:�U 6���{�ԀѠ�a�>�a�>X�36p//e0J���5_F܍w_������<'>��s�n�Q�"�r�h�.9�UN�rQ&v��ʋ4<N�a���2��dܗ�u�8�6v�����p�TK��F��Z�̀z7#�U#r�Yȁ��;�'r�J�8�i�a�'�M���g�������e\�9O(E���hՉ� �Ac�S�	~Λ5���>�W�=s�\���C	�yy�������Q͵����|��Jέ
�Zz[i@@�(T��T� ^b�P�%�C�ۖ�m*mOH��m23�`�r�':u���|��Csnv���̪fi����~&.�s���p��h4��ӫԨ5�,��tc+R�����<��%{ �*���᷆ۜ��Fa�T���E���l���b���n�ENj�tCy�2.��[�`*,��T�A�.Uv;���;�I����c,���E1�#�@�l��I�����Xę*�_�0��h���4�*�0�8{�=+D>�DZ��z���S�M�҈?�����*�چ
�~}����nxɻi�ߵ~*W �~E;墼�����~*�S���vO?�$с���K8�ۉf��;s��$��-i��yS����	U��+|��"*ĸh��+˔�_tؘ�-2�
��[�:.��Ӽ�����������%���q��3�S��<�-{࿶�zc�-�r��-��`r�(g6"z����\����Vfr��}[#����)1�g*�1�٠(A�DY`�Kh%m<�-]|��n�����WH�ۖ��,W2
�����
a5��<�����'�$���r�b�d�ʒK�~u��l��?ߝ�4r�H���M�A�T��k>
�MƆ-|j*kۢ`���}���]L]7�窧�
I\�[�2�p����˜�9�q�q���s��+q� �p!.玒����Ck}#�eiV�@>�?CP���m�$��Tb����M�`����uEQF�)̇?�#����X-��B�A5ZA/o���5*ؘM�%)���J��&7��݇~���4;�M���j��6D�q�� ���A� �]�����<��{�<{4�3�X,*�ͮ��� FSÅ�~<�*S��x���z�N�w������Nc�*�eM�\A��\�'�����W�/��	 ���[[Ժ���q�PFa���o�J;���|�:E��(�a�W�w��%�O"?��<2�5�7�)�s3�����mYJ ]���_
!�P����gC�(��!�i�_�D@c�1~�_Kx�7�AL�R�k��T�V�ٌ��/�DWlȊH�t<�	m5���?�n�C����;`�����2M��!��ղ���]�ޫ��hv@E�*�Z9����ʕ�;;�8�b�\�D�� ���?�2��=z_�t�e3ry��n���!�����x�L�b�-"R��*��>KD"�%�
��藚�.����c�3���A3�N���6 ����i5��n���`V-�T��K�:�̰��������m�8K�����-?�u�Z���+��6�#���RY��(��X%簫�_@1y���K+\I��8��c�3�e�ʁ#d���	�[�w�Q8�܈�n��Q �H�?M�ߙ�w��ݙ�s��C�'�~XF�����Z;y	Z�Sj�h?������\T�~�5�!�I��7\�ch4�|c�.HJR3� �ɮ�8	P��|��� �)t����^�]�,�j��"kx�N�$�h8��sE ;~��6OfF�~T�Xn� �8W�T[�\������`��-?@}�מ��@�≆m@��E�����L�����`�v��s��K�O�᎗���i��V�9�{*d8!� pZ�[t�cҐly8���ЂMQ{�l}�*l3 ��Ƥ����<5�t\�=��/�L�
`i��P!�^�L���wW�:��[�P,��7�1"���𐅨F���F� {��e���{�<��[���t+��T��A}1M48�Fc8���gR�F�����]B��=�Xqr���rKJU|5d@#
�ְ��c��6��L=1hũd���B��@g@Id|z]G��-���c�
�X=b�bAȬɳ�Em�,��](���n�86�Reb�`˚�)wi����@�"�f��A�ׄ���o�E�K�ת��{��b������&�R�'�F��u��E��9u|�h?/���P�i�	�1)k�,������,�"MJq}����J(*�U��r�&0f��v@���o`&���Q��V.^R�g~��ɖ��S"���~��uo�5�#�ҳ)�1B��߶�i�>Dѡ��>~S�i��Y�U������\�����U���* N�,�}i�^�MfE�:��l��ءwK�>���k�?���M�f��O-�W������j����鿮up!Z�Fz�7ϰV]2f��NC�5V~2�ށ*�TO��5�X�YD�G��{�'�c���3����dIP�Q�)���ܲ��`Cqv���Z���\V#{�?-_k�QG"���u�j\\�^M��BGR���o������?+_>�`�|W��}��]	�� �-�Y|tf]$����w�
u�&s��1������L)�P����rk�����L��P���R�M��X��]y�e<!��B��Am�e�m�5Qlm�G����7�;����'[�v2�eg-Kf�(<�v{����1(��Ǜ�Ζ,Ł�+4�����yNG�t�6:v>�ċ�4�?������o���6w���tȒ�Rep��Zz��nN3l(C@�(��2�3E��RF�,|�Z��:���t�����1��=��V�J%�`=&�(} xK�(�/Ե��s�	9A*ɲ���gD�J������oc���N��*��{ �h��{����\`5�M���׼3�=YN��Y��=-�?�ԡ�w g���i��dCL�^A2D��:��Dv��F��x#�1�aH�NW;�\�xBʆ�0�C��g�`�O����&��O4�+��/�?�W��-�O��Z�)���^��:-�����x^�GAZ'����ւ�_��|}l%	9(�4(�:-J%�B24���Z%�`���f�)��O�hC�^/���R�9�*�s�rK_t��Y��/~8^������MĂ2�,z�Z�h���5}��_N����b��x��<�;|�N��ܑimz���u����u0O ��;I��ϭ�z7fA�Y���[.+>01%�T��}�y��:�,?��8cW{퇀�լ��R�boG��	$��ߋ���m�DH���ϜR�p�����$�%�KX�=|W��T�Z/��.�s�Ϛe��~�UB�}J��� ����cnI5�n����t�b��ߟ���qӡHw�P�7���4g]�@��q;̻yr�4�J��#�Z��l0j��a�	;v����>����A�ޗ�.��3�Xq�̤���B�.W��$��
D���1�.�#X����7%�/W���@IF����_N]�G�~Iq��n��N?�K$a>�r�uk�RL�z�DՈ7�*��ur�# ل�W۾�<W�C=�Ģ�5q���j4�ȠO��gut��6)M�����;50��"9�YT�;x.!��Z��#��lp��3u������e�����{�ݗ�� �1��_^��6���W�YDU�����I���mQkk���[D}fc����J}�yAf�&|SRI�R������Gst�l#����c��<��A���~��� \��K�����I)��f�nr�ɴ�XI%�JD���p�kO���o��U.�LuRl�� 㼸"٥>k�������j�J�ʜ�%��VLT}4	����I�Y�б�=KS�GBO�UTd��%?Tw��1Q��B�W1���0��gZk�y�LK�������}��vk%�f�`ԑN̇���0n��)�^QG�L�����i�(��_���U�2���Q
�}/���\��Y�]��c��Q�Ϸ.M��u��E�4�}��5q���2�(����.�"y�-O�AUߗ�q,_oYI�X4�������s����J�e�4����F�~~eLlr��i$.�rK��k��#}C~��1H����{��e���]�/j��L��ǣ����hb�Ŕ|3=Ԙ&�@�E|#E���DV|BG)�$+ټZL�n�q|���e{9�8`K�?�_�A���.yϚ��������Z�=�vSH�N���T'1�]�pn����"T@����c��]0��ngWh�PKS�:z}J�7�/�3�S�;�y&�)I̹���(K@�g�	{��վ��Q?�ޡ��3�|����ߏmT�L�y�s2�I����)�P� �cD�N�sf�mL>������� v��ׇ��0$i�gy�S<�X�iz�V�!��_n�X��������
�O襗�Ĭ��Y��fg�e��	���L�n�SX��m����^���������l�@NC?P������@�d4e�XM_v���䴪eRɩq����Fv90=�'�xi��^����a<$�IA��<�����h G@����k,8y'Φ�Ze�`��?7Y����k��H1�WM�l�D�F�I;�z���������l��WQ���gU���t�@΀?�_���Z�j�)�AYC<�J���|��h�������|W`�� ��dy�o-
���#Mj ���_0�elY�x���W�~��	eTg��O�Y�H_{���!u�y$�H�&��
���T�K��^�����WAL3�c��yh�.����k6��W�B��~X����v�l_��0�]�Ï̥O��p�X�9L�kz'�D�6�V:=t�4�}�t�k�o����A.RQMz�j�Y��0iZ~f6G��8|��W5��Hpfu���x��QMIU�	L2*�&�j ���x��D���S��[�p�ԯ��,�{tQ?nr�~p��-دТ6E�(��2�V|�6���u�����l(�{�w!x}���!G�,m�S\�1�S)?���"��%7^�yJ�-���-�4�:d.3�a�࿎	=%|>w�O˓j���P-�bq�{ωw��>�P����B�|���ض-�{|<-�;���\A�5�ofn�wS���bA��@X��h��Kg��^چ���x.�>j	�F���:�91Ly�?�\�F����J�A���º2�4T�!<'1Um�*mÑ���Y}�Fn�\�R�NAM�V KY��~�!T. [���3�ʉ^�h���Q����LO�4�$�4��
����@��p��vE�@5� ;���vE"�Oq�Ya�T�y ���J�1�;��9Cxpr�r���4H���[�K�;�=̷wT���M��AU�>��y����`P_"b�;}}�a��F��J�j�.C�x���ԍ�0�>�ة�@�wwGxk�z�M��X8�~TgtJ�D%���&�`߷k%w�nex���e���֥.0I���,}B�A©C��e���C|�$����9>ͬ>�Hɪ���	\�)��%�~As�yRY�.���b�l���9Մ�CY~�쩲T(d�y�U�����~�pXP�6$��ւ��j#�R�@^8�@G�����nc�5U�i�+����䦝�P�k����]�4�v�x�	�n*��3��D�I��������ϑ���$���̷b��~���w��Z騂�4�K����2���z\�- ̖MPsU�z��	���;1�Q尻�Ʃ�e�LU ��RG���� Tff�))��3R�oԞ�lʄ�����6K^�`��s�u��k�L������y����u��J�qA�U
9M����$`%Z -1���{g8��8�T��Y!��З���2N�)��
�)�b��U��`䥒�q��0�*��&ώ����.SB��#2:JuدD���u��w$Y�B�Q�	���ȶ���Y�����p��r��*S��?�
��59���Ӿ�lQ\)�m@�"�
¾����6�&��S�=����"���G��]	��V��p��UE�G��w{�xJ��^[�a��#�K�~V�*g�չ�!w�W��^s��O:x`c'[�G�b��+��{��ɚٵ�����0.ȣ2�N�tXѝNc��7�2tz��ZXg�tŰ������h;�>*����e�K�^��E��]�Mq[� �i5����j�#"����¶������(����C=9@�oN)�.Z�7�9Su=Ѝ����$Qr�z~�hf��9��<�
��ؼ����x��M+8�.��CS<��o�9k���?���/�Vh�;"�,����'}�8���*�Yo�.���L�|���eB�|7/H�R� ��A�
|�/=2�f�����?��X��L}$Sq3�<%E�xZ�Z��+�ξp�S.�W�+t�!U�-{Ϥ�� �}�Z�/��7�"�@����:�1���[R�]�,�/�7���Ou�0�c� ��^�YM7�hʣ
}g��[>a�[�ѭ//+�E��l��}��&�]��YT�7c_�j����J>��x�0>�u�%[H�I�������kt��7���J|Ec��'�~XX�� (R�Ot����&�-6|��&��[�c��,YBX���L��f��§�;i��!bk$WS��w�C��q���֖�9�	����ֹ�)Z90O�������dя��o�z�Z?BEx��ze�P�X���Z�;rTL)�|�KYHV�Y��̮�Ք�6��A�B}i��@����M�z:nN��� K�M�j פ�~�w�(f�'�*�^?˽��2�A�E7����l�h��'}`��d�_ �Z��V$�8������Pya��p;�;����o�1���Ju�Fni�0l�D�*3��M�T�En�ϲ��d;ь�崼!��S
���LB�|r��7
�6WE3&� �M��E�fG�X��T���}OA��WԽ7�y�`d� ���~�m2�yS���9�mfB- b��d���Vq�J�0s�g�ͤj�n�^�#��^"o�/��(b��͓�ǃtK}�0OW��;��S,�W�R��U��[�u䦅�3��?l��p�4�ܷ�1�fZ����ѺY���h���'�j8Px_���E�/0�M�F$��:FG��ώ�[淞ͮW�> ^M<O�~X��!Bv��phAǄ/��Z�]�������&BTj��ˮ�I9p4V*N6�Ըz=��Q�'5��\�R�1��>��8���!Id��G��A������W�	i��sz4���RFEX@6��]o�+0z4P��6���0��-Pgz�5(Hw �1�U��q��VL�����
����F=h�Z-�Os<=:�I�t��y-���G&[	��ՔSG�z4��Aq?�k��>jۮ��;�g�Z��Obst'u��a�A�]ꬴ���?f�g��3J�a�U
�mξF��L�
k�;���`�6	y}��m�훌�q"���F���z����9����[ʯy�zb�M6E��M�(�ywro{���b[�RV�[^�bQ�%5�#�����`����۶����y���W���zn�{Se�c�&a�α��q���!U,{�6��38B�x����}��j���t���}HI�s�q��ui���4lr@�\�ki����Ǔ��<[P$�h��4���#´v����ũ���	��|2q��~���6b��f^Y:�����<�ޜ\[�%'�V,�������{�4j}�3���Y�'}9��08v0+LK�氡s���tU�)c�w"ٞ�CE�'sāS�1!������a�/7+E�j��$�]ַ�E�!_����a"�._Y��ν�hl���|�I���I�����lnUNE^t��Ev��W�ֿ���"��3�M��Q�Ze�*^�����-6<
W��.y3�g�2��#Y�I^�b0���wUI-��,�L}�z���h���L��93��W�﹆%�H��d�������V�ve.�eYnR�I��)ܒ�긿+(��7�XwD=�y?�8�ZTWC׸-=�@-���.��[��s�!(R/+�{��>�M ��2�e���<�j˒mFۆ�AH�=��-��~��gσ��V�tNN�.IU�l�
{���s�[����r6�b@>S:�k	�1e �{k���;���O��xؠ�?�R���7�}�ӝ,��K���JW��U���s2���j�����GS(�tU z�Y�e���9�e�����6X;��Z����(���.��>3+oX��4��(L��@��%]�4_����u,v塊��O��R����P���������p����=�t�z_�4ܱj�iL�:�\J,���0� �O�sH6}Y�� �Bo���W�˩�>�<��QV�jłj�d:��"��B[������1nnl�O������quX�;N�������X�>g�,ѹ�Hu�AΆe��.���S�
0�E�Ss�ol���*CԸ� �x�X�bc����V���rAu?��Y{y�;�Z����.�*mHwb���m�p��+BVZ��"�l `�`;��� ��c���	�ٴ���o�e/�ǆ�j�xo��41I�6p�t��a���=��n�ͻ�s���Y>;�V���b��4�
��0�n�n	����D/��un�\ٟ�+�:�r�Z�Zova���[?ƥ���l�`�O.o��8��Ne�ƹ;���ӝ?��b[\���Sܥ��w�u��#�F�����Me�B� �K:;ݗ�$ޚ�T�ͬ��LM�|�!��[�!���RO�� �	�R��5��5iNS���I��@Gg���Ԧ��02fg	���=��4�Z���	��s�:����[r�	W{}��]4+�,smu��:��^��F���;�iȏM� �����W)��UA/&�c!D�������* \�-Q�B3�o!�ϬT���OV�֭���_>i�����JG5������l�Sc�CgF�����`��U�Ҋ��T8u����.",$E$�����/&2��fqazxpZ�-�w�� 7�\b�7�&}�rmd�� Zi��t}�w�H=�@�t!� �L��4
!WΖ���@�+k��	�!�d@���W��l��;+<�䁹K�n�jUн��;/�0��y9r�mƿ8;�O]*��R^"7����D�k?���m���j�VDx���B���W#K�D4����j;�Ħ���r�q�D�N�%I}�Wpc�v��G�É��y�K��^�z����d/LZ��U*�h����k}�Y+Prn0��\!��N�q�+鵡���W�����Y�:�G$�O�,@1|E׷��f�s�=!�T�q�H��,�P݁��Rk�~R����>��ݞAĜm�aP�8ɱ�v65K�M)�[Ե$�>B��SÅ��� ǡ�����*�"q��$�Ѭj�{����f��S@IU��xג����PYJ��5 jVrC��eˤ�wM�0���+��<Y�E������D�����o��YcHd�҃M?(�H�I����Kv�֓�q�[���N-��7�
�}�C3T��J�C����鵪\8鮭��wC`�?�FF�A���Ǜ[�_�~��P̯�� \��Pb���F|'³�Y��֭��p��&���.�U�S���o^�&m�l��G��`]��چ���l�V�U��֩&�z�X� a�Jd��߾0�}Tf����?4�T�ްD:ŧ��9�a�J#>�L�)v�����B���l=B�u���j�'+��'����������C�ؠ�b�U<OW�d���u�p#��Uj"�z��Z]=�BB��L4��t��6mɭMb<7�1h�;���I:�E54	��Q��(�dq�ue �p��[,����r�s�t�a���#�D��Y|����F�@��R���A?� �=�e�D�������9�)q
�h4��`��g/L�P���{w��q�R�d�q�F��y���F���bTbE��hv+�<	&<# �uF�0�^%���<*��	V�?�z��qM���4&T��=k:j,~>'#|��+�)<y�eͥ�E
I��β���1���[9�QT��i�ɋXKfa}��g�#}��!A�����K�&*˷��fď�v��ڇ��t1���<WB����@"����A�h�ֶ uJ�I�{ۛ��_L�'b$�s��}���{��x����"啼�P��zn^~<I����k�֓��`X B,n�H��Y�[��ݦ�Λ2c�n��� }5�\,e��陛�M�%��0�хYī��)�̊9�
��-9�`�b�!�]��W;)�Q@4�B���
�:1�AC�������qD*ˎ�b�Ow*�8,��'��v�&��߁��X�	�%VD�G��˱�S�l����@�8���T��$�o�f2�D����!�o�XP���߼^�t
G���l��Ú�G\t�@�+<�e���[SxW�'��E�H�;���U��
��U2DN� X����8ao�h�p{��b���(e�j��e��2Ǉ(��-O����6 e���X�����,��l��e����O����Glr8V�^�̀"r���%�F�h"��,��f\�}���	Nѱ�����K��-����<�*(SK�,��r[i� �cΐ�"�v���1�.j���u�:��`b���pt3&O�~H"��{S��5k��ηe��L��L-�QV�,��A��s���^�0�Ǐ��[R ٯ|�_βX�;��W��R�Zb�|�C��Tޑ`�9��z>�Feڝ��
��k*�x7�X��9���������c��FEc�������~�������1���z.CiV<�ʆ��T�C�B���Elй�ܙۑj�!�[��Q[C�ڋՑ�9�]ל��ȷl{Ǖ4�_~�uo��a�7p3h��������in矋Il�ߐЋC%�׵��c�$ �����C&]�YLp�)��A��c����-.�k̯)��ͼ�){B̴���>ab��7�R��X`wI����vD4�>I@緱K�!���{=_6fg=l�O���C��EAO,���m�����+��&Bq���&����ߺr|����wIs5.ㅎ:Sl�MXt�)�O?����!Uh����l_4�ƃ�s2|π���Ͱ)�G Ft�%���S�|�c�8�R��l���KY!Ȏ0�j���V�'�"Q�b����,Е��U��ͱ�q�E.�.0
�Ȃ�
��0<��c�ME�Z�:C�X�&d�[F?�B��xZ�Q��4�DV/Wl�}�,���͸�H|�׷IC�Srp���4��lsȥ@~�i�K"R��B�/Ƚ��1�ƻ��%��3绚�-b��*D݇���������m�`�D	�I����6M�;Km%$dj�.��@T���.u�5��3��x��s<���4�t��J���M)?r�������~����#X�=1>r�̈WM#�\U��x{3o�D��~���I���0���7��/�+n.��-K�y����L[��ߥ�lU�f	�orE`��˾�1���IX�v<}yG@�����;��ޘ�Iܕ�!����oG�'{-�ֳe�ˀkl+��:��b  ��H�?�f�'�&��|@�4�O���*K_�1O��|kngRo}u���o��X'��EW��;mІ
��ng��V����,�z�DIAs$A��Pύ=���|=�4�փ�ߕ����u!! ��N B%�C��{�A;��LQ�(N�h�+�l
�)"�2��e���&��	�1m�.,�z���l��I��tj�FW&����	s��y�,1q+��Yi�.dm������xpPQ�l���w�Z�s��.��i�	�;7C>ti!9�Lس�+՜�.�S1���y��i�q:Ć�N����ˏc�m(	�@� ��^3ے�(��ݔtT�X� ��:��ܦk��`Db��G�+p�fˤR+�'Մ�#P�WB�
M�z�K:�����́��`% ��@��㎌��9F�K~`�=��e�8$���ӺܔS�1{@`��:���3F��q�2�y��؜1˛6C��Q�v�~����,��l%{M{iSN~�a�D��"P��\}`b[�|�+̔��+Ab"��}���w�K�J���3�	ou�]�Z�^�p����χ�EnKx���~G��ܖ\��+�F���Z}�I5�.���tJ�������Xl���l����B��f�wץm$�e� ����w�|fL�?[I�:�PGd���f��k��?���S�����*p�2���$lI^y��z�j�'g�G��.� M*|a=�Wn����3T�I޿���x'���9ѲQ��ػ�.�>#����Da���}��#%���P��⤨}�;^ԁ#�ȡ���ޥ���
�I��Ӡf�ʍ^������1���q6Bۢ\��s�>�o�3��.Y��"����>���1%^q�����ީ�ٹs��xI�ܧ��Ѝ�4�s����F�_�Vg�C�Dc��1�D�+�(���F r���O��t0�;��4*+2���|[-��ɰ��Fm�VWO(�(^F�8`��P`�6��GP�=ݍ�S�q���ߥ�b(���TP.&AV8eF�I{�hf������Ep�NK�Z���^��[�ݘ�SFR����pG��%��TO�����F'GA?D1���ւ�|t?b�6������t��FZQ�Z# Vכ����,wV �G����c��U�}��������5����+�UJh�Ek���iJ@]�Ѻ�2���O]E����{C��)Iw(�W"~>[eZ~���"Q	(R9:��=K�\�D����rAg�J�~*���0^F�>f8�1�g�}1w���0L���5��(�'c�v�*���9�rIw��i[i�U����o7xi���ğ NS�<�vEUF ^q�1)��0�ݧr.)�����Yvݽ���B$�����?Cp����Ǌ}�<�m����o+�j2��t�L
�p��k�=���R\w�X	%2��a�oG�C;<�u<����y.uK�i���$ �;���׽�����ǜ�58��=f}�]�݂���	�����2&5�`,��]�b!�V
X:s2��e�B���Z>;�9@�GIA�`Ƽ �&�z���5J}��0gL����@�>�l�`z
�|�6  �����{��enL���/����3�f.�{c�d&�wB%^�$��*�*�H�1J��\������`�GnB.��"�R��'Юܥ������1�����ع]�ʦ�x��n|^!�^��N�-���ȏ�}�t$â�ZYH=����c�4M\I8D�I4޻�A��Ӗi�.��|1	�
'<�	 :���#��˵��ʧ1�[5��M���o���>\߹���0��*��d
h���*/A����<]�'S�]$����SƵ{a|�Z̹L�/�?h��Y�^x՞;`�j'��,g����E�4SύwJq����46�+�o�L��O��W�g�q"T�χ���(�-��A�s���9���O�қ�P��K�k�1���F���>8\�t�A�㲧O�g���eX�"�o��������)q(勻h��E��g �?�T� �L��v���u��JPX �̱�o˥����4@��B��]���T�ud�Pn4f͸���W�|;�&�����Ɣ�o�D�mj��e��j������Fw|+N�JA�NT�q̋ڕ�:VYj�#7���IƿʐR�J0#?�P�w'�'��i�'C�<��B �IuK����L�`���vI�}!�&�|���a�ݽ�/��� S�SA��|�5�<3H=9v߫�E��q!���_״�u�gUQ�&�禀i�oL���_c|�CC���}u:����Z�$Zŋ��ۤ�����N�}h�T��`��D?�%|n�GC�t��L���o�fC�i����L2�<r�����e���
A�~��x�fo9F�s���"FRP+P��KeJ|�P?c:z$_$�=�D����8o���<Ј'�?��\5���=����PZ��6��6bY ����b&�9���e�1
	KЂ~V@W�hS�j�	�(��I��(����"����Ҵ�x�4�EF+�X���Z�U2��=W�}dP���z�Ӟ&2�; �ys���}%�6ȌuCa�(n~NIg��XDGaZF-�O��Vo�HTN��$\�r�"��E�P�Ψ�Z��NPD�U,�X���F7�fD�o���j2�c�;�>���������Ĝ	/�������<�!B�ė��nC`=�u�:�'8�E��~���vK�_D����R�c���q�a���������{C�c�{�M�|����d
���#Cq�G�|�`J�������<qdb�]� �aY0�x����k����U�٧�9�1����jU��j�&��3��Ċo�����݋UZX�鉁��;e�x����Z����@��� 5�����]�-ﱌ`^ݦ\#��wiȴ���)�Į��H�d7J)����[m[����N�GB^H��K����=�"�#���,x뜦/���~�q �	s�uR���2�@�����I&�32W��*�L?�*�A㱡�N��'�#JB*��@8y���ZOl������}co�.�P޽A���M�m����M�Ԓs�\�����h�V� �M@���P5{�rͧE���;�#�ǟ��Z�r�%�}K^y��[��[��sZ��aÛ,J2��{o��.x`��Vc����#��*�͖�������蹭�5>���W�Ts�:�����H1.�0v�l62Q����1;/ �ƞ<�4��k��ț��۴ݙ"#bJuΦ,ݹ����&����-�xB�)�Q�e=��Ђ;eם�uf+5�r��OQY���&��Ux�b �C1��5���˕�ꬂ���ZD�Ջ�Rv&�;7���y �3��. ��r%Tߢ�«����#>�?yO�UV��[�x�`�؃�q�9%��Tf��=8��չ�x1ɍ�����M�A�KF��2��ͫH���
x��:ް������S�^�}>��9k��ՇQ���R��� T�h1��b��!�>$�ϑ-���͖���M��@sfM8�Ya�S=@�q����sw?��ͭOq�I�߶��O?[�-�B�0#6�Ha[��/4�G�F/�l�IW��ҤUo��<qc�����N[��M�[g�y��$g�h�U:XS��,��xi��')
�Y`�O����>�#P�Ҝ�H!�M����n'�'�t��q��L�`��{�4n�S����p���M�=�f�2���Պ"�?fUl ��s \����@㵍��c�*�����v{zxVxӟ\��G�UaH']�0�~0�p�P����.z!mP���Pt.���9h�ў�t���8�-� �	)�{���x2�C��e_����$�+5��խ��qs���!ў2��X&[�<��ELTs�j�ێ�Zd�Xc�^<[��t&g�w�n��},�ިkP�o;* &���Wl�ԍO�V�zpE(p�������
7W�Y2�1̈́C���� @�m�gab��f&�w\�2*��C��C��oFB,)@�gGacF��K)���_�X_��R�O�����`{$v��,M�as�!f��n��-74`ʾ��7���W9& ?�d�����隓 @��,ܳ���)Ԅ��F�1	Ŵ���w`C�щ�\]�B�[IK���S���T�I���r=)tn� ���' �4�k������2�dʲď�1.�ٸ!�@�n�P����W��8�������e�Ep��V~�����	2sxI���g7���z�'9���^[��7�˺��5I�4<&*W� ���*+�tԊ�/ҳ�Υ��`��<�����Z����,_W,����l��/��2;n=FX{j)Ȟb���5�!���Y�Y3lp�N��4i7[S�V����;���*F��I�*a��Z%*^�;�Z?��tj����2B��#�*(�O�8�j�k�f7H@��o�n�ԇ�h�7�RnR304yټ�[�I)�!�䕗��v�/����F��R���"h+�Mwǋ�����d|&�H�Ud�Q%+��nbĩ�C��wF�L�`y	g��qܵ3W�	#�~a��C�"�"Q_��HZ�q��M/����(��.#'dG ������;��-�i��yo�;A'-�/D�P�Yv�w�E��(��T�&ݙ�y��o?|_�g����,[u�'#]�y�tDDdP�b\���Ъ���8�
���������
���d!P�q�ڿeG��r-��{����e}Qsx��mL�U�B]#���hꏐ�i����K4�e,:��*na�7ڂe��(n8O�/�v��,�����So�Z��WO`�;#�zUS�^,�i3F�2�����@n��?��|蚵ᅭ6ȘZ�TظI�]6R��69�^�R��c���IR%���^��YW�+`�$Ք]��K��R&Z����M{w�Rc	SP}\�
@�ǐ�5�vh��Q�;m_�Kb���|�D�E��۩��h��eO_�#���XQ�*7X:ᶞA��]�����``�zfi�]��t�ڻ������SϤ���b����j���3��tt���(
�g���&t���'Ȕ��Ȣ��[^&����4�M��Be����s���2�XVe���?�7�N6��9��ݧ��*�h F���X�؛�m�[b�N�'R��U�:R��S�q;zF����PG3�ک�sC$�L�>ɖf![ɫE�ӯ���7�W�A�P���hv6�לd�B���`$��t6��͍E�O���9\�}���Z2������.l����B�D�����K�a���ޟ�wPd��`~�>�'������½Օ���A���G=ŮL.�SP���Ċh`G�Č@s+�0���-���!�[,
�ŋ�h4c�TҵD�A�r���GV��ڐ�Y¥=������ed��Գct�{9~ٗ, �ZK�G��/�z�Z������?6��	�
�f��8��XEJ#C���Tez�
*/�1�7sS�7��������˦��RCʞ(2�mK�����/�d�XM_[q*o�LD��9��l?:d��ui�q�E��⹣\�;ii�ݬ�� �MԣxY�k	��˲���-��a���`���k��hg��\�P�TUB.��%Sܪ��hB��<Ig��޼�
���R���Uw.I�}'g/�ޒ����������鬫 g���z��P�!KB{��϶��"
0�06���^�h/�)�PQU1��b9�E��>e�V�C��g��=S�A<�xے��X4(�O�f}ܡS���+�}��57�eg|[F�rC���~�t�����m"����:�����=5o��@<l�X��v?��8� T��By��Gɜ3�j\�늶`-�"P���S��3SOl-Șn0���51~a�`C�4:mNr�Ƒs2c����N��L7Q�=�O��@���s!�=��ӓ�QǊ�x����*�e�=�>D���9�rK'8�#��EOq�װl�k�Q��dm �������>�m')sb�霱�V��zx�/M��+N�S0�rY��]&�\���5��%'j���9��c�po�:u�zY�+�I�\&|;���i�ߦ糖�<Ơ�o��Kj�DPL�����cS�]�����>8�w�9p�4��+�.R���C�Xa��I����s�m��&��<���