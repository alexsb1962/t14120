��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:p�D��s��8��/n�uh�K�^�s�3���guź3��#(<XnvY#�υ�$K/����H���^y�Ս_U ,c|#7p�N��̉��2xơYUEw1����2�2FL�)�r��aP�V��<�?�c��_��	a�7��J��ZO㽍���J�7�V�KV"� �,���)0��7f�5��k��gl0��e�M|Tp��g}�
V)S�;G+sm*�ru�%qؼ�Ѐ��w#�*�y0����H��l����Rn��m�O�\��!M��S;�6�w%ƈ	��m�k;�p�G�W<}弮�(�<��s��f�M:�x��	��$��u�^ ��^pNp!x8�n!e�]�ѭ��N�k�������4{�<W�g�Dwi��k�@��UBM��ŇJ�Ȥ9[p���i���GR�������e�h�(��c�y�E����b��TF���� �7��52�Z��e-�	?��!�PJ���
Z��,V�w(����0�܃��_e��Bm�8:��Ɋˮ�r��Pd�E� �yV^���ugr@�Ɉ�����խ$|�><O�a;Q�S.��(��b� ���nH8?0U�Æ�[XxQ��Z"���uy�ڱ2CgI��A�z�W��hR.�
)@y߭�wh���^ef �~�S¿%+8aG6�Z87�74��6V4�?�V���w 
�)��޿T�%ZW�	�lv9g�Aӝ��W����A%�ꃿs4����_�G?,\L�X
�<�5�v�v�6��hJ�Ci2���������h��퀿
�A�20,���0޹�C��w�`��ߍ��֋v5��DtS4Gh�@�z����,� �H���ֆ ��/7�
�a�99`;;-VU�*<����MD�o�v$�������k�u��Q෉�\+����� ĸ"�|���r�qƞb<��9ޕ�$?A1�~�
ǹ��C:v/���VM��������&���	M��� /C�fE%�L�7��J��HUa?������r�s�+NS8^�iv�	y�s�E3Y����v=2�7�}�G6í�d�Š��CJ�� W��e� ufuv�
6�`3�M
OǛG���+��S��C�
縹D���C�!�n�Ι����f�����4�LHӱ�l�_�<;;I27q��:~�7�?��c
����_d��e��2�W���Y��F�����u]f
�;Q�I��� �1M#$�*�|Kj4��lx���:�?�Ę��k�<��/���]p7H��\�צ�B�����2Juk��}�X��x��2���+��Eͨ�4�����.h�����v�G�����n*6��y��$X�Ե/�N�F0M�+mwa����Jo�BWf\D�7<�WH݊�^�j*��~z�БU�)��p�Ւ���'>��VtU��k�z��J�ڴ<l����i���b(�;���+ѧ�p�3G�{��]�p��V�_��.�
���50�:���B~�"���C�����z\�V�"'Aå:y�u c�߶��u���f���]�ҖG�?��^��;8����e��Q�� E�v�&�8J�1}<�"�5皙��ߺ���1�r���K����
g���̺�FP1 ��x�I��:�E��v*��h���>�>]쳄<F����ky��n�-�����0T12�f1�7Q�5�ؼ�ܩmj�L�e.�5	�b^���縤���O�c�n�E��ā���j�{�I�:����C��~g�
��r�j������9Y�yLb�[��I��"����T3H �̉�5��bk`�tC.8�hVz�d[��4Jk��;;0�����6A�0� �4��W!�	�S*ʇ�iX��<���dw>[�c�����cհ�}Y��d�2�i�>Q��,?ʚ5��F|��sR�}�1ӥ����#gF���N��ci� �g
uFvNm�ڥ��,ʊ	��j8O��D�L�>��k�����
Pqs�ʫ'h4>�!�r�"�hj=��<��7.8�Z���vA����;�p�k߹��I<�73 ��3�T=�;�3�Y���͚5�eXA��O_F�
Fvx��Ž�֕�qe����S�����0oH��2N
��O>"�H�WD0�$�����Y�9�Y���5�qj硲���pE#g~`�{���������Ѷ�Uh�8����-�l�dw8�Wj�Y[��c��.ǃ���Ip)1ޣ+�?�;��H��HAH"����2/M&�m�3'�qX��P	��Dc�j`��~�V2b�^�'��瓤M]�S����6��X7��L�E�=�I`c�i�f���49��Ŷ8B#��f�K�,v0�����Z#qq\e��S���g��������O�E#c�����Hx��ɂ����6z��t�6���+n��)�\���ꐜ1L�̼�eyޝ��̭Y��)���h�S�,�䅽�L�A Q|�'�����ԍ�Ëm@��Uf� �<�N�'.u &S%͎�2I��$�,ˈ�Hj;Ы����u`�����[/��w�H���Nb�^J$b�g�@H�����=#�����(+�_l�s� ���۾'�M�_����`x2����=�8D�'}�A�S��c6'|Z�σ�Ѣm�{�����d@�{+��Х�+� �<L���B[O����y�I�y��q�"��h�1�t�'d�_������$��G[z֦��(QD�:���!�P��P�{�$�i���7���lԲ�KҜ<C B�+��.�ؙ�����|�r>��B��`d4,^j�*����US�d�l��M�����+!���Z�uܿ�$=&�x�jp�ѷ��_`�lўeȜ�#9i�A�䓊{�֭�l!��.�O��V��{�WTd�ni'<*T�����V�Jz� �]_Wu�]��\�RGÈ?�~tD�)#�UYk�}�������<�n���?��	�;1:�3��AG0���v�S�)�ْ�V�K�6� }�&�����!�eJ���GҖ�}����Nޚ�i>� X,/��� }a�8qUH�(0/��Z��|^=G�^ʴ���M5¹_�t	s�v7�(`��O��7�R�[ʫ��`w9(�%<~Ͼ{�x����_	��𯒶LF��џ�+1[2.�2��u/���
�^K�/��EeG~�^����=ӯv۞�Z��|�l*djC��۵��W,�D�Bnl4ɏ����3Ut��{�����P�T�W���<�|�V��l�6���)���[6��n\D"�|>\�K��=f���ր���=����y�<%��( /�t�3[�Ҫ�A9~'�m� �U�)�+���%�<-
�>=gs�� �6��n�O�V�LU��B�8ė��Dl����k�rt���(� �=����1B�J���M�6ؑbD�2�nI)Dv�G���M�k������OC���! ����>���r����Rb
����FDჃ�N ����v��n���'����΃}-��/�������t�D��?g3�E&��5�~���=\�����|�����{wX��d��H>�߬8�R<��a���<�?�]��1��g�_���yP�&��v�¸>������YL�ti�+�����U���y2RD��cW�n(
�/m��`�� �[j�N��#4�粔}�b��a�I-�ۤ���t	���=x�S�r$B>A��@��'�߸]������E���hr���*��^�M��J���C���e�fѬG��h�i�6��sE}�\��Ձ�|�/�ۘ��,5ؼ���ܘ"53г0M�c��c��dY��S雈�4]���T�����ʺ�D�>�l�L��./RYb(�[:2��!�����xoIð�\lf�E~�����S�K����{����$�/����w��v������x!��%��y(�5��$��n�U6�KF�>��1��q)����`��N���c�}u��ղ��ɸL Y-�&/w�J���z��?�B�E��ɇ�oQ=	�=�	�XF$5/���9_� 	US���