��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^��������yDʨnF'{�l]�;�{#���?����,(G�Y"��.�I�=f_,�
� �|'Pw�q�HQ�	i��_���H���Y���a�s���O��yO=	b�FU+�Gy��G��G"p���^�L�ՔF����ƅ�A2l�]m�k6�p�sn$I{��nW㼻�Q>�̟�,KB� g����?�*�� �v����ٮ,�����5�zݧ�����=�>��j�|���N[�C��ｒ}��@��ӆ_4������P�����DC��+*�J�%���,_a��GO��R����R�
tf�4���g�����7.9�%� ���S�ͷ?n�n�?;`���U��S��26-�%4�[S<�h���U ��;i#����P��N�zh+�*/�bp����峨���_�4f�~�s�qE��o���L����[@ �2}���g�r� d�/3�L������:��w��a헫�G����дn���N�(,��S~M(����s�Q�m���5�^. ��>��}�Tr�)_Ŏ��yB�=��s]��>����u nE�'�7�'�ވ/W��mH�_����5�h�T��
>!���}&������A~�2���(O�6P�����jr��ޔ����v9��jz18�/�H1e�F܀��sY�R{�A��?��.��@�स6f��~Қ���:bc��r�ci���I�v�è���t�#���Bq�
K��VW�c�q	P���w�1I�k5z�N��W��FR�sC9pZ���A$O�,N"�.���?�N�]K٫�m�=��*@`cF㣄+=݇	�o�,*+�:�ZM\�$~�]�������Xq�d�O�x�����ۚ�m��R�,�?��T���؄���߲vyc�T�\漙y�Z]�)���Q�YGs6B߳$����Ku^��k�_��a8ƛ��T�n�S�/��ڒT�YBJM�'�zˮ���eժ�����<�SB3���K�m&�)U�^��m������9+����!�X�<M'Mnlg�M��[]<�I�c�_�ඍ3����8�+�sM"D��dt�$�_�����de�װ���N��mLKx�_���@�I1Z��ߍCÌ�lt��VGWt�� �,�e����$�`W�SBx�w��44�PK6�}�8�S�`�$�
E�ؘ�y�� '�14dİ���CB[���kHoj
��D�X<�>7Q8'�`��Uc9s��,�qcz�Y�OB�޲���B�~W�99b��|�W�/`"��,�JE5C��� ;��BR��# �r1UB��#�.���i;��kY]Ȑ�,���L�e����+!	�B���0}]F�w�D\u��?+�@Øb��v����!\�}h%�{a�;s^����<7��h���p�O�LEOb��ӝ$�_,���^5��Μ�-f��o�s�5����|���Z5m'��Xg�e��|_Z��RO��BX�l���	�1W_��
�!wE@�QRC�#󡥽�6Ğ�7^�5�bR���sW�|�Mž+*!p[�?� Y&�&$�� �:��I,,��C��y[����	1���v����P��������-с4(#X���?���2K��aX�WBW�=2�鿡(qdR<.U���a�!�a�����=N�I��w�����	�[��W3pƲ_H��}�F�y�o��ĵ;X�1����H���Jpu�����mD� ��k��-�����L�lQ��qN���H}����9PI'|�|W��p���e?'խ��9�,�S�HF�t��	~6(��%x���|��_�l/�eɖYw9�����~��*V�E;u\A�Z�	���T
q�z�&�Qg�69���9VKk�'8�if��-���(5��?��7�B	���V���� �?�L�GO��ޞ���;���P���,ׄ�|���)�J��~�!HS꠱)�Ud$9̾���ဳf��G�谄袺8o�<-�!�9�I{�S�j�����F��tC��T�������f��g�ɘB#�j���e&�Hw�Y>8�@�u��֍�DiE��
X�s� 1
����$;�b�0b q�?�׃�)�%�/�1�:Mj���/��*(��*�K۱���硬� D��"�A���ׇL��Q�[b{d�~e����B�'.λH ��<���:جy*�[�\j
�)G��ܮ����;��AQ�T�$�O"G��/����&Ш^(7L�{eu��mp�0�e>8�Td��r��4�kXL�s6%���%�~�����(}3��p����xoؾg�
z@�6�~v���k����)`�ʟBRI<�� گ�B�]0�a�RJŸ�ݯKy�y�7�Y�hb�j��<*L�7I�M�,��e	li���cm#�)�͝<��%@���ʱ�ο���w�I�4���Z��Sw��K�O�x֬��: ��,T��.���r>�׷?̹ͪ�
��7����`0�7�����A�p�-�m���Ӏ]�LW�U�n]cHɅ��"n[s\	�<��=o�R5�Փ`b�.����: �ԟ�uK<�(��ԥ(����j!K�.�O|*1H��!r�((��[����vI���j8��z�z��� z�Y���l���]?q����\(v1�8�<=�;Yq"AΆ����=�"�� J%Qr2yŗ�[3��JV������)y�b�2�w~�S:�_Ρ���R7�s�����;7��m G%ecT�m�w>�r��CW�a�(����R��j�l�!jߙH�$���� aoY�8[r�ѝ;O�����&�����\Uq�F����bW 	������5(D�����$��Cp3$��]�$��;��?G]��P+�C����Z$:�N�a�t�9
�-�gj���~���1��k��į
�����S����T��>q6�g�bE����x������o���.�{�kK�F��˟&��HD��-�M�nrt��m�Fv2Y�~���.�l�!�gb�T@B6ZR؏��K�`���g��L������
ҋ2�r>�t�(!�ez�i\�4A��fy�i�2�"�u�xŉ�� G�X�F����i�x"3!��D]�p�h�Q���17��W�T����+8�p����HQp�s��\��/�Y�y�q��������FW�K�v@�>Y���=�Uz�M��b	[��1ڙ�vxV�q��f�ȸ������ZՅv&[�����'�_�ǋ|<\�����_>5[���^ó�&�.�I���V	^g��l��J�2W�����=������2�s�������><uo����y�]�45���#�r��-�~�Ch+����?lOXf{���+3���N��S_�aV:5��sv���g�c�6
Vu���+��n)�DgԜF/�$O����ע����~�9O]ھ�d|��\ ~f�ӗ��E��o���ggԫ��LŮ,��<�;4qM�7m�����^5�r�����&�̚����8�ݛ�̞.E�c~���'¤���?�o�i� -T�;>@�nߦ�S�ټ�
oc��ٸ�ٷ��xx"=37��s��qsg}���	�%Y�o�ܗ]����hؼ���~��p�q�oɓ��pJ�V�3)D�+;6z*�ӚO>L�Y����{ޜ�bH	3X�cZm%�tE2��e�/��Q�f�Jp��ڑ9�.�J�Ѧ ��&^ƞ�ڨ �������U��06�ʄ`37�Z�t�N?b~���@��&���(w>��r^Tp�1e1�Ơ��o!��x@����.�����*��Y�8��U�t ƍy�3� �-�D����O���h�fO�1Kn��+���bVԋ���<�� ���\6 ���Z����}����%�o�e0���(�{A�)���ܜ��Y��3�N�"���*Y�L���l3Q!h�a"MA�؇��}U�k���]�GHHB?�����H��!�^iOE=���wP"}?,�j���f*w����心�A���3<�eK���˕E���a�6ߓ���
/y�-k�&fUSF�]^��!�3���|M��Q�-�me!ݴ"h�bD�x�?��h�LP\ƻ��U�)xQB,� zb�[6"]i��q*��	j���|B�����=Dh���Uw����RZ��6�̬�b1������+��Sk�3��d|�^y<�)�P$?�3�L�/7&
���i���ܹ�إ�Z��;+�AM�9�f�X�th\E$��^�C\f@�B.�B��ЉM��;̑n�UQ&�����^"����I]��vm��)��D%'���8_3�8�V��
�>->�@�Q(��+|������Lb�z�����\�)�����dn���ԗ�Z��SO�C%��u'�ST���q��!)%�A��x�2���'��v�	���	`��yT���2_\�0Gf�j�3���n��^>����ﾭT��|���$�FEN���3J0�
4y�&3d��
DZ}�f<�6!nc7 {N��[��i��d`��W̯�Q�L�b�I���9�B����������D� qP�0��ynys�y��F����Qʚ*�"�jH���pL�~�#����u&��yLBϬg����e�p��N�f�_����U{+d�_S@�$'����/6j;C@�9�E�1CBO���o(�֩{�r��h�����C�^�?V�#�%��k�X�@��<����ڣ[�1�hy,�5��1(����`C�)��;7T��@� +r̟�4���'m�x���%����&c�Fm�f� B���G��s"SѶ����O[<P9�����Z���15�.̲��C��=Λ�p;���Nh{J@��w�^�s�)IUQ�vs0�̸Q��ɢ>��,@�e?K�mp���/0ns�-ɽ�P��Pb9�!G&�u�$�C����8d������,]@j��ռUE[��B���H}wZ��N�w��0�%��L����=Кb��7 ����nɼ�9}���rg�,4!��X�y��)�{y�qz!5�\�_m�g�9�Z�ncY$	�Q�[���,�$�8 �B�ܖܜˠ��� �"����J�x <�&��~o*R���Q�9���Y��X�kְ^~��6��N��T�0� {;�7#X��obj�1�eG��Qನ7v��hQ	-�� Z:��y�:M[|�hp�n�	ۨ[����ܤ��Q�A����S�85Hr[�k��$oY�����4��|�\�}�OϕS�y}�9��v��Ń�S,	�I'��-��e�~}r�7����jU���3oP��3�.ef�8���M~�?�&u��]�/[`Ф<�	J�=̃X����m>n�A��E�I�����s12����B�7(���4�z�Nz���T�!q��=�K#8j��j�'�=2�gC��䦃{��^� 9�'+N��i�;&��r��!�P��(v��>.�����fP����*�I�k��:��缒��}�J��]���`���5���$#�:w^o��F&|�K1��,��o����@�"�oAE�[;��� w��`"!�S<l�%���K�f*��OuU�uz�)�;l4�Б����/��7�4�����=ߙT��`�n����}����	�!'�M��_&Kp���W���/y9�d�vr���[
3�c-F�Kgȃz����-ݮ��80�v�[T�����U£�H4�4�Iy*�^�ΐ>n*��`=d@@:�Fb��o��'�O�z�CKEx��t�Hݛ��wf3ݝv\`��(�����Ga!9�ص����Y��L��%٭@W�W�B�����>-ՐX�������Py��t�[�,D}��3���G擗1�dѠ�P���k��@KWRg�zK ��/
�7�E��ڱSt}�Dr�奼�*N�{�3	8O���N��݃2�_˅H]��P�E�.$S��';�H�޼7؛��K��	"ߺ� ��������sW��J��o�m��@-H����)�����d��@��{�8��j�=����ѣ��?���]L_�:`VzEezB���E����Y�J�G��rBoH>�H��Bn�9�T���]�ꆔ	f���:Big��no�z�1�^��׳�"���P�5Ǘn��Мr}1����>�<xe��a��Q�S^6�Y�����MO{r�RHd{���C����I��ڕ}��0-ف U�ܶ�ƞ�2������R����21<\��_η0��EJ7�U44�����<%�N��T,#��q��}���)��4K肋^!��i@��>��C�~��j&�4� s��_�j`���}<ZՍhfr�XXm�s��]���d��(=�^k!�5u�%Ց��^����kt�1v
���J]t?�d2}����2�F��P��U�R[�A�I��j��l�.ad.��Ps��'�oQfH<	e���L���Za�x�ƿ�K��a��EL]$v� ��H�w�td�R�${{�8�2����NшA�Ԯ�g<x
1���|;>�'vhG���8��~M���P&A�rs{]i�~�����xXrq���ɂ�"��O7�kb9imN�"E6S������VCb '��e�-��nfV	%	8WX�+�����-jFa�P��{jz3;TYK��9����ۏ��l������y����ܒ	���!M��M���)JfֲIU��.=9>�e��}�o�Z�dp2\�X�q�[ͽ�����9��� ����tʏQʙ+��,�	?2����|s8��Y�S�YWF`�gqԀ�����0�V�)oZ�G���z%�,��N"Oeb����3�]l�igD���6���+�Ӫ_d��Iq?�h���m3�I[z�n�Vr�W=x�jn��`�+A�)����&k��&j�⑋*���z+�=`�Qa(DH��F&L����JP8fc<o��\�fO��fi4a�����cfݲ�rz���R�s�����ɷ��%��si��tJ��ރG�'m����Y��ϱ����s�������D��ԶX����zJ*%�:��e8�����n��sI ,�-rd��ӐJv��O�y�uE�_��6<v{q��m�߮����5o��X �Gw�����9Ò�hRv	���-hj8sDd�o�2~�-G�i:>������t�=��= :�xv���i�D�>>��/��2�����v�����\�o���X�`azP�;��5�=��X\�4@�UEH��H��
}�Rr��l.�r���C�D�!�#�iY���"��QJ���ca�����w�K�#�#�9�٪�������� a�{|�t��G�ٹ�H�s��X�ʉ�F@+a�E�B���=0v�Q�Ќ���0���v��$}mW+l�o���ktŒj
	�	@��?��|>��20Ҁ���RP�z0=���7�n��\�[Ϥ��Е�'g�#�BE�k�R�����L�r3��W�4'�y`��#��R��܆�eJ���΋s�#Ц�Z`�du:/�0{��= ;9>�/d�fB����ɣ#IE��5����k$R�t�O�A���5���m!�c�	�;�ͦ�N�#"�1f�E�4"�a5S�(�g*Q����?�[P䚘�(���K�%��)��]r�[��6�jϓ�г�:�߁GȄ�D�8��]�d�F�S��=>.��SM��hú�?�b'�B��C�V�������Z"��;����x�Q���-�]�΀n�:�����G����[�6\C�JL/)���F�/"!x���%����8缚��zh���
e��	�8�d�q�4�~�?�7y?M�w���rqY�<��%��~d��~|�B� 965e"CPJŖ'aJ���t���#�{�qI6p�zE?�`r!|a0#Ίaޞ8^u%�پcM�+x���{�%����$Ln��lW&�*����Dk,x:,y�-�xD�]	;}����꧀�����f����̥u�'ԋ̠��.h�=���+w�z�'}���8�"1_,�]�t������Q�]�n@�&�툿�,FS�0��=L����K�Qz �Y�9��۩�I�	7<��px��r��ˀ�4">���j����~YDr�Ig~���B����Є����|��t�΁��4��x~v���Rf)�Ga��c	�t��e��3m�U�1�B�R��ÏQA��l�(�����X.����Һ�dP��긂��[* ;�D��^lSud`h�n�^7�`�Z+7�*� .M���;e��nLdO�=f6�lH��*��ȼ��Y�X�I�hU�{g��+��T�������8fZ�¤� ��;DI���7A�"�N�x�p��W;� �w�g0����˕�rC!g�:��x9u�Nl���X6�i��Ō��,�SQ�C�zH��/������
���p��������;K~��	r�((�h.����O�9�a}����e6g���:8���+
�B*$K�`M�i�~���4x���v.-��s��eu��S����� ����z���w��Q�,�{�(޶�Q�������`8�s�[v�Ez�M&�^pX��,����9���٠9!��tM���C7�nd�ٴ0򿃈~usƣ�L`���зE�K"�:}�@�����!?p���d�b'�����U���Q��.�^2I����\f�K<��e$�%>�[xͷ4Ɂ�"�`�y�S�{�>� V��f^\�NR.|!�t���fu�d��A��y����$��*k�L|ۧZ?,���g����KP<顳�f�6����p*%"X�V}[���s�i��'~�A�%