��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>�� �F9!�/_g�T@_hm/a3^��(#z�dZ�E�����v�h��|���-�>bkgá�G�j���zA�;h��Ċ�k��ׇ/�gN�3ӟ����i�� ����4��m�"��]��V��W!��J乧1�u�M>w��;��
�̗�E����@<S�ǿ�α�7C��8��B�TGEM=[���b�#@sr��C+�:�]d�}��.��{_e[��9#2�_�IQ/���*���ڥ���Z(4:�	��k~a|jg��ӹ��dY+@y��k1%v�J��AW�m&kT��v��	���lT�I#-�T��-�L��kRv��ڄ������s��.����``uc��
���ˢc�����Xr�+��ů(~���,�k��8���3o���'�����tM���B��~�V�m^����n������Ȳ���b�-�~B��=4���
��.T!E�|��+7Ik�P���.�uA�Wķ����Jgd�,%��u R�*y��Ŧ_���,��I~��Q�I�$�F�����S�&Q����ǝ;�AS�V���h��.�M�����Ԁ��x"��Q=J�?8��/�Q4S�������R�P�#���C!!8(�0g��C0�\<:yg�I*�{��Ur�p$ʧ��B���\um,�`�,�n�w�wCG���ec
�O�����Aa���6T���`�c~��#���h��׸R����k:m��ϞLy;Y6�*V�ڹ��^ǣ`3����G����ߓ��N)G��pAm�ߐ�=����e�փ	����(��)	�a$@�3Oj���UqOe���[zC�V�i��5������޺���@��D�s����A����ZO����7�!q��h��>Vߞ��?�@��(���:͔��܌�oJ[��_�B[�$�M�"�|��!x�0�te�F#j��2�]!�	�gS�wE���iKP��E�[(�M����kd��_k�w~0��h�>!���I)\��4��[��9��W����bj�����v��h��T��ݣ�u�!��]�x<X���F��6��~k��1~�18Ӽ8zyX0rS�d��ƌ��EGƞ�q ����j/cڞ���6�����˯DsP��4zf�^���r�>?�X3
���Ίw;��&��vi.Ȝ�ֳ:o�-I+7+�)��U���},�v^�kp��G,m�K��l]��ֳ>�\k�_�/��J��$��0�!A���颇�B}6&|�_q��gqD:�hmP�g�Ĝ�A�-�Iۅ2�_���_�i��E$����C�G������p��6{��{����� ���9�<�e؊$�,���2u��d��f+@���о&���fTKȖ[H��119���]�o�|���D;�c�˶���N�?2�7@�Ϥs&�<�I`�'�#�ͅi�)"� *Z�l��q����)}GrI�q�.c:[�ު�YTD̖(C�G��{�'�;<O�_q̷ϼ(�_�%T�k7h	����0{)����N���7$�E钌FZ�g���k�ԅNzJ��ɘӃ	I#���R*|1.{�?<k�,ﲺ�E�Y�7`���}AE����WR7�o�sX��4��&A�-�G�P���V�����:K�?h�nGwMU�Մ.@l�+ʵ6'�����\:f����m�?1w�8�l5��S.cL�}Q�%}e��d�!�S�OwJ��;wp��d(�@j�_#�术�Eǿ��RT�Y@C�d��܆��M�(r���f{t����0�`���A��C1�Yݔ�ꆵ�^W�q��ۇp�$+Ж5�{�L�6�	����(��L���p�}7Pj���o%��,�V�w�D���u�2zt��ނL��L�"�m-D�;i�G�[�\�~�CV}էC�9��H��[|(�G�m�9���څ�%��G!m���$��m-��׋�A����'C{���+�[���I��q�7׸V��S����f����F�����8
a�1�V��n��:���A��fo�㷱	��ҬC"{�	��W�\6���ԃ�XkH#�KB���$r���V�Ikg�	��c�$���ذ��Z�3Ĭ'������LJ�1[�LJS�Nq)��씣 ���1E`��,�Q�l��z�N���2��S'i?Ds�O�t*��ܮ�<:�h��s(u"�2��i��U0:���9He�4�h�D�S��F����-�g);d �ܼ�[EL1�!�\2!�� ZϷ毇�=O9��>�Y����.\voZs���W��'^<�:�C�PQI�E1�������@��R�\������e�P���k��_�>9A��t׼<�6��?:3���?�HW�g%���oIU���vR��G��}(Db:�I�wB�%�?��$�v����$4Ż��	w��_�aǐ�C�]���b�k�]�b4dZR�3�"J�=Ҁ�״����e,�-�䫓�T��:�$./�kD�AU�%�bQ�v@�ջ�	(rw�<\�)P��r"� ��B]RJ�K#ؖW����e���݊y�8ބ�:��%���Hh��u�o.���Ev�KOw��Ƃ��$(d��0���K�x�xqv.��	i��:�"��~w����T����U�����k����ί =�d��q�+���H#�b�� ����\6�����+��� �Ͷ��&�B�⠶���0��Ѻ^���6���bN^��<IV������ �\���|Q����⛞��?��2E��Ys	�xCF�c���E�z��g��N�zwNM�n����}Tw_j�bH�S��{у)� ����D�=.x�ɥ	?C���	�c,줺�3�n�z���APa�Zn��e/�R.�IX�b m��L�O���^�%8�kArζ��F�;^���J8�#�v���Z/\#oM��k34ؖ(�CJ��=s<X����(��m���+�:�ñ�)V5�������gO>�2n�DXk��z�ʠ�U��/m��F�:���C-�)ܙ�E����V>/[�����'"j�ӝ�`�K��[�p���5�u�������g��Q�5Mb��K�Xhn�F�9|�Y��i�rk{2B�p���tÁ�h�y�����1�uX�<�R�w�;���h�H"4h�v����*5���ģ7����El���g�B��l�!����%��,f��{���\G�'�RxS��?{��4Es�a�������� !�H���y3[�c���2P\b�����J�وG�!<{d��$u }k��Gb��C �d�?"�V�d�b�U׋'Um/�o����8�N)�v<�ڤ(�Ż���\���z*(�GĂ��yz�+1cK(3Y[;� ���x#�_͕�o!�������
�y��
�eB��궃J�k4�B�?�iYa"�.�3%�&%��ѣ��z��	�	vp�G|��9b����=�e�o�m?�v# ��[�"��YL��yr��Z���ξ�����Zx�8�u6Bv~�Ka�9wh�Ff�㙺�$%�ME���"w���yV�Ta�� �WHJ��B�s8|�E1��<mHB=��tEE�hK��IR/
��yz>����<��:��k�&0=��dy���!^>�\��0{�yϫ�ů�j��#��u���*Z�oa9�È��T�T�K�}^i�'#����F�&>L�/��"hU-�Q��|髈p�H��)؁��gP�銢S��qI_˧(7����