��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������L�|l�c�M*3����1��!�\��kj������C3:��ϯ�e�aͺd�����pO,���J�0z��h�x�Р�X�����OK���p��F.1�X�˔�a�7�Z�M����q�����/�^nu��Ay/֖�K����r�KE�n�Kl��o�6�Zͅ-=X���סu�k��;ע�}%�Q�r$o����^G#�lT�;�H�QS��Xb������Uއq��{f�N�����i�ֶ�s�nJ�f��C݁��\�0p�Ebx<���oF#���B���)�}��p�ľ�1!h�oT����D��쳇z'zl2����D�4��F�\�n��va�Z��D������Yz�xv�$�{Ex�C��-�1O�χ�y3Ex��(u�S����K��,ҽ�H%)�`�r\��z����3o�hM{
���TV#f�;ZCb��p��<#��^%?�J���_>��G�1��'�^*!��q���H��_�zQ{�4t6p%�cf5҃�y/H����.8��C=�`ō��+�tŖ�a�g���}_��d���!�׽��w\|�<��~na�Z���H��_�^��֚�C���Tr������D�X`��T�X+J�<c���3�`�B�X5#(�0��/��ٸ*� L�]jDU:�o�HM~�A~"�-��W�s�J�l�&�������WǜTc�OU�e��	K����v�����?�y&q�P�e��Ĝΰ"�&s���$ջn;+oL7�tĮ؆���!-���V����H=
�~(��V�L�s�|�+��k#ɇo�y�b��f��K3�F&��/j]׆"��~��BT��2�@2#�����c�Q��?Z��p�M���q&\s��&a�v�����1W?/u�e>z˿�y,o�#��֨��;y���biĀ��:���{y)��-�E�������ґ�l����4+�+�gUS����r�\� ��#�W��9G|-L��=��+N  ��z"L�������{�|�q�w�q`1G<1cFx���hm�L�m���Лx���rMT�=��G������1���S'�+OΌ���P���:I=a��&R(��+�j�E�6\�#�`���a��Y?Q���;���������+�M)�X�� ��ի��0��\�r��d�V�'���_�oƣH5�Oa�|Ϛ�&��'����P-�y�C[2եj��h0�JU]\�<� ���a�!O����%����7�G��j*K"kM�3r�����{�92iEh�_-�P,�P�w��w�Y�}&�¢I��I���+�J���֐ 5�������}�eخU�.c�&�b: �m�)_��!�ą;���<�ˎW�J�P���g=}��rtBBE1��Z#�����I��گ�n� 0���~�K̖�eE�����<�_c�]�������l���>��2�!�B�_t��ԭ&���R�sU���k��󿅜.n�ObtN��9u��ӕ����Q��K����!�/�M�{����N�b&cEK��N���lX1� ���c&�q����[n�/'l� ���?�Q,GRU}G�L����IÑI��Tƕ �%�`��
���r�(��8=mߖו�]S���D��+����J�@}��0+q>&b�p�x�C1�
|~�T�Fƴ$w�S8o��S&���r?�	ظ�h��p`�[��Oeo���t���O��c�b:Ǻ�z��Cu�Ig�W�T ���v`��e6Ś�G���,���#�o��ȹ����Ѐ�	��D۬5�ɺ�Ǎ����-�\���l�(4��e��6}3g4 ��}uڮ2	ѿs~VM�@�����w�Y<�X�сGn�jO���{��ؗ�u���'!4�SZ����Q�W2�K���P�aX�j@� ��w������v��E�9�̈́�����'��&WՇY� y�((��#X���X�#�N��8����[��K�_ �eܲ��.�D�(Pa��i`8�=(bq�v�.�S�9� �g�C4�fR�G�>q��Ϧ6��I�RjiU�Qޓ���0����S��?���<?�Q����Kԥpn�:��Ss��4R�(4xl��^���s���k=z{wN�*@�8[Bv�g'4tF�7�/m]��~�dQ�2i�����#��O����d��r�:�IG5~�����&_X2U�ʉ���"�C�������C�8#<���P�v�e�� ����~Ԯ�h���9��R%88�{6|d5��N<���W�Cǫ�Ff{|w�o�]��k���׃ԙ=^X��k����톀BUr^ʱC��HuB[��
�7�5iUY��)|�ݼ�F^�]d"���� S��D^��BKԖm�Qj[�,@L�r���1]y,��q��^g0#>,at����kºuRTL�A#�j�d��IC����/Hs���NH���F,�V�>Rɽ��ܽ�(>���g���%��� ,-�q'�m1t�nKr�S|�.���CN���^�O�G`�3�#��]<9�� P��:��5���|M�/+�汷"E;�>�_l��dcZ3�����An���з�
���ز��zS�7ӡń�x�|�)���=�Е��=�^���O��Б��g�����T��^R�
���8cn5��B�b�t�%�@�\N�`꽙P�R�҉<yAc�Ϭ�O��+_��}	R��_�=���M@�R��X�s���m�yi���+�C����I�%|D[N��Д��^�����A�H�/�jג;��� �_���8����K���U�+�4��KbR��q�{�tŭ���0n�g�1o������闑쀓w�!�	�7<;�U	^��j#z��~rʲ�����q,ޥ(!f5*^JT	ͼV��~'��F��_,�_���˸��:{�X��,?C��c 8�)N�RV����`領�eգ��]Goې]rSHj�g.�b��k�ITkU��ާ�،��"(O�zOx��M ����u���^4ٺ�<�&4���M�ݨ�[5�&*D���:��4Y� �� uڄ7� ����ê
���Ŷ�A���AHHE��rJ��x �!�����6�>�Pl���[ƲPM {}�❃��>UTp̉����@Pq�g��h/�+���_�>m;B�������0eK1kQ!�J�mf@3�����*{4��%3��A92�Q�.j�^{@�ʨG�� ^W/�=�Y>��bm+F8+4�0�I4��0��ʘ˃b]>��c<:��,!�1�~e`�YɁ�5�@3��������y��ئ���qf�>��N�*yqP?ul�����M�&�=���|从-hFHH0��d �t#�E{�Z]8���(�t�I�BXS���Y�� X�i(U��a���|5�|X�J۟Z����"5�VN�����B��K����M�.3)�����q��\��0�_��wx���w$6�"�펁�l��~��w$��3�ƟM˰��O��L��8�,�ZoP�n��y`yC�bSO�Q�"��=Wۅ��g,!*?̄�Y��U�sA-p��5���D��|C�R����vZ�4�������9F��$(�H�+�"�/4�n].��g��.*�j����s��<J��Yj�"!����u�4?��,�Y���K�^ڟ�b�o"��s�C��3��+_D���s�%��<�w�2P�`�3b��Υ��h���w>��.n�����砃v�hPr�8(=W2�zd�&Nʽ0�{����{i���ސY�<��`	�߹B[П̯�x �=���\mn.�v��ch�oW{?�N�	�$�~ �\<�Ol�>(6ճ��܃�f�nB������f:�'=i��z������Dj�TJ�M64��O9���E�����P*a��v�Hv�<�=�M��"_��=�Y�p�;u�Ϯ��`9���^Ӵ5�#Y,Kz�#�3�Y6��>;�"V0}#Hd��|*����R�d���F�d� ���d�fڂ��{8��x��� �8�Y%��4�y�v%ۯ׼3�T�	��J�x	Ζc��-�x"�A`�/|Q�44H��Vs�P��n�ŏܐαM�*�E[���ӡ�����f�������&*}�Q�i��lmL+��U�#��a�2���f������<F�B��1�Z��Sf�LnG(V�;mȐp��~8�$2��G�_�>L5m�9w�]M{�E��EL[m;bG��氧Z_�#�ƫ�*�fw9��U�ؤ^/�g<��$����W�b�M����2����&�jL��w��w�p�Y��j���N�.�_@^��F����\
���<+T��!bm��j���q���I�k�v����E��`�/i�̹�ƹ�����!�+PZ%�Aa��x���^�����eE�7�X��w`�x�S�\���
�iJEZˠ
]t����h���̾N���yo����9w��<H���v��#�.JQ�\n5\Bb���ie���F��K��E�#��*w���iS�ݛ�}��2���R� �]7�ڮ{E(�v$���r
�I�/��g|\��˿�x�_��LTg�B����&���?���;�y���V��5�I
`I�A��!aE�iU��6[B��0Y���6�F��0:gzS*~Q�
��ag�Q�X����a��9�%�~%(B���-uw�;x�TD`�BH�MA6y�ҷNE�Q�pUhф���3�ElIȄ@9��h{��ǉ�p�E�TɲA��Y�Ȧ+8������ˮ��!����N���TN"�����c�_�ص�TMF��3L�ة�)�ؤ�Ћ)��)E)6�(��OLYς~�)����t��za��A��r9��v���� 7 b]g���-.`}
GD:�h%���~E��bGnF�1���P�׽KmI���|�i��'ė�
>2؎gKO��ߛ��DN#/	�l�Q�<ﶽ�͛��q����Y���FVfeNT�������#R�^�wu_��m��Jx;q��6��PX�N+�ɺ�PT4q�1k�����Rn.l��?��0������Gǆ��V��_�@