��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����Xͺn�Q�ʐ�Я=��(J�9h��]��8��@��Fэ�I��t�,�'쬱9j��t�yC�.ԍ;�^�m-�]��R��"m����	���ZF�cX��V��t���P5���W�W�k�$H�\���1�M�h5F������%^��n?NO���t}��`3]y�:��O�s_�ڧ�8�:�M��H�ߛ��;�7���D�5��u����'�����oAH����a�8��!�\BP��aV#��G�J��u��2�*�p�G�>�@Zm�f�jqj�N-���9��*��qb�=�ۜZ���RN�T��R>�czuyvg�V3�%�I)T杄P-�Z�1h�SRz֘��u��"�UU\�&��-����&Y+�fTgV�?EϬ�@��������O�aH��1�A�V��+��#��D�nO"�ʬ����^���0��q����z���	�r�n���[�H�́,�y`dD`�O]s��F�x�q���\�ঢ=j9��8�ɡ���8Թ�F>$��X�a����o�9��2�YY��E�@���ɑ��Ij:cw�]�I����d�m7
[qW,H��04���
��@�
>i��B��`��{5o�6�<�d^׳��n�G��������1�հt�� ����zI'-3����/��*.�Č�q�*���������I�BAf�G28b.LJt%��/N�{
�g�Ahx;���p��g�=�v��� Ϸ:Ϥ�����i��!�;gu}�^�I�G��.�Ƶ��	d�����0�����|���c�ׄ`��DA�\�06m|�0�,�kĠ~�lC����f���rj�[��M�p�= ��0���l5U��z�3��I�IS1�£���P	\���A�P��ůtC.A���(��}z�o�h	����]�I��h޴�A$f�B^w*�-��
��:��� �o6�'��U�+Q쮒�}z�tNL�2�oJ�b�7�v�t��m�gø�C_E�}�9z�=_		�?��
*���P��L����r�}��Cg�v<K��&˗�B�^����&��0N��~�u]�t��I���X~Z�'��bN�N����Ӿ�*������~�`���QT?�qiLh�����7kU�O~,�_���n'����=����2�_��^��JPl��y=�ϵ!��\O{���%}��h�U�7�ч��k��
U��;O�u�B�r@s�Wj���_T 4*����ʶ@�Զ}Tњ�|C�F��ΩhUd$���3�}`q[�}�k�wn�s��<	��
!�c�
~A^E b��B ��f\X?���]A��U�����y,�d�&����ɓ}���d���*���Tr3E*X�|�گL1:�h�o��AM�r9s��I"^Opѓ#��VB�������)hҰ��k;b����V���(?O-l_����km�/3`�=-gƳ�M� �Հ4S/�*)�)1�-�X/ޝ$Y����>(� �v��eW�'�k��> ��; i��Oւb�/�>�Rl,$k9�O�fX���;I�H+m��Y<��Y��k����~_-\6E�uȖ��p���Q�a�St��v������n���-��g�J ֱ�CQaD�����?�x�V;�-`HF���Z������R����P�(��^^�U�j,�bn�����A������5<	��K+,���O��j�.Ԭ���21��7"3ѓ;x�|Q9�n�x�����{�9j|:���M�#���'Q���h-��$Nt�θ+d:�1�dHl{��P#��=�ۮ��@������|�]�a뎗��ϯ���BTTQ���	�u��J�4]�������3��Ug���`��w
�X7Fp����X+�4�a)�ޢ,�U�'i��w��:0�u��o0l�Y��9�:֋��<��j�F��$2S �6(Ie��c�j���/��8/���1�W����E�B;�ŹP�G����Ԥ��V̿ %U�����DZ/K�>�Qz�g l�p�/��\��ѵ���BcuTs�$�,�S��������"���O(�a��K�=��K�-d��'�֟�"�=��~v(�z�p� �f>?1|�wM�iPZ1^JO���qU��귕v�ر�b��H�q�2k?8'�.�=P��VE�p~�dB8վ\G��x��l��hS���h��[� g���>��v��&D3cg�K�j+��Qۂ|>�TPJ����W�n�)|l<;S���ˊ�Z��Ȟ��	����'��G��PRa�$L�s���W����^��!����fק����r�6���U$���&.�c��¥�����o�W�z]�$�>��3Q�򐲹�}a�`�m�N
g���p���=�P�HY��anCq�����1���	�.��='����|oi�:�kZ<���P���8��Gl0���U�'z�u�?lb��5z4�O/�v:	��i�.Aj#E,&�lR��-�&��2��m�pն��O�B������5=?d���&���j�����}�Z.�:?:8��+���c>d�T����!��� ���8̵}p�g4`6�O��F���_��MnG���Y鮭"�x劫��y��; �N�k�6=�1�<Og�x�b%�ɱ�O��μ-u`߉=�9)@��vKkG.��H:��ݷ��K)���p�P_=���by�0�Z6L���� ����"b�/h��1#�X�M?S=��3�4���Z���J��l����g+4��]�@C����h|�p#A��R�Ϯ+3�d?��I�/WR]ia@~⏪��!���{��̇�`�`x��� >�Q�c���iM,��4^�	��� ��U�4�.M_눧Fd<Lůd�ډi�r�l�-l���㷱bvZ���kA���+g�}OpJ��=������A�I�U� ����g�D����<2��_�5����N�I�[G9NRuh�~�aSG�n"�]���cĹJZÓ���ou��&��|Fi�c�Q�~�@9�KH�xT:,J(F��a�F��bP�z��H4OMұ�Xq���k>�C5V��dd�Z�B�L�~UA���,��`�%�5�0o�&���^�a�fQ�sgd�5���\�53Y
��	y=	��=��<�So	�ư���$��_��TF�2P�G����k>&���M�K�� �ꍼ3QF.�ΤRQ�Ƹ"UCYG̹�1ÅM����^�?o�T���ly�X�\����p�O�.��B
LEN���c�+Y4��]�Y�}�oU4��$D>��̈���(밟�؍|����#�<����{����I!�}[$!�Wz��E
!�(۠*��c�:��Aa�y�EK�V�x�Q�l�(|��=��������]d�HxB5�d��-#������"�
��:f��<wd0O�o.|�vXM���Ҟ��`c��<���c&.j&n��Y�YL���	��N�FP����`u�Nh���10����?�Th��I1'5��!G�O*?�a��H��>�ߓ���"���/��˖R��V֐���3y(k)zbw֗� �u;~�5�.U��I�a�`��~�=B��&-�kmo�.�� �:����: &w+��_��s�˘����s��;Q��P�`������ ��b3��o.�+Qf��&�`O���d���*^�+g�ǌ���0�?�J��tX�N�Lg�K�~ �K`��c�Tћ/|�+�ƿ��^;��c�b-U�Ɣ���<
s�:̆\z��)5[PvW[��[��ʂ�c]y|Y�t��:x��%�s�2�hC��q����c^~����d#GhV��/�ϸ6C�u-g�WZ��������O�=�c �+b���]��(Z5L
X�E��k���7��%�>T����Q�? =V�3�Dq$�W�,-}�SƎ�ְ�&���l��R�m~ڼ�;{1���5��(�V|��;�R��A�ߨc� $�C�<��ӽo��BQ���C�o���Ɓ�#q �VJ���Z�4!6#f���b,�v��b���K}�� P�fb[i�(�Y�ă�Y�hE}{�_��i4E+*��]���H�����CY#��f��.�� �9huq�d?��'z�x[F�$�n�����/�4�@�Q�vr `0���8��l��W���׮ �Z�����ו�#Vj�ٸ��OX%���h
���nt����|G���%\Ń:<^"��yX��p ��M�?�N��V.�ў,j�ӕݏ�$8zo�	?�6��)�� [�+����o1(�>��B�����s��8{n7*
v}���EL��+���H"y� GToG�+�q��ؘU�����������W C������h��Q�N	D�N�NぱQ\}~��?���I��b�\�!ƽ��眙ׇSzO`ק�穰����>�gUk�&�ŕ]����Y���"����>���\���(�Д�E���r����|�Ǘ`��u��僴[|Q��51jGw�Q�3uly���kFEA��/XJ̖�q����B�H腻8rt:�(���xa
�G��?X�
f��^�kۍ�����tܦz#��!���]~y��y���B��4�R���ݡdX��e�~>��z0�t����C1H�QL��b�Å_x���;[���K1�r���z�2w�tPރ��8��$s�=dkן�,�l���e��%�+�u�ʃ��Ń���O���?��8�a¸EW��(�/���]�2c�G�4���\���t�~ܳ��wga��]�~)Ԣ5�z�V�?x��1���^�޶�t{�HU`�f����-{͉dm�!/�,K�y�!ٜ$-j[9'��B!.sC2g�'�����~��HM���_�ݸ���c.:)�
i5{�wQW���$,t)r�X��������H�xQ�	� u�	m��k���{�<���k�P^�f��}�D�_H��g"��;�sY�Ǆ���y̓��!1W� �]wq����M���+<�� ;pJ�RL���bf�c�03�H@"�����S�m�w�I�>4���I<��'�2̿��
��/�;�m�M�-��V9nzu��o�E2M6�Z�_�뺮����P&�4���!��e��I���s���QU��X���/�{S�	A�ռ��ԩ�D� �`S��&R3?��|u@��+�5xid�9�˰~4��dc��N�ܖL����T	�D(#�?�hb��X86�򬮫�d쪡����6F%^ףF�o��/+(wJ���(�6D��w��i�\���\�%hۋ�G�c�=�y��i�L�ǟ_���*r���z�q��p)��]db&Ţq���T�n޼�`y�Y�_H��>�pE��%����`�D��h����!��>��oU܇�kK#�Q?w��l�++��{T���0�S���}��nV�o����������䠴lXD�#��� 0	�{�J�Ru��F��ܺ�HU��ˊxC��G#��'�6�WH�����.�P�X����u#@4iBzYS��S g�¤�{�j�Q�ZogL�%4-��
UU�g�cWE\�#0T@R�N�T����˧�2�+�y�R(�UAJ���"� ␡�d�b{��vz�t�W�3������R�sc&��N��͘�.EX
">�+*��91s�*ؖ�����:G��m��W^=���~��4��V�ޗl�y�=��$yi�`W޿ ��ө��m��Ln�ڣn^nk�v*v�I�p�YˑQ�y c-`_%�����1���6�[}3�{�7��P��F&,���9��?��~��;j�����g�"��㽼ڏs )������=�*p��E/n���M�8��gv���`PR�FHI���G��-m��- �$�a;�'�(�j��z: ��m���K;�����I:GG���?Y��-<��m�~�zܘ U/f�5�)*CkUc~<o�/���T�~'��-,�I����[^�_lh\�2�P������	"��Gf�6d�{X��V
���P��'\��������
���'Іɖ�6�C�����gx�c1��'�6�o�"�0\v��:O�)�����̒�s����q�)/Y&�����H ���n���t����|N�^�����|���3���	��wšʚģkxƩ��iM�CK�0�Y&�ۘ����~��1���H~o�-ྼme�R\�Ol"�_8��den�bp�3������-��e��$s��U�q}�����f9|R�"	>�hK�kI�腳*X�N�<�;ֽ�<=�����X���k��I�<� ��G�ȹ��s���x�N��LO��A;�7Z��i=g�]i��o�㣷�Q������ȫyT6���p���{g�{@�`p��(re�~�$"���Cס�_�lV�\���\t'��� !JokF�et���gyt�t����v��+%+����RHj�A�kd˚&3��P-g6�W�5c��~)D����m�V6�FS��FMDۺ͓��=`� �>��ʼ^�_�Ui����%@fy~?Я��!gx��2��T*��o����G. �}^D��-f�A��׆���1���~��я�tm��r�ޡLE�b��%FnO�١�'x��NB! �Ę,-�%G�ߦ_��;rY?z�%�`Ǌm�JG�[���L�����yE�|(H�nQ��l�$C�h�lX~���V�݂�_ �l�]��D���/��Y�"�>��y�aI�� Z�f�z��»1J��h4bfp�� b������f)��)3M�2����g��.i�k�	�+s_�5^!ই! �8�HdA��=��V	�i�A_`~��N�D׬�?\S�������ɑ��Y@1��
�9H�ӳr{"�XB�\谻�Ѽ�T�>%ae᧐�z� >O��|/$�i���
�u��W2(�ث�x��Mj���5�H+���n�%�����={��(4T�J�hw*�j���S�O�C�F$��]�+t��\ �wa2��K����~&-��%��_������ΚW�M�B�ee�EbH���ԁ���{� 𻆫t�E,kɠ��|ĵ���E>�U�q[p֗��� )٠�
�V��?��=s��t���u�d!��B�anh�X�Rw�P,R�qk�(����M#����W�c�0�'�-$�@q�8����&�IC��.��#��>ZT���ʮ�K`U��V/�H��n9 D�y��E��зVA�v�rq�*���a$|��/�CQ�K�="���c6�ʚȄ��o��Yq
Dҋ`��#묎�!Q����sd6�ƹŇƕ��"IN3kdB�3S<�ڽ~��'h6h�UKqh�׆�}7��-�Nq��nL�qk���+`
�j�����^�)����� �:�F��K�!2���d�|��i�͢�?�T=�A��FT].!�f�_+/`��y;-
Zo&���lp|y��)�mH�5�mHe^
:�������Ձbc$03ߪs��J�	f�y� \r�4�10��iVL@��w��aq�)�)��m>D�����[��e����-��J^p�����U�H�K���V�:+�S�x���5!���Rf�IeEF��<^?�<�������騀5K Cm�k��<��b�W8	��ϴ�uE���Ö�E �����W/�~��a��uDb�W��b���U�RC-n�O3s=�ۏ�
6S' GB�\���wdbk8�Ch��o��� O����W��
�t	��^o�Μ�tv�/c�PD +�%D�Ղݴ�T�:<2��a��]�p�-����I�Â�r���6��-�O`���D�۩��Df�S��^��+g��#B�7R�� !R>�������~i�>�xȃ��gz��h-<�7��:�X[v��0>��Y�<���Y�OV�,�#��x�:u��w���graU��)��!�^X�0�Ī�U���5*w���@��E�Y&x��Xs�*Ks�D�8��8Si��B_�8�����r�vd���Pa��H�o(�N��y�Θg��Fkd�w��>e᭡5����R��>Ce9� ��RȮ"GR�T7������7{Y)�:�i��`��ꍘ�jί"�r\�������2(>���+X�,�MF�PeC:)ΥC�j\����~�#���?����.@��F�/	��rq_�9�gOUu�h@Cڞ�e��	��gՒ*��[�����z��4�È�	��61,O���O�6�0��a�1���
�ֿvđ�	d�p/�"ї��LA��yc{�߮��/ċ���p�r9���|4�\��8�����Sz��AE��4Nr�������ko�:����4�M�d�	����9?Y�ʐgE��k�6�G"��
�2�D�E=�䃯����4����-aOK.,���3G�����zR���G��,�e"pKn�au|z4o�}��A�o\�?��k�)��Bp�r�=�������݀�G���P:��|��|st��|���66y�vZ!�}��:�]a�a<ӵ*��%�qN>g.M=@�?
�g�9�۾<�_5�Й�����\6cԎ�>���h�;��07�C�7�`�T>/�2톕�p�U�	��㹄7Q� �O��������#�2vUc�N�;Z�/��8
����4�¡��F)���6���R=}�E�j��1X(f5 ٪����v�ݚ	�LƏ������J�Iy�Щ��^���JL�|e��%�~�D�.�ː�c���Y���Q��A��*�Q=M�|.ҳ��	_�p&�-PmWّRr'c�[��1fԸ����S���bd;������q�J #���n�:	{�D��>���Y�TP��E��`(�]o�Q`6簍o`q�D�
S��k�]�c�{�7�u��֭��V�,�߲jC�ismل���ЖU�+�l� `9*u���_ˆu�Zp�����DizXcK�6������e�1�)0��H�o����<?������ASu��9 %+X<��0S�����< ���A��5_�t��[����R�q�_�Z��ey�?{/����ض��b��	�əd5*��K#�h�c��ԗN��KS�h��B�)F��hP#���yD�+��d���m�<���]��p���}��m�7FJ>��M� H����vq⻳��J逇��K��Q셜;EX�/���+S��g�9'N��J�~M��	�@����@^����V�Z���Z/�N�epW�̩�e�{�ׅ�~YUܓS�ى4��#'���bs/�2�˫Y�7Ȥچ�]/��}�+{�����āc�`�V錃��ћ���������,r��M�s�g!eqQ��|%	!%ov3	�fF�]_#i���<�^{.����_N�zg�D$��oB!�zj�a���i�ґm���IK���5�A����5�;K�o�����ٶSX=TfۄI�
l�{ӂdי�:xܞ�������Z�\���v3t�.���3�a����v�,2�8�E�Z���c\���x���M1���+#�ާ?�p^��"�LpG1Q�4PØ�D�EkG��ԛz�}Wt��X��#ޘ:ax��uU��)���+��S��/��A@v}`1SFM����e4�{��&(�h�����LL�{�Im��O3���J3ٚ��y�r��� q1�XZv�*s0��2Ly[� X��X]�zH��<��]���3X:�ܫ:Cf� x<��T�n�����3�B.�~n�#Z�����!ND/,�m,�:���u��ԓ �t5�i؇�w�R��e�%5ǩ��҇��΢����]�_�!�O�х�oWc�(W�۠B3�[*��Fr5���c�n �k�:G+fn=0v�Bw�|�� `j��[��!dL��{9��E⢔r�zb|Sʞbՠ�Ktț����Hxb%>�ح��'�B�]u_p�Q�F���S�h��[�9@X�i������m?��
��J@+33c���vb�}�1��A'x���K��ێF��0���h��PP8�{ڼN�M\{0��m��8�������0��J~���P�r���t�P@MT��;b"C��+A�N��M��c뿌���G+K8/5Olx�D<��p� �N��G��O�Q��O��}��?<��k{�FVV�zvUw��+5K�\eǊݝWZ����N@����)���)�?$i���	$��L�:t�al�d{U���]�r'i��%��A<s��b����W�(�i���{�F�9~���C����k8pQ��o�4 ���.�b�Dx?��T H4� �U}O�S�>���B���tn��� �0���j;�%�VS�ib��K`I ����T`r���v^IL,"��2�ۊ��j���G��)�{�[0�:�@0�d����i�����k[(ON��V[؞�?y�\Yi�j�\��tʱ]�1��Ȩ�zL��[h§ �PHd*Q��C3)��r�'Fu f���*�Ն������t��e�<�B�s*O�zm�XkG���;��	�g�{�@�(k8E�63OpoL�����iz߾s&7c�K:�v(�˯G�Pb�7(pf�T���ҍv�Qe�יn'!_)����<�.��.��r�+���в[�
�K������Zd(�(tt�Ԁ`^`_�g3�Y�l��2f�z�?�vS���N���c����ž��]��}��[��k�r_{�N�Zfz���;c_�+������E��X���3��
�$,��L~6��u9D�G=�t�&;�(E*���?����kX	�w�m��W)�f�:$��H���џO؆Y�NEJ쫛�����@����K������6�Tb� ��3F�n���8��.r)"����g�٠v�~�s�.��.J�n(���ϙ�����ԁ�b��E vO�8%�d��C�+���Y�o��l��0
��r��W�����<h#�t+���-���n�M�ܟwB��3��X�A+t;�6h��=�V&7�>'x�Ʉ�PEɿ�����gN
O��i��� k���E+�wIJ҉�΀�;�&;�τf>�9#ˤ�D�<�"Vm�FgV'(�9ٛ.�F�Mו˜	�U�p�0CN	�%	�M6$��>R���Mf����I|�k+�D��]��)>��B�Hhc�E��L0�˥��ҷK#o���������E���7�r�ܠ@�	���C�8y�j�v���9�#�c�V!je��:���A�W���SlsSUȳ�ݡ���ŴTz�j""����L<4#(˜���[ia��ʠ��aw�s����)U�h�z{���IUPހ�QFb����{#7��:o6�?�z�������7?&��.�:��y�M�hb�V)	�0��C�\<F��r�go�j�a�b���_�3�V��&�;�3?��ˌ��EYl�l�żM�:'Cո�#�� Ȇn|)��pwM�;���Lw�k��Q3Wt�L�H�MA�1�{���Q�f;�A#��l�.�è�ֳ£p���:�a&I���G��v��A�<�����lxx���t����+PUM������X&�}�,1����ۄ�j���5>δ�+rmV�,7�����j+0�u\����NQ��^Ӛ}��Pμ���U��y�oq\�S�{���ɋ2`۟M1�9��ѹ����r��p�a�"<�'V���̬k@�>?*�� Bx�^��@cC٘��������H�f��&��(smͫ;��U�����Þ�]����wI�B��k2��$eD�Dx���<Z�q��n}��*}CMn\��&IR�.�@ݰ=;< s԰�`�����Br�]X�.	H,�I-K�9\��wj*��]ޛ <ͥJ�V��D]d]����L�s_��D��<D+T�_|2.�K��?N����g�|�.����	hPplm]锋x𻡗��\*��+�=m��(� 2�e�O��,ݔ �8��%�I�FL����LV��b���9W~�Yj���ؕ�[�O]A��>��`��z|�,9x�0��)��Fb�x`�>����b���qy�U'I��AX<h�A!�;�QmW��:�Q:�y���ib��ۍ*�:u�f� y��I
����S?�:���%{�������T�Y ��YrD<|�816Qj�Z�4�1�D��]�ք'��!C�ć@eۦ����o�ٜ���ͩc��q/툡9�V^{�5c�v��v�X���j2fk}�������m!�Y�[�ftf��~D��=}Q_r7D[9�c��\M���8M�"�$C��ѓXq�g�U�J�v�x�����:�c�n��\����(�a�+��"������� 4��k`��`��!���[��6���<8,�UЕ�����_4tQӹ���n��*����R�����=)��E=y��W����
Dn`@��>T��1�k��QC}M���l��M�-0��3s4?���A?�kEF��� ��(��S�,񰞺��˲��W��O��ު�q�F�dK\�O���Y"�
<g2����a���R�!5V�eˊ���6f�.���|F���vU��b����|��.}N�Q-�JPt�~ǒ�\������c��y�Rmn�Vs�ȶ�|���'���r�ȋ�j��"����P���`<-p�a��������#:����988r^��/��ot-�W�RJ��P�3�f@Ŭ�$5�c:�e ��w�[�.$��L�7��,/�L�����1� %J�UP[{� � *ph %����D���&���i縆�{�ћ7>�9!�4��%��6�^ؼ|�J�S��;�I�<���In#rs9`z��ʺ�8d�Sz~�r�.������1�����DQF�q� ���Q��6�w���ζ^�\��-�zu�h�w7�MU����Y ��NƩL���:F�z�x$�Fd?�+�if̳��^~���[P#MV-ȣ�x�c�O�ޣ0�/Ԧ9��1�z���a,���Z(������DK�K�"�� �C�5
�+��}�*�QK*��o�xSW���8�ֲm;���}�5Ӻ���YMV*4�Ȕ��Q�	��0M���q�6[J���\�-�Gׯ2LvH�����0A��#;cZqeI<��Aa�O,F��u��6��-lk��DY�*�Y�l�h`º�?�p]|������y.��{�X�*�c�z�\\��������o�����|7P"�w4��#L��G<�;�"�y�h��	�b�F�]Ì�w��xW���/.��W/x�{���N�+p� 9)���vf��¯��1nL�8�]��/�3w!|O��3����X��U|��^�2��w�4�1I_�l�e�@�S~���[����͊~��������'��\�bG�X6^��9�]�-��EO-7��XC�r!���+4�����G�P~I� �����&��!���a����\FH2
�5��c���ԃx������#�I�vL��o�*�_���%$���	c(V������R����g���c��/��ϥ�FY���5}�r�pꤪ���73-�����G]C�TH�@�(�
ƌ����Q�& ����)A������=v9`�g
�!P�i_��`���/GkǪn�@'�C_��5r�$"wzx���8M#2qs�_u4v�d��37�5�&ހ�%� ���L��h��;�L;�H�ŨނH��w>�X��GL�w6�����eV�!���x,�F|�iP@�����_p.� �$b��$���+����`%Qo@?�7Y[<ņi����W"A��E��F��2��)��|vL;^T�[S�k��M���\�?��-��ᇣJuU�0e7������l�_0��:X�.�[:.s(�,���3Nw�i�$"���7�:M�틠�#�
��R�Er�h�5K���%�EBu�9��$��!i���{ŵc��N���Z�coE�J2�a)D���`�Ks�1*�j��sǊ�����(^�v��Y�ͭ�h��40�<���<���hݵ̎���@s�H��)lca^�z��G�5�`���X̚P�q,p��Z뮍s~�~(yj��A�:1!<p��ݫ���e�O.�+L�tH�.ʎ�����ͦ��B-8M'E�ֶ]���Ǟ��U�����=��~cV6�������{7�%B�����s�3�"�b���ٓx��y�BT�$$3���tE�V���}��S�ňHs�<�^�һ�X'�t�6U̜�a��*�8Y%��Ɨ�]��֮�7g}��E*���1����f�ˑ�eݩT� �l@t ��P���m;��3�C���:���<�<�� yz�|�,wUڨ5�p8`��X���m�Erեғ����)P� 3C�x�c����z݋���h&�A�Y^�4���9q���]{�|�a�����?U?nH�����Vz�!U�~s~�=�;q˰��=�[���l�S�N
�I����Bf��i���Z�>hvd:ZH0�b�R�J�Q�畢��K*	O!?@)n��{��:q;�o4�*�2U�f3c���<�c�ݷ`���(�=���E�S�j��X�,	��d�g_���1_��+�d�]�5%.��7���oC�`���e���= �G��,�I�$�D�WnBI��^L� Lпw�R�Vx�h���q2�Q?e�n�/�m��)����]7��y�_�����0�I����9"�VpKS?���K�|���vHA(�\
[E���6�R�N�C!;�N�uZI`m��[��Ԛ��.#Cr�E˔��e���/�HYܾ�-%I?�~���F��m-�hڽt��ju��eR�i�ځ�ॏk���Ĭ,��p�7���B��i�!��y�6�?_�!�&�6ZP��"����R��[y?��j.�UI�&\��T�/Ct`�ߔ[O�h�#;M���L-IAus���+����O�X�f����0
�8�屶:p2a1x����g���B��L�n�P�c�����7������$2텲�Q3��,k�i�ڷVdh�����l��l^�	��a
��xb�	)NY�y�� ��
�a�=M�t��/9M$ӗ�ޯU�]� �/�N��o�e"�n�~>�
U�U�M�{�C?Û�<�t�����(�<Qo�sU�Zv ����6�
B�Y���I���L�X�0�.Hz]#�@�;�u�e�i����}b܉�N��`��;���4��s)l�`��z��V>�"�0(�gŔΖ�ݛ,�mm`y3{�Z�C�,aEnҹ��Ņ��o�L � ��}�;MKR���)��n�Ǳ>��K;x��2��+�s��: ��D8�W-.Ջ�*<�~`}qD�Dه�y��'h�����fcC��~?���@o�e��uͩr�"I�R�e�g��ᐈ��uS��(���*:D��]���.�F�t�Rq9;�;�H�ɳ��,�I�����S'�ȓ��0H�S�lY�*)���KWe��q}��C�,M�AR苁&��ocxZ��WN�@��:��Kn�VgO��x�ZcV,}v@�)�Oi�~26����(C���8}Y3N��v��g2� � �e!�4�$���c��hm���o�l��>y�8vKC8 ��3��?��[lZ��Ly3��#�k��
�^�'\���Y�
T����xouW}h��A�댛�Py蓮\���$�c�߫te�\����%#�k��Z?YsvI6M�$j���-Cc_ȸ(m)󘟝�T�K�?�|�F-��ަ���~�
*�ZB��r�/������\kl�S31�еk���F�j*��þx��n�Ī�.
����Y=��V�!��~���ně��F��8/������ݏɎ�8r!;��PX�� �"(�s�~��^hg���P��؀���S}ԏ@����tx�����F�WV�4}})5I����E!5�����Ulut�+�
�������j@w�j^�q�r�Vpl������j^��A���Ȭ͏c;4-`D���ʉ�j[	$����H0�����Z�X4&w�+:۪�E>�$ϙM�ؑ�25`�gԈ?K��9�q_�g��쓒�~�y]�S�:���RGB���_��Zi�/a��"+�K����TRE���sXaI����)�T����{�=�.�Bs.~s�-�Oኧ�N�:�a���0��jR!��t�hQ�f�J��+�?]��BJ�+��&D�l2@z�,�b�X�Q�Y��0v`Zg�j|��T�������9��1:r
ޯ=�$sԇ�9��,��Y3����5/�D5��[=n�R�J(#�ۓ]������A���DA��1�UI��u�e)�5������r��U���m���� ޷�(��C-��iv�V5/IVN[v-5@�c!Q�Z��JfL��x߯<�R�j�z�	��?|b����#~=�Z!�ޥ��������$���+�w�hZ����E��d�D�l�-d�Ԕ5��Љ���&��H�ڄZ1�1�s�ُ��P��`����-�4��sJUC��lF>��(��z�,Uou�' ��K� W��/R���'2|�n�Io���,�we�<��*[Nx���ʪ?�@���s��hF�æaf2�?�&+�Q��� ���.���Nω2"������Ò(S��1�������`���R�g���W��C 3L14���4F�J��IrP5�*����V�4sD��3��a�V�	H�빖�}\�l����̒+�3��v���eK�T�I�k�����@���tVn�0� U�Y�d��%��}F"h:��Y'��!�<�[�շ��`��RP��˧���[t�O�������ݼ�mj����0W� A�׉ʻ"��D���}V�(��}�X}&�I��y�*v��Px@V�%�Y}]��$4 �)@�4~���o=N�羫[��%�|d%�G�Kcs��<2�5��Xو\\[�ސCܵ����&Š������$�A���=�p�*H��/Z4k	jR1{���f�����D��җ	�e��\7�@H�����	�	�S))�,I�F�:�4�᠙���E謃��K�\�ߘ��Mf�ֱF_�S��ġ#E=�O�>��M�0Hk��.P�ț�@��A� 7f,�K�+��{6l��k�df(�u�y����`#�
Q��݁�Ӫ�� q�`��n���ӷթ�ͯ���b�{J$=�ڳE�af5 1�4�0�<3%V�v�+�M<���$�2�V���-��};������2k��_іR�C�!k�^Nq���:9`����>�Wĵ�Oq�{�~��B���lp�J�^��
��%Tb�!�#w�e.j����o{G%lG�_z�,@�t7���V�ܘ���R®���	�/P�R�>���Le��"��M��CM���q ��s��+����p��QhD)-�墺�M���T�Rk#������[�K��I8�b�K0	�VU5{u�+H�D�b3f*�I��0OXrDG�"��"#@��;n�Y4^1y���9؜�m�A5Υ
�}$b�k�����u�@TNb���V
� '���h�>�+�}k=zC�bC�6N�p�`��mЄ�`Ib�+Z������L��,jBX����4M�6$�C>�`�O��	��P�
Z���E�~֕%.��HY�UR
bW!1��a�r6M9cğ6��&wJn��E�l�c �2�����.�AS�{��H�13���Q2w=<�
�`��l���q���!"ɓ jf?�"m|�Ne�j��^�O�D1�>���U˦�ԌMY4]���N#�'DR������0V[�p�cjsW��ĺ���)�7������ �
���''l�({�{�;�s�֚h�aC�t�i�L���������C�J��1��?M�ËK?���Z��8�ܬ���?i�Cv��Q��J���u��3@=��'�T��e��X��Q��`$7ȡ�SlǇp���vS�h�7�F9�'�5/wI��*��L��-O�KDRu[��#�	���u���u�֭x�-�����bJ6�(��zm��	���ʢn��>Sp`�(������}��8�4Z�m{��YH��=>�Q�]U��a���.������w.����ۉd'
A��	x�1g�j�6)��X��1(��ꅸ��&?�*H�PW�%���pLz�vnD�p0�'8԰(�L����:�<���S%�Jk� ��i�oͼ�W׀���0�˰Av3�QRrD�8/vR���. N*�5�,7y:Y� P��˧ҏ���*��������-rm��~�i�
9F7��@�q���y^�z�R�]��N}}4aim�9NڅmB�����5���t�h㒞���d�=�e��4-F��[�)����n�#a�A}�T
.��*N��&w�I�a���N-�A�l�I���	���=�~�}	]O}:�dW�D4d�r�JX2��zG5�Y��Q��)��~�r���dz�ɓ�O�h�����J�s�Y����`�U��N�`.��Ovj��t)7�
a�p����کӌ��������<�r2���x��.����;W �/���O�i�RsF�%{�TQd�NV��������D^�vIU�7W���.-^C���E�Iӏ�b��Kj*F�i ��_���ѡj]@I�SP�c��P�e���B`���*&*�X��#��)Ym5?oR����h��r��ȇ��?�#,i"��Q�@�0����uA�����NX�gQ�(�ٱ��N�o������0(��a�uX�Y�㥇2���a_b`����sӮ�������g��&� �����Y��Oאg�M8�~��a��Ɗ�,X?�6�[�@�Ă����DJ� �u<=����˴�D�W�#{��9$��JgMVʆe�!܂��%�ZJq�Dl ���%8�JZ�D���✮�/ �q����Q��-����5 ��d��j�]�(\�=Q�w.�f]�_��f�S�-}z<�)@禉�5��֋�:fd�����uW�^����SB��\�!�a��Nհb\�HK9�B8�����%���	]�%�H,�@V,W�l�+�L����4������f�*�^W�V�a��]*���X1N�y��d4>�=�l��ȱC�j�*�Q?�S
�V$�jZ����m��VP��S�n9�i�i��g,������v���2�$�[=z��3I��5��Ӻ�#.�Ppcc�l9-	��Rg�T�� WC�aj��|��I�?��!��`s�N�*�Y��3Rcc��Z9LM��ˮt^���WH+��p7�iR*����0ڬQ㽦�����Kt�o�/��o�HȅU�� q=ڶA�J����$h�>�0�V�^�p�>���T�����2~k2���Hf�i�u8��;�������^{XM���l孔�Q�����v�@��r0_^�\<������s}%-���������*Q�͔���a6Q@��[\AO�U�䶇�Q_Z��U�߯��]n�=�l�G�e�J�T��~�ӎEU��@c��[<�C����M����T���Hp[w���-W� F�$�&+�%��T�T?ވiK� 'Е
OX��{�u_)���z9�y�����e *9	 �8w�si�U���*�e����Ȣ�����~�M��Ei;����q�x��oHR#�}��fZX��؂
�8[:��t	�!V;�Fu)Bq3��+��H	���/��%�\p;7� 8S�؋n2�:W��F?��IM�Y)�'n�źTTKn���5�eI�`s��,4�f����Bn�j���T��3YR��=)�UM]H���� N�a��%v� �}W��`�Љo�:���b�ef�z��vk6���><�r7tXP5S���������!�Eg4c]���b��z���Z��c�i����J�O�T�b��񺙕�m?E���(d�_��?�s?{9� �)���FȔ�I����\�AI�����}�A��/�\��{�)y�԰ڄi���K4��Y�0�#@��_�"���x�Z�Ī?"�+�.���.эkE���Rq�D��F�$#vd�xEEw���+7}2�H[�[I��"�׶\|�A��\�^��N�gz(�Q��=>g.�cpF�&�M�N�DrC�����M<g��tb�Op��J�%�,Z2���IE"o00!_^WJ��x�%z�[ܶ���2,B����珪��?U��C2W�z����W�M���s�F�R�t?���Embi��˸�&y=W�� U��T�RZ.�ל����,T��:)ގT��_�
���;c�o�8;�1:N����q�4BZ��)Si[`R\'������PT��֟�"/�t]�ʾ���+���CH���� �x������ת=����gw���=�&�蕰䲱�cp0�;���f����6|�B��'�#��f+LSSqL�;$Q�����~3�K�k��ը���q���GD��f���7*��Qgv�+��^h��i~X|$h's��#Q/T�B��1���}t
��ʵڊ���(�h���zB�)��D�8�����xh�tp����r�����Y�k"&��J5�����vA���ۮ��&!�L���A��I'��6��E����tʥ�@w��4��(�Q#�����$� q圍��i2ߙ�n�u��|{Y��7�xb>�l{�B�8���!j}7f�@���8]7��6�q�J�0R����������$����E�"du0���b�C?�>bhߒ��CnW��(��YѻX��6j�uYBM���BG$���0���L/f-�W��%��hJ��>�����ʽDĽ�Њ=���F�G@bWQu �e_t�.z�3��d���63
~�w'�fOo���n3b�1gǻz��لx�NiA����ݢ�X�T�r�S�RQ��>����`M��6�t-4 s��F��5JYOh�@9��ꔑt��WQ���;���L��!�]�OM��K`Hs���ABW0�D���C�#�����4Q���*@[@�rqw�
+M�,5]ْ�I�����Nb$�~����.Ƥ<j~#����W��3Q����@�G�ki���"~�]��I�P�&�6���#�}���v}>6jm�i�����b��Q��B��VW-q}Ss59�X�Q�%��i	N,H��hD��)��F���?�2u�I9lf� 9i��ȸ3x�Dr�I���?���ۉ�s�W�A�kF�5a޹h#�w�L0��b�9�n��2�#ud�UC�=e	Q�$Q	sk�/�0ɛSF�����NrR�ɡ��0{��rf�N�9��E�@�0�:�0`�/cQgi��\����
u��W�k���:�7��?�*���Cѓu�Jr�]�]��y&�'A�'s�[�z�d�QX�-�6��Tc#ъ�����q�PE���5gn����e~N��K��l�����
>�/� ɿ����H�a)����W����dF}_j
 �F���侹v��-�rD�i$@�����43�.g���6�H���E|��
�i�M\U!t�	��6����e���ҟ8~-[E���,����*Yy��7������/��T���K���9"�n�C��#�V�4F��a�:�4E�P��m�����>���N����Ĉ�e�
�=$��W��8N�U���Q��s;�t�;;?��NWj�@ ^X�H����5Ogwf��3a0M!��d�bv�<��-��������/*
J�r��'_$Z�W>	%� � �{YyǶ�U�A�W�3k��U��J�N�	:��)�Z��F�XX������G��rwº%�N0;�eO+	�#y/�|�C\���GEw�^�^��?5zJr����3Ef��LD2�1#*�Rڠl�L�		on��Iب��	��h�&�v�h���D^WN��hϴ)���<½-�7&+|S���Vģ5��!�}.��7�h'��f<���X���`F��}���\�Z�%����:g��jê�c��E�H�E+-�_mV~	�O���v�(��"M&��Ч% ���|zɸi%um���ZAb˴�.hf�~ĳ��{�9c��L� +�)��G%�c� ���74p�7ȅt	���!Z��O"���4ǧ�q�!��}ea�f�m��u�P穖�C�*���sEk�g�0��#�<kڭUa��Ӡ�i��=�$mqD�B���6f�y�L3T�i��6�!�@��=�3F��-��!ɨޡB�+L�����9��(��X
�d����6MB� <�7�pW8������3*ϻNF�n/�Bآ����y��Y�a��Վ��xH桵B�y��eȫ�|��pHR�#�|8k�pw�@ao�WqIga���<$��e�5g���i1�?��H���<w���(��'넴���c�i��V��ud7)�w��E�� �f���)�aL}����bf���;�u��'�C����l�n�9��ʻ]�WFint޼Z�[��1p���z<�fȗ�`$��U�!?k'���e�����1F���L��^�J�� uN0�W;���8g�xu�+�v��J��i�ɠ_�����ۊ��% R�n�D����.� Gv��&[�Ye���b�ݺ�¨�eޡ��>�ث
X��OO!�-0�d�kO;��|k#R����/���)v��V;re ���4f���dq)h@H��E��ӂ8���~9���(�h��Q�hB�l���bK
r����/=���G�%�c�c���+��h��fwVjm�ztp'
J�r����,�M?5�&\>9 
o��H3���(2�0vߑ'ʮ����4�%��ǣp�r�)9]XS�%�[Xi�T\oF��<�b��uSDV2pI��"�Po�ѓ�.���T�v�3�����w�E:�c����h�����%ZƔ�+�8C���ǐ�*ҿ� �_;:�%���6���j78U���r��u�����;hl��=ǀB_��ę&\�0^a�s�ȴ�����[:�W����V�%��4d��f�L>�y�h�E6�?���6�:Ÿ�-T��z�!.5؎�yJ�� �ۭ��-���Ǌ�q  ?;��[ ����M�:ul��#E���g����(��/`��^*�G����T�BaI-�0��pDr�jxxx�Qɋ��
�5�Vh%>ᚗ�����K肔���B6�Et1#�w��=c�$B�����eYK
Z�U��s���^Mr�f���� �NIͣAW�z�Vj�I��f}�Ԓ��C��6��.��NO�;��Q��xtЕ�>"���N����q�r�ɖe48�~tePz�(���z�rv[�U�^m��x=q�	�����G�Z���&
�avNF(�M��&�,>Xּ4�w���9G�!pW xJ__ �I���=���(�F� 6�Aa?�M#
��;c0�z�ͻ%�%��&XO��?y{��@D�K��K���8������dO*C����n=B�T>�98��cN���2)����ʟ��A�_b����:N�� T	�����ݴa>5%sji���;���4 9{����t���\�P��2�qǄ���*�L�FXD+`T�n�|��44�B'(}�l*��լ�G�\x�"w�B��*YǙ�#�Q*��/�_�̭�B����D����,��R��?B��F��,&��/I_�z>LI�3b��H��䓛o� �ڧ�n
�y_M\��>�],����6��K��� =BJڊMH#���w��϶ �/�e�����7Os]���=� �MB]�"��p �&%d))�!z��Q����?%(Ӻd1*UE���[}w��b�l{NŌ/��Z���*��٫@g�\���8��y���ܐ�1ˤ�]�r����mQ=nKFHn�H��[T8X
��(�������1z`��M�-����FŒ�!�����w�>*I¾&�Pi�³p�å�˄W����*���4��&g�R�'�m/=^\@�����4�ֻ@,[��d��PB��� �&l�B��{ٴz�E!PȜ�L��en�@:��bo�+v����0`�	���Pvߔ8�|ޓ��	��<���5�r��]�:��6vB�/�a4M~nF) h�x�`�O�X���ǎ7z��S뜧^@�?m[���r�J*C�oA�.�z���ILfJ�~�P�aȥ��e�^���$a�����M��{���	f��7m���.[���?G�0������LF=��o�B�`���0��,��c�vB�'�鿣wO��;�X�(K?�F��KӚF�m;����w*.��ް-�صH#��m*���d����%�葃���x��+�/J��":�~�ag�\E���,<M�G�%�`&�?��|��O�G�IMc��j�ۋl��Đ�ߗ�^��bq�DpfI�7">���t�JC�����е���RmH�;�d^n�qi���W�ެ"��1��f N9N#��#�<�h�T[��-g}I�-���0-ՔVj��Q���m�G
S�-zm���mxՅ!Ў�U�Qa:6�>R����qȞN��`�i���v>���h*�*- ;�2X4���$��t�q6U����f