��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4dտf+����ؐ��7&Qa�z���m�ࠧ��3`����8s�@M�4�s~��B��h����&����YND��b��1Ü�(_^�[: Е'�GK���c����i�};<���k�.j1���a�����e}�PN��_�8���>=6�eK/L(�#�S0��C?v�>�-}闌�=��b�7��-6��ָ�	���8/8bWbR�рI�5�� �!VX�`�H��-jw�_�W �T�2��@�w�E�ў����q��Jx*YiEW�f�<�P^���hሔ]�:&"u�Xg�ծP��齖zd���u`�l6d�zh�L�Z�͙���z)���i2NR��uoݕ�W�y�U3)}�C����7�g��H+�X��6��e�f
��,���@2��v>P�ۉ+�\��@v��$%]�+�����M#��.-6`�F�ǹ���X�=m2����v�]���[�_>Z#�2�VLXW9�{���6j���r<w5 ���h�^���O4��0�;rw0�1Hb�&�q�	@�ˉ�9Ȧ��|b�pJr��^X�]�dG��)����<��"߹H#0�.b!�ޏ�
1ir�g}��u�L��Ӆ2.zb��pY�݁%��`���>��}���.�#3�e�(���*���Ѫ�����6j�S�&��vv�3���J���F�h;{#���ql���[*������b��:xh^"/��D�����3S (�G�xC��èv/�n�b����W�|V�,�\C�%������1%�,�Y���T3�W5u��J����ډ�E�&��z�
K�� -�8b�\�T�0&��*�Nk2�N�0��M:�;z�bӾ�|����-��փ=���[����(drl��B#�#��%J
�ͯ5ׅK՛�Pe�/^2�'^25�Xs��6�1�:��8	��ex\�Q�m5�oL�gzK��P/X΢F��~�z��c	y)�:�9�-������#<a�x�XⲒ$�3؂�9�����he��di^h�8����S�3�����2��xko����}����& 1,�������mM�XW�M����G�,�fMA8s��LQ$d�?���p��#P�t�e�a{��6��PD]weh�0�*Ӻ����6_FĜ�X��#`�oV��V�+�����B�tC��x�#�KT��A��a ��^�uNoU�N��	"�mH�)/IǬ��n�hU��r_T¹�	�9;]T/��������-��>�5�\�\e�L��X��ː���l�u��f����\y����N�[S�n�:b����(�P�"]<�
DkJ�Lɓ'���Ω������eV@*
)��O�!eo�����<f��^!2�TK)�K@]����#�,ճ�,R�������,5��x� 5��A���36��~��?ɲv�[yɕ�M��0<��ɋ�/?�f�P�7�����%���/"��7���%2B����>�r�8��%aި*�ѳE����s�<�t�CH��9�Œ���e�)�k*��B�� ΰ�yW���0��z���!=�4���� u�������O)����c^�ĥs�v-�e�I��a�x&�o�+AO4k0H7'>���.��l<\�?��?Ԑ^)�9�&̘�H��[��q?PN��`��+3�ȫ�4|��U!_ ��|N,�R_�Ӂ\F�������[� $A<~�O�.��X�o?8�y��)@m��/7�e$���U��A�
U
��\�M3�]�n��t�8�Qs!w��m��é��T��q�l�؏��j>�Wȓ2
:�{9R���^�vJeH5�?��� c�d�,��?VK'�23�n�Xc���G}97zST�ﱚĸ.x;"9m��9�[�+�g��� ������%J���>Gx��J��e�_�ɽ %���k�W}��E]�*�s�PԆw���k3WLN|���n���:�\���v29x�1�=86)�,X70����N��~OW(��F�t���V�̩��'1���Y�vj�~!��<8��^&)`�������_���� ��	̴�:�ucR��/.<� ]�s�kAo�Z�<��v����= ��� �U��ŋ��+M`��MW�=�;Ϗ�3������b.dk�����A�^�k���~:L9�%�:3�FX2�k,ƺ�F�ny����f���;��`��]xzUF�y�"�E ��_�� �'P{ �,%�h�|0mu�P���3)S�mo-�:=D�%���J�n&��s�ޏ/A�c�.�|���u�����%�ӀM�Y�*�Ȃî?�Y9���;8�U�0Y#j0������ĺ^LY���MR����<�0b��W�$W���MN�S)~hD İ;��-V��w���8��, !r��)0��Ϟf���;��1��ʗ�[�9�3���i燞�(䌅���w�;��poS�w�|6M��Hg�>�@Ē�]���N���s�'Oł�j����Y	d���31�p�Iw�c�,+J���.X.��j@h��1���݃�S�)��x(kC:��R.Q����xK�q\7apBx�$�^��T�9�{p�R�H��㟔��E�	����J���uM�e^��m��g�R�|$`�>�N�!1_�"8R�c�~
{�iV/��ma9K u�̢5vԕx��V��tJhq7��!΍�.����|@	ϔ�����R/�����������02���.����*�G�h�6Xu�n�`�tu��FJ�Ջ�ק�:���_�n䠒���9��<w/	�Ί���v�^$J	�g����2RG)�ٵ��h�F8a����O
I7(X�~3N�ڐZ:�|��|_i v�^�H��Q@bz&��=DK�_�nx�5�AMJ�
1hvB���F�}"�*� -��rx۞��YӒ[biWqu�چ��KI��|�w�#rJ+��|4X��*̿^q�V:2H�� fc��U����광c���K��\�2���v�ȣ�.ہ7m2��T��s�`���lg��6�T�ZP�pF�
*Қ��U��8�UD�?�MUx�a3sl�}XTw��ž�t\Cg6��,�3zL�.kх`M���&�Q��u~y�𿋉�����N}Z�?�x��> �D�1\���yb�w����S�q	];�8){�k��wt�@ۊ��xJ����`�=����`�&��7�Ÿ�9=�b�_D���j'����@r8=�Z�zT�z�qDd�XFU�Q�L���lE��T%B����q28��7\������2����y|�t�[{��>7�������4�2OF�. Ul�?l����j:I4[��ʰ�
���5얘DJ��B=QWw�{6=�����z�U<��*���߁}z_�Y�x�W�C�_� ~�^ؖw���;���7#uK(��+���"�ꧣ7{&Q�_{#֒J��`��k��:h�mi��N�:nk�����~L�Z|�L��D+ט�<�,0�P6nF��O4Ku߰��Eti�Vƀ�X'41]`�̎`��w ��?��N��~���ĝ����MM������0��r�Q��J�H6��`2��S�$Ӣ��́\?�O��+���6,��h��}���5)�eؐ�si�>#�*��J>���w�q;O �˵(fH��<��@m0|tS��P�n;�����{�֗��t珜|�]��u�X����7l���=l��P�:a Y�YGi���^�UmV�7]���%�<&D�]�9q�J���}M��d:����3�߆P��*w6wWMO0eO7PaͩyFڙ�X�=W�8������@�K�rpp6L
p �����C��]|M�F��*=d ��G�m��W��ݐ0현e`n[ K���3��A���f�n� [;{?8��a��:d���Y�-�3�u0Kf5s�{Q�#�m�Գ�&��l�	�d�;u�h�v���tRVϟªdW&H�oL]�L�Ģ���Ai�>�R�Z%H����J�;w���	�J.�������o�@w���%�P/|�fmg�U��I=�ױ�0�V�w�P��mٽk��fE?~v����FJ��T����i�a�]�#)>-ze�d/*����LlE��L�5I��G6���(��+D���2,�{�Q)�wxy Y����~XA��a�2�Ρ�_޺�g��G+�Ӧ(z&��M���;�7�s��;ݰ�!e�P�]��a��o�D�@��IP�W����UV�d$��/����] Y��5o�	��O�k�&R�}<'���m��1I�_���^�:����j¹盦���3B�v((q(�ɝ�p"m�������9���X�=�8�r;�6�2��}�k���g�3���,���x.�Ly�E&4��J�<2�O�CAA����J��@��`��\�)�Պ[��38�lT��ܳ�o�	k��k��E��j��xDn�8�3�P�|#��jRu-g���I�Y�┆�3(ւ'ɮ������M��۳���|�Iy@��Mw��q�*(�:rB9�Dt^��&� X`��������B�ZP
>�