��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�������@�wA�>��)�A�����F�����l��`�0��#[�Sj��2u!�b����@B���`L�����o����d y��_Q�LAn���'[����H��J���:C'���+Wq�>�Ԩ�"J��v��쌢0��d3K`ۗ������T��LRR�+�Z
���{<�e7��>�Q���Q<�Q�9i�0�\��8�M������
���kc
�*�b�����}��� -��j6"��dB|�#�8��ͯ-�E�Y���;YD;�}� 6�I(��h�X�"`��B�|:�;VS�z� }���ҙ3�Ev�/�Gr#{5mPc&������_x�e�\�=M#ns��YpV��NkЏ;j�i��Z�c��a%?�l�i#�?�Q˗8�}�٢,SUz�deDo`j5E�j</�/���K�#�@��*{�둥���ۓJv�����%v�Ƽ��;��{��e懮4,>k�+�hŗ�Ŋ�p\v��t���pC���	q�G�'V�;�x�'j�᷎�S^�]�4a��_
����]zQ��a��G[�]�Z��e_�-�'���>��?4@u$�"�ށ�J�����>l�������q)�c?TK��ȥ]F�G�:Ym�w��[�pH���6� �_�aC`G��~��DBH�R�@i[)��,$�L#j��W�?!Q��:��Q�U��C����`ǚ"�_Y�q/�N�F�AJ��Mn�������k�CR���@hS44(�3�\�;������ox�((n�y��b=�Ѻ!~OC��dË"6M	��s7�K {��v^��ѻ
��>�1�� �� <5I83��}�[>�O����bG��E�l�v�bK�2�!�2���a]:K~�r�~��F!C��Om�'�hzDx��`�{A[��*Ko5َ��YP�y��L��k� ���ٻ�T�jk��h��%����҈���ƥ ���5L��!�8\�3C-�9\梦g�l�I<\/��J��iD�Pr^�)~�����cr���4���|[���Jv�3X^~����a@�f���얔�Ё�kb��"p\]��]����������#�l^}N��v#�p�'^� �P��m�JP�	�P$��q��D�����݌�.`:SxA�b ��M�VH��z�]�,��0v5Z�A�|z2"1�E��r������r�G"�3��>�1H��?o�旸\\F���1����۽|r��/۞�S:�p���S���^Zp�d3�\TN�~�Y���m>���i�}!�"?���ү�;���"�tr3~������4b0��iz�@�_���C�ݤ�a�X�:�,+��vRn��e&�M�����<�����Ew�V_;Ka���A?���ݖ�hK=ħX��v#�2�^�ؘ(���!�{�憴��/��yN��0��\.$y}�u����Z]9��(7�?��w���8)�`/��t5�o�a�b'p��\���VQ�S����i�_
���H�a�PJ��Y���y��C��Q�0�}/X%�����(��X�lyt*e�Xw�[J{���[�-a���pw�͜���|%t��d���0���bI���7VVw�����J�7�����v|���v88�R9�Uz�-+8����O"|��غ��	�?�Q������E������ >��N־���K��˼7��w��^g�^����*�A���E�Q>�	����˗?���*'���?z��x/.���\
�e�S�Ix��NP+y���{�CR�-cz���(�^!����pm�T���W9�9��r�V��9V+�q�ςG�bp@ƚ��oA_0�����P-ڗ!@aY�j�we]ҬhQ�����'�p�1���zS`C�݊�T.`jw7���.����J戼��l���D����d;�f[���@���E3K�KA�;��L ff��`���a�׾o�@¯J�QG�]FءMc;�+���G�N�26�v�BNJ��H�zu6֒��������;k�km�
�+!o
n��"��J[��5��%�p��@+�{��(&i �����v9.hq��!��r^T"}K����Y|W�֯�WR	� �Fu�I�3�=:�)�7b��T�Z?�p<�>��~��(P����"�^��s��B�-~<���qdۍ(�iL N��ӻ��^�'�'�����v �M�R�ѽ��3>tS,F���YK��@f��=�P@��4& �]�je	#]AY�a�琒V��Gf����������I5�4#�u��׸!�vq�'��5���U$q+`̕�|Yr�oo�N���I+�N���w�����4�$:N�q\Uc���J{Ԯ��l���B"U�ibw���^O��X��bxw�.��ϡ���>ݙ�:��dkYCu�ǀ�{c�c��,�O���-��/������i0�'�l���zx���Ļ.Ѯ�i����bU��#�H�oXd�)dtn�pY��9TT�n���2 ��s��L�;L�5 Q9e}�Ų/U�{�j�g���$��F�����[Dv����?���	fDqv/�I�y�"�I��`�����qw�\cj��
�f��g��� Af��؁
͟���%J��L\�O��Բ���70���2w�pI4f���wr��y�\@��3Dٲ��Q�A�UC�\O����_ͣ�Iw����	Iq�Q�2:���#6�^�-b=�u���↧��槏Q @�DS�W�����.���?�mp�$;��o�/0?NN��Q}�"�bߪ򺮈�sG�u��'d���x�)�yu�@:��Ȗ��+����wZ��|k��u��H�PNʆ����+�߼�"h�zŷ;�Y#��V6.侈�E����u�ή�F�Z�����Q�q��߂&	'S*�𦻪|3P�`'�C�����1̯�r`�샫���8�>=��']j7u�^4{�����G�7������fz�tl��؊�B֘�'~$,(OG���M�!��x��V$h�u$�d=�֬9�x�U����&d&�9�W�uT% K�J^�l�V����O�h�S�W��#������\��7;����b,��=H���FK��������ފ��JL����kӉ8�v�d��9ME��6Й�"�I�`����(58}2}��:��H�6�wJ��׆!�<�d%}��MDK���O�0�4�Յ�Q�9H��|d������7l�o辳Bb��u�L��	�B�l�^v ����9�"���7�}Z{f���q
(��x]���[���t�f���X����.�xά���ҹ~rJ�>�AƆ_�2gxd �>�j����,�^�\Ɩ�Nأ"+�@<h���}.Fޤ��o��\G�z����Tf�ʺJ��̕d.��T��h劊[�D��4�c#�����>}��%��ѓ� �4X�jl��Ah���[b��熛����:&:���cuw��:�̷``�����#�;�]?!����_��"��ؗR]��.T	���;:�y��Ġ�����7e���-p�W.�����-X�􌡫Oe�R/�z���U������`�����Bj�_�d���{�!����q�~�<D�yV���.�4�M��ǔ�3:���]�{qI8n��� �"#/6���2�8����A�h'�����H-i,���#��o�\��o�.��Sk�P�-w�g ��a�>m_N���Z��x�q� D?����`$of5�G��mKY�Šw�Hlo�Q�[���g
~8c2�
5{]k��y
&X��~�%:4%P������x�<��3t���q�D�d�C�^�q�SJ�+�5~�O��F.'�/6$�������4���M����(⌟��wX{��G9��[��g�O�G��L3u� e�p)EҚ������d`#-�n�Ji����d���T�K话;�u�嗌.j�fo4t}DYcA�JWO"��cNX�W��۷A�W�sـ��8����y#��+���	0�����S�hx��V��*5�&P]_�����6�A"E�����t&!R܃���"�قz�)�����{AD؎]Z �yL0�AAL�Ǫ�o� �T �vޘ ��G2?]�T��aF�L$���i��X}ݩS�A=��[ງ�P��&[��_!&��������Ҥq��h���BG�fm;�0!�(��8����_��,�*'���+L�|XEpd$(|�"va�+�2"{������A���Ks����e'�2�="1��p�C��&�G��c�>�F,|Q� �N���P;ў�.D��y���D �7kS��{2�/&l��0��Ќ/�Q[�%���<8+���E����r5���񅦊�U�)��!UQz!��&���q�I�s�2����hb�(+���y��.*��ݼ�[����!R[�Ä=`�Fx*�ϓ6�y�9X{��"5(<�AZo����$��I1A��F0w[w�p+����m=��T%x��qtlf/�(��*dU���i�?�f�=r�:J�w�/�彅U�4��8�#TZ� #��= M$�3<�ޯ�.s��3��C�j��b{8�Rl�j
�Tq��蚙�O����G��Hu�>�G6�����6͵�v���v��2����	���i�Tں6�v�d�S(`"Ra��.k�R/n�T��6	/�p'!��9]4���K�H��_��p���\�|`��aOh��P����w�Ʈ�o�W��Ҝ!b�E'�L�% ��-�7�_�1Jj��/@����2;�`����Z׿(&�r�!�0���Fk]�W@���M�揀:I�c�����;��1�k)���A��%���g6��/�	b���\E�~�Z�)�mVCw����W�^�.�qFya8�2�ۙ�lm�$:�%�oiX�*�E@�����#yǰ��G���1�ɰy0��!߶j��9�}�#�#�Ð�4r�jak��/E�� �h��͒� ����UI����m�Pa��U_��T��T�I�>��f{.gm�iHMjɯ �t�'z��ǉV�]�4�#���ۑ ��jӪ���W��e$���N�@�R�l��6=�*g�7����Y�*A�x��RܑUj��8�ʭ����1�1H_� BU��D��CH��~���:�<���|MM��$zb��X֎L|��F7O0��b �^K��l�=Hf�R.v_n��y�roL&�B�f�By��Ǎq_���h�:CQD�m��,�[?���n邤C��O��� z#��ӯ��V��R����(Đ�a���(8�͙y�[���i~ݠ�n���UҊ0��vā�R�9�(/ݯ�1�q��|������1̘�^�v0���:Ci3[��}�c���J�E�A~�����ʣiM]��џ�qԁP,a+�I���'ڎ��t�:v������ �.�=t��n���=	1	�~浴嫹�'?{���I�����H���,)���|[���ik�߉��	O����WilY_��\DR}�'�m�D;i��7S���脌��9���P)��w���\����.�'���A�p���L`����,�� 2=���e�\��z�Nژ,�s#�q�P�Z=���	��s�cN�,'=�L�!WO33�;~nr�GZGO���}�]�a�Ω�2�w|QͶ<Y�F7Bs��#�|O�N�_���pX֙נ���چ�&/X�2��"EM@�v� 3��*��L�E�^�b��AS��jz��бL:�Jx�
_	�`�}���`�<Y��W�]�d{�Ҡ
���ؠ&�RS��մT@1к�F��Mw[D��2��y��N�(-��$��d�{����G�ս�9�Kr�ߧ?��!^_�4�iл�.��.8�`0]���ʂ(
�Kݫ��_����ٟ=�d;�Lgs���a����@�9��z�����dPH
�\��6� ?�%��o!�����'�8��$��ҰPI�>���aXJ"�G��-�מӭ �m ����xqX%9��pb��&'Ppux����	�^��{� �qC�xXǬ��&���Cû	K���
g��y�}�%�pxJ)��tDg��#r�*9�1D*;!�D��.�!����$y�㝜�d������q^s��������J��w�WM$A��d�ɯ	���I�O��M�����T�ݵBP��{c��3G�����-WxVV�g���$��z�C@���z�Ak� ҋ�	����iT(5+^�$�	�Ü�5���G�<O�Z�B�#�X��IV*�,eF>���L�ه�bW.�!,{G��;V{��;af=�����V���]t�o>LF��xJނ�4l޸9W��}x�0��g��\�.^����	܉��5ʚ��g�����7���;���]eGI�ުp*?�n��(T���6�:�DEߥ�V�]��d�}�3v��C�Sӝ�Qu��OA� ���@ ڧ�WO5x����Av�Q�]��'�͑.lЩrկ-�A���mj�2��̫Վ�A�B�#|�n3�6�dk2��E��.�eU���2�Ĵ
D�d1�@�X4��D���N�h�yYۍ���B7�G�/Ճ���r�<nA��ǅ�`��U��M�-���ޭ��E�^@�͏��-(Ek�������۟%��܎�|�ǨX
G(qh4���5��u{���qyw2f����>���P`�9ܓy63��%C��㓒�`+ix��`�ʡX�U���*����bW��1���g�A �Q����E,�Z��~�=��j��s�5�R�;%�`� F���r��P[��V�����C�k�^��Z.l�*۸�}cJ�Bvx�����9����Wn[�o'� �>��,	f������,��6�z0c�����%)�Ǣ���:���b+����VԻ��5��ђ�Q/�.�����ج|D���a�I�#Ѯ	5n�&y8�$UI�QE/2����m��(��r����,k� �s�<����Q�躿1�Z�@�T�kX�ƐƑ\�l�G�)�
A"���/OX�6zϢ�Uw	��ch��Bo��ME
�G�X?�-�D�ҏ�0{Q�Oy4���ۗ�vَ[��Nm��&�TTXC�O�2ƫb�#�4gL�b湯,7|��ޝ��!�
xa;G[���4��Q��8��h��e��˂�>%2�c�	S刢w!r�.��{���
n����d���9�ir�"+bH�K��\�y�4onL6#��I�a�^��qdi�]�6F{�Ϩ����"|�S1���������Rg�#���W��+�%��BwMp�����Wt�}V4��V�I��e���U���SW
�w战5�p�Zx>}]�߿_�<Ƨ5�N�%��������D�7�c��3��e�Pa���z�gh$=��n��$��, �.l��=G����G�,�=�$��ݗ�A�{B�c
�r�<	���Û��"(NZB��J�Up(m�����-��
ˆ'��G�7��X���m2�e�@0�v��_[�	*.��~v��	����T��EV-j�=��$!� �����~�Ϝ$���#s\����N�~�R�~$z��]wY)�ä�B�����N��uk�_���,H� f���3!-`hm���٬���k��z�;��6�-��pd��8�Q$ޕ2���j��m��Je���h�L�s5X���ʅʇ����D/L��A����YXb�
�,�p�D������j�=��������i�p����B��@����8���~/���f��	H�[��hT�gr�y6�>a���,"��z�(ĿT�,�+.�)�͟��fR@���7	ϯ�ȼ>>ZM�ĿE~��t��(	��/M0���r�~^{���~�;���,��i ^pk@}xr���|�sݫ�����Ѹ���)����71��4�4{�OZ#3�A���0ץ\���n~O���\!���<k��՚��➸s%����zs,IU�d􉬂x=1_ �s�\��b 7�~�$х�r��+Ǽ�9�](��9�p�p�H5��r.�7 �|�SQ����(��P�-���k��ۦ0�p5e�4a}�F~�y=�E}���k�#�a6tw�v"An�kx�W�s;ae���`�