��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������T&|+��J�ʄ��*a������A[tFI�2�ZJ��#��!٧��1�H�n6�4�0�>�NS�	���C��H����[���qE�<���oRn�*�sF�6\=�-����0�ɠ��m	;�΁K9GN���Ho-}�Bwɷq),&|�?�����D�ī��&ԛ?�&#���\`�(��R���q�zg8'k���>�LY�V!�Fߔ]��=ɀ��]�O���k����N)[r����ʡtө>�z����;���V�4C����,s��>Avi-(kV�=�\%��Mq�N(~���eX�nϡX��6�oq"1�Z��2��O�%woj�Zd�|��W�N뉡��H�"J�i!LFlÞ����g��d)�-��g�`�!;y�nG皇�}�nIEⰵ������<0L��L���|Ƞ�et?���6���)��ڮ�j�Rk�J��,�50��YV0�&t�f9Ou���F� !�Ǝ!Z�����q�@�!��>*�1>�7�5�5MN��_6����h��䰰���D��Ns���(�)�Hjh.� ��Ii��s2IY\����	�(�9��$��1��+e-(p��s0zN�XqH!��L��f+��em����M]���%`o݃X�{�i���jM�>�O�T�g���գ�i��s �ʵȟB�=�zGb��N(�
����dn����m)�b=���9'�C�s|�
���U�Ǧ��n�.KېV������w���Obt�x���!��\���D��k�z]2�L�KI�fY��6��_'�� �Ge	�B6�JO�q,��!��w��e�C$��+�w]���$�!Բt<rៅrA�_�[LU����L���vO��~�$O�:@��7.�A��buѬV�'I�g@ ��Xt�>J��cYz�\J��'�'w���`�������3ŐCX�|e�p9�F3s�"-z1�b����k��-���_���|�/�GH/U���'I�e��8�Chأ����s?�(�� D�K6ӛ�p�����xN�Qc�~�m�)��Aa���{u�dt â�R��x�8'��� ě��يVQ��O�� x�v��8-6"�M�s��E�N���P��b��H�����|�v�u�e�o�u�Ɗd�dX���3{��-V�N�J��4t���G�'���2ʎa��W�B��7�T�O��gxmX	y�c�)�ٙ��&�,�%`�� (T_$05�&�i�����d���68��ߪ����1��׋�r�L��޷sva����
�QR�����D6�5#��\M��m�i��U�a������ϣc�}<�p�:�:�]��G)n�4��k���y����� ����ﰳ��m+��?��$B,�[�=�|ie�0��i������6_�ja�̆A��ee�|�0�����m��B��l#�w���R5�y�;�g��q��Q��Z����ܒm��5.�g��!����wc�?�($=zB��>������!A�3��aQ��K�f�6~c����Eih�B��p��ZJ�e���i/^P�ҡ�I���jy���U>smj�꼎)��ޝHŨ�=���a�azr��t'+V�:�<4���{G�rjI�-�R57�*��'.8)�Ȧ'<D+ ��T^Z&�H���l/�Q
=ar���9���r�:�HO���W�ύ�GFim����l
�#~ʔ��;���g���CS��%�Dpd�7M6;���&x��u ��#��v��23ʋĶ��Z�d؃}��8���D(�0�䙇,s��ӄe�4%�ØG���Bo`'Z:���Ѕ�m2�%�)]ӸE�Mـ���"������Pb�tg�K|[z.1�ڦI�|9�~�3�����)���~ǘ%��F|'V~�C[	��P��؋3���C���w=����O�Dr��Z9�����/��a����4ʺ���Z���s@��G�btX�A�܀ޑ.�u����ʰ�0���(.����7�Џ��F�PQ����6�7�~��Yn1��&��M�7���38�#	�>����{�EP�Y���ۤ����V9��ñ�z�P���4�9~�Ԡ�����)��`~�ͳ��n�����>>s�	p�~�N��L�u���%Iú��`E��> �%�P��m����u��ZA��$a��I�?6ʌ�jr��I�M���G�X�8"��v"�����	����d��IT�����Ab�|~�x2�bz��!�]kj���7Ĵ+�)��M���?0-��Y�̪ux������$�@SZ�G8E9��/��!�S@�E�J`�<<����S�.�H�T�s���7���;�^��A宮7����;�b�R�t����\O ^1Ϡ����Q�O|���L �Ə���S}�h���Aj�+M����v�韂a
P;���^Is�k�t����dP=��+�b��Q��I�5 E<<��c(ֻݣߢ�y_wD� r~�xV��ۛn���+k�D�b���h��+�Α�� ȋ�o��ъ4���"V������Sj3�Bl���^��s(v�L֠�P�;~Y��U� J=�Z_i^2�.b�g���� ���!(fvH(��p+�/#��4v�j^Q�l�ʣ�W�rG�f�pJGZSi��ſGt�oh��f|�j���'�����d	�%��6�ڰ�ĸ�,�'���5ߞE�9sd�D=��ۓк�m{u�&�R�U��b���ӱS�+L3ީ�vBH?UJ���Bh1��䯎Jq<�T�s���!�P�"��)��1�:��s���e0��'�V2XY��	�kc���X��;�E�=��xW��,j��	mW�V@�����y��E����YLK͙�XHT���0.���}��H��#m�B�:�Ε*u	�b�;yv��zj�FxfN2�oZ1��s@Ӿ��)�E����%�L�_n�g�T{�{��$�.�y3���q���8f>�A��&F�m�������vj�J�j1�a� �.Η��K:_���}��P�N1���Ǉ���f��c#�m�7�K4Z��Q
S�5�N�c	��R�<� ���A���
D|D��tF)��KGƢ�Q�nn��oye(���
a��!�(� �#�zK�(x2��%&#)�w
Teye�g�`h_�������J����8��붞�p ��5Em82Dl�9��_|<Gjgk��I�y�t�����"��9�W�}�xZ@�exY�.��ܭ�7���>V��n׋�"�lw�o'-�A�D�W�&Lؓ]U�̠sL���p��_Y�V��33��~Ɉ��(6��Y�:�}�J�F7��t�ie&P�\�o��0����po�HF�%��=����>����e�Z�*R���`�c��r@��>�6�Ѝfg`CGj�8������w��N�\�+C���U����I��I��T�f�Zr�E��-��-0[�(\�>���C�g�@�7�'ߥF'JO�!`��)(Gcr����N��]����T �E�	Z��������`�J8Z<MH���Wc��u1:�~��Ӵ�!~hIjz3���s^A�Y=7��q0����c�(Ͳ|�~H��8��g���<l���vJ(&��� �N ��ȿv��\r�����ۿ�: 6癝���i��e=/��ӷ�蘀���CC�ަT��g��t�T�B�P#���+��� ꈝ��[���nn�]:$�:<Jݕ��'ZF��X"�Ret���&�z�o��3~��N�Ȅ��#�j�6�qKO�PzU��5hkb�����	�y#\go��3'�DE�<68Y1�f��)�(�l<Q��ޱ���ai���b�(X��?i����܊�(u�u.�B�ͺ����F���1�YK�5��I3�[�7|L/W�G�3h�i��*_qJʜ6�f�����Ol��>�D�����$&��Z�H��X��>�J�4*l47��׻C�ql�>φ�`����՟C��Dv�*�#��&r��^$��4�&�g�}��YԼ��U]��h~F}`U��	���a¾�@ַi�M�*g*�]�H����T��b�>7�}o���bn���W%�>�"��l�0*t{�ҧ!�V.���!9�sb����K�����.�ؓh~�`��m.�dL��E�@��*���p�C�]�5�l^mz���ðC_�3&:�e2yҜ�*-(�8p>��5Ieh.t/<�w��ꕒ&89v:VP��#1��t�㢭D��oo5��@M��J�*�@f\��~k:N��%���ב�9Ƹ�*�ac�X�:�.�}�\+�`�^�U����M\�V�>��Fyci/*���;B�[H
 	��P�;d��[�{�F���:��"� �Kd�U�|�����'��jN����i!Ë��vv���Z�YyJ���c��O1��J�[-L�#-���ӓ� FR<d��#E/S��I#X�妫� ��L�ڣ�ډA���olCD@�Dp��#mB{#t!�0���oR��3E��k�u�`h�'w�j�n
ޏtc�X�Z�fu� 2ab�b��0'��}ªج��FsqW��Z��@�^������wYl�2�<4���i�D{�J�P޹�"/������R���x�TI�L�r~�����08��"�l�k�"�ڭ$s�Gt�|J�e��E����������՛�ϩ��L7�3T�Q��)i+��p ׆�q�W6�UҴ����F�>Z������8��Z3Si`ǻe��_J@���Mu���dؤȍ&������F���ɵT7��� �:Syԗ��%�y�mY�rHX�"։��&M^Ey�'�?���fP(� 8��u���(�x�'��Rܮ��׎����2o��~+ax���*�������7n�e!��Q����J�_���U܍_�=\��*�?+]��r�A 1`�����1�d �Z�ޣ�J�P�֡������jc�2L1�����R���L��}7����My����]x!�2�6l�W� 3�����\`uKd�~~s�qd�,�^����Y@�>k~(z���X�_|}Ն����_�8���to�.�\�o3'6vH������̵0���s�3��|���'�Y�jdla��ڴX�H�����>���\�ݲ�r��s{A(7a�i���TX:@��F���[�`ߡ^F1���涣�x�9�K����s�O[�E���.|����<*�w���6�zZ��ce���1�ZO]�1>v��K_g��H5 �t2&�8�	ɇ3e�{��S�2���J�&�]aB��C�2t&�9�L8�\�M(7���[O�֯�[\��~��V}8���V"�WtH$d =.����Nm&��c��/oĶ.�_�q_�W`�'��K����sж�mE�dp�L��͓����~��\�����H��	�c!��=��sJN���y�s����7s���#	ҟ@~*w��C����7e��+kV�,�|���;.�'�zc �������oHj�)̡P�3y׋ה����mڠ���I8 �/�-W�97�:����t��c?��m�}kj7E,V��wl���5�%<��f�~�H9��+7О�ɟ�j��«�vEQ�.���TS<S�o�=�����;+#E��Y���J�ć�h1a�.|Vr�����a�e��u֮�c�G?db���c3�Og��V��S���LU�E��Н����iC8;��);��Z��u�����E����`���R��&�LSxw8�\�7pI��aɎ;9�"A��Ԣ�K�l�p�<�*d�o�"�
!YI]2w�j�NI��9����nB����=y;@\�Y.4�mḣ�e�B�u��ވz%(u�oh��T����X�����|���I2��A�--?\}K}�ˮSh�<���@�oh�&���0Q�J�Q<�(.�ǁ��y4�}�&Ι0zHA䑖��U�H2H�N����wp��b`�9=�����j��eWn�{�*%���'�s���a���o�?��T����¿�8ĥ���I6��n�=������Q���1Jn�R�]4��u4#����]L{W�ũӶ}`b{53����	��\��$̹4��V��me��*%��{p��\�5����h���MSz�����h�N^�b�fӦ ����8�i�
d_�R���P�l��%����Cn�[Rr�"�U�I5���_58�`'�oj���aZo�:��lStQ��pm|m�����̰s�a���6�n��~0��Y<��*{0,}k5�����|4�^��M������OgAN���~zY�R��✜'�V�AЧ��"���]�/�3}b�&�+7�Z�7�(���B�̓JҬ*�
�̾Zr���,�RN�.�;����}��赶�γ#m%��glQ:�e%C����� �`�M���K���`��$�ʛ���c����8OOD]�j���$<�#��|uz����ç���"h��;o	=JC����d�l���1����Ȟ��c�U�ִ�Ú��Tx j��w�N�Q�$�i�-��<##�SsQ��!Ce�!VͲ�j��i=vZ�a������dy��|K˫�0'<���+%��J�4�Xf����t��-��*1M���7J����։A1�躬A0��\~��7`�4�|1rH� ;}�r,��(x��U����ugy@�!�[?
陕�Ͱw����"
���\!
�\�e���bn�1�y�Y{����OG��C�����e�n���V�Ǭ]-\�4����爔B!��}���ٟ/ֿ
/G�����Sx�P�b��@#)4W����",�<@��-���#}�I�*|��� �\��)�I �\��9z��RI�i�3�#ʢ��p�yP�w%H��Xj�`j�$�5��3l�V��'�Fɹd/u� ���o+��Z����_�J�ϲ?�*R��M���aɀ���\��F����EM0�ZE��3��:�@���mtVAl ����f7|+
5�Q�F�LuT�;��a1�FG��1�z	U���nX}-����wT �\����m�ݪת���o��pK��9�d�h$l�cИ��D���_ `W�W��hV�ٳ��͵��Q��%��v#7'r�w����J��.���.E�,��m���'��(�}*�Fm0%˚��w�����K<D��˶�1�{ޗ��7�A��G~�������=5�K��:`����U;!��5�s�T�?�=O`�U7ㅞ4V�����mk��3Y���8�~�$bS[���ފ��htr")G�ϴX���5vx~ȡ��c[^�I�A�æ���<�q?���`ߢ=z�M}�a�k���"���JUE�Ʌ]��V�"F�v����U���r����h��H�=��<:���FC=��=��NB�O��4�eKP��_���;��^h��gYl�ʣ�t6`=���Np�z������t��4]��?C��x�$�S� *C4��8�ߓ���/�ş�ڽ�W:�O&`��4GŘ|��0(kw��NdG{�y]�����fNDO7��K�w�+�{a�w��^;����s�L�^|<o�Γ?��3�˩tQ�6��(Z��� r�Pc>��o����{�F�>���^B��)�����F����K|Ye���He�5c�Lo"�0ʳI�q��6ޏ�Z�����L죭�8����vY\O����塳0�����*l�?��Ȍ��MI�e�W�RrZǔՄQ�6Ø\]
u�Z�������%�K2<�&�d?��[W<7	���a��K+o���ϻ��F=i��Q��4��=1i꾭�&ꘐ����Xq����Ѯ���r�0�1���LT�W �O��ca�8�ٗ�	����X4���m��x�F��G*pn|��m�.1#XS�<��j�`0F��i�c�[?f���.I��v�[�}�nNc��}�	d��R�ȱq�U1�"�
�_)+d�y`]m�ƻ���(�[�tR_ڈ���ꓻ�r3�en��3����^Z�Z�j����hХ��RrA"��i��9d�]V]P�v]�*�{��������b�X�n+������?�1s@$��#�ɷ]Dsc������~^��!2�벽~���4��̕��\A%߯�=g7bO.664���{/X`���t��f v�6�+�x#dB9'5�QHؓWApQS�헙�l� ���RX���Y�Zf/R(fza�����y��n-�$./d�O��=��;�Ë]�)����P���M/v�ɓ;`aM�G\��Np>�����)��1�X��)���=~�;�c"-� H��d[<���D�(�2�Ȯ��D�E{�ᢘD�d�����de?I7v�]<^|uL���ɚ% d=N@��-+��ch���Ď���p���|Yw/�LC)���,<��L��r�8q��>'$O��H�[F��C])s3>''9��֦�x�5���HR�Xb�K �8���#f� =|摮��<V��D�O�p���f3��"����*�.ט��8��L��2����9��:.E��0>��H��C�UKj�|�<�ӈE���~U	؎uU-�L��,����������qÜn>��m��	�3���ݕ>Պ�:Y�~Kҙ��ciF�#?�E}��{�I;��ɾf���_F�
q�P��tV�1�s�o��w�qɔq��}m��r����rg5\���(�k������Z��j�^ܵ~��{�_������K<�>��T�S��&�]���� �丿y����N!_�ļΊ�t��O�������:��E�L�[ ��܌bmi��b������cd��2�X���$�F���y!��I��U{�!U�p�쀗�J�в�9%�X��+�s���1��%�u��Q���2X��� ���� ���5����m%(l���*#M���<�)�g�P��j6��v�Fo�t}�i0�#ؤIot8Fq*���U����P	����(�_w���F��	�}#լHwJ��D*�^��P0|0�ݭ���+h�I[6�Z�G���$M�!M���>�I���#X��­��, �Qt�S�?;�^�h���T�
�&S���8jMc�*��aL=�e�Ԕ�!��$��i�K��g9#� ���̙��=����0o��v>/����/�R!�O ������_J2�;qG�{G`x��	���K?�nǡ1�z��#\~����"egu��V]i��e�7Je�t0�o��0�S^�A�9Hhhj���Cw	e(�<�ϙ�|@��
�!6�8�7����]N��C)�-y�r�BF�MB�r��pUtl���O3�Mr;�ok�u�^�/>��S8G0eCR(;�H����`\�gH�!��}��|�v<��~<�8���3�	�ס��N�:�@
�h`���E��o�N�0��=W�#2O��SSh�q� �v��:h�ݣ��袈��^�25<��X����Y+�e�k�A�n� =�����ŲzG�+��|������m L׀H���]�]�%XO���[{"�@z�-<�c�AΝ��W��{��^�k�D�B,�Jӝ�2y���=�|3J�A��� �����<*$t�5�V�Ք��g
�л׮��aR*!�/�sg*g�BxǛ�7�VF�@#��{\[s7It��m�z���%`Rcʖ���R0#��ܞ����rqq��Y���5�yH��~iS�@0WV��v3M� +4���pœ�U�,ba8-eH�Gi�^����3�p-EU�`R^%h'��������q�
�1��y������) � Hq��/<�����NR�u�H�܆#��MH*'��%��3�0�j]�o�H�����O�Dp������	��V��X�������\����#��m�QF�ӮEl�i-�C���y2s�G���Zc��<����)�� ��F��"Ώw\�1D=�]d1�5���:)==ˤ�X�|9e�L�m�}HYb�Q2�o:oѽV���:�h*�bN{x�Z/�,��U�	�&>q��rFR"�"1V���aӐBHB��j�z�uPI�`Qj�|WA5� V2dRI���,�"Wy���
���s�N^�Mr�u��6��m��5�t4��q�4��A_�[A;��D��g�]��R���o��|�a��#/�	��s��-�[/%��4D�����#���W_�;$|��9Y�ā��΃�9b�	�X\-����3���)}���Q�h�x�i��X�@��"�H�1�3�!��ռ�����ՎKIEk÷��Ȩzꥪ�o(���Z�����ƪ=�֬p�@~T�����mm���)��%K-k�$�:S��Є#:��<S�vݠC�B*<�6TOWa��X�*a�f�\)��٦9��4UR�\Z1��=	�d����%!i�����x�(������:M�I��<!N�0�Oc[V�Ɠ��C���/�1J����>��1���N����L���)g�;�h�Ȯ�~�A�Q��I���Oia�6l�%�5�Tr�e�L�Ǒ�[��R��y 'V�l�I��R��Mr����y�L��+�urΛ��g_B^��Unϻ%Բ�?� Ec��'_B�ry�4�� �ݣd`ܩr�|iFrd��#шQMrz��}gW��\4v�a��)cK���w��V+��s�L�	NM��rN���iB���P��sm`�(M��?A�o�A��.��vOgJ�;\֗`T�
�F5T�W��"�P^��!��
Mv��)d��g�ֹ\�hj5wO��rU��w/�K8&	'�/e�n�I`=1#Mi'����1��."�aV"Mª����N���s��1WvfHͼm����8=� ����8l���R��é�z7�0��F7Ŵg��V�s���2KXD'�7��F=e�n}���K���х_]��S��� (E%Dc� e��h�3���\����ٲ0��[���#.<U�Z�:|1�L �Ӹ�U�Zg�Yo��w��B�?��d?��
���c��L��YK7{Lj *.7����P��϶�h�ܠ�ʌ��Sk����Qn_�f�����M��o��b�S
jh��&���{����k�
_�<[#�!��\�*Ng�J]z4��to��nF+Q�R#5{���k�"�t]�n������Ō�.2�׈��t3���d��;RTY������Zm�U���M>���i��YV4R@�ϣ:�x*E&�6���޻������F2Qi�w!���%�\A�`t���r����{x�k�־�<@(|&�=^�d�5�3�;`⒊��T{F-׺>��xI�$Isg槙��Y��Y��B@R`��`�j'�����y ���Z5q�~K�	���d2-0L�h?Q��BD�����r!hbu��G��X{���1��$[�0����:v��Hc�>��w1ݥ��2��g󠁳������O�K� �����>�ŲS�^}Iu��Y����h��# ��Ob�+K�w�Ehvn���E&�:�T���Mߠ���%=�Ys�C,�L��s9dG���h��l=��6�'-�.�fc]U�:X.��׈P�����E%?ӄ�?�$�Z�\�UY7�+����u�� �o"Nև�p�������S0���`໹�c�����C ���r��\��ꐨN`d��~�9���M`]��G�ؾ��}�.>��daE���1����O<�^K`篡�N��s�	,���:4�����˗��l�I�e�R����yl�>�F��1]�\��Y��>�YyM�4N�D9��g��e������ߺ^�7?�=U��]#'0�h���P�w��.�a�X!�	�q9�6(D,���	,��s\
�7�~D_|��8W8"�#k����ek����@G	i���o��@K˪��� U��>ԡ:/q�4R�N|TH��7������
>�S���+p.z�3t��HG�ʋ[�01�*�Fg����? ji}GeiC*�w�d/�u��)`�Z�o�D�\�e�uVf�b@��P;*���EG�%l'�������70~0X��k�J����G��(1S�ĲK�ͮ|��9B����c���>粸��[�B'��v�4�Ȉ/�C���.�c�m�B�X��@��YT�ܢi?̺G�q�zg$����q��'ƽ>�Xet�����9�������/p�����G�K��6:�8��c��}�R!5k3;��UVK������ErA5n��B?������^_���_4ʭ�֬�D�a6�z*-�@�Gw���Vؘ��F��{!����w�4n@�`��L�a�4֎���7��GF\#at�3G%�WI���=�����ܔзW�)F��N�����g�" �a�s��`-�r�曭-�v�����a����8Kr��ݢ�b��0�k��V��(��s���d�����~O*΋��n�9�țF�����:�3n@� ���X��`3�Tg�����T'��	4B�K��~QG��j�sl*�� i�`n8~�Gb���h?�߷��p��z��$�{@U'i�k~x8��jl����%\�8�����58S�}"Bdkwnm�_�8���G)QN��|�EҺ���2�*xo�����M�� �c�v�Q��tgק1($��u�?Pf����Ε��MO�"z����M����v,�0|ݯ�:8���L~��"���z#=��w�C˯6�*ԜVS�D�p8�g��EQ����g+�3�ُ��ă�|�mշ��i���ldt�'�0!���x���-(��G�8m@�	��2ůyQ�bc���: �R��z�I�x-�w-���=���.$�n	A�\�(�t��I�'�2ԽC�4��U)Nݖ�|6�9�~dO�s���C�@�F��Li���_dBf��xՎQ4��K�_">���҆��� ��n�G��k"͑sߺ�nS���[b��t����g���p~�v�Ek�����4�vD\ۼ���r����4�
 ��"q3�f��m}��t|�N&�5�mY���*�Xj�N��2�ߑf�X�P�J�3�u�MF���"�����'��c>���&����>X�z��$�!Q��׽K�D�7Z�3�F�V��p���h��T� u�O(��K`e��l��[<�u��	�;�ы�G�:$�g����.do�&��R��;�2����6@N�XX?��LNR�UWc��H\i n.�!ZW�s��O ��>�/2i�ˀJC	�O@�"�"������R�� p��
9zLW��`5:���1HL��E6
�_sB��g�(��Fkϡg>w�_ɘwI����jڹpD��]�\'��;�6��H�);hs�:��
v�R��K��Ô=L��K=�bAG��B=���S�Ө����]���P���}�v����@��^yaz]:���FG�����=���&�Ȥ���o!�Z��g�3�<RzYs]��|"��1j�ĎQ��vņv.L���e�3^�w\�@L�b$�^_���zqrߨ�r�Y����{lm�XcP*U�W�J0y5C�2���\�vw�K����:��e�>��Z���ٕ+����ත&��ZZy�ڐ�;O猺����[�u�Ov�77C�uI�~3���j�"�*%�
F[r�]�� 6.�9n-��V}��[���2���U8�a��L<ot\\�X�����0�[lL�c�s
�迚bk=�M֒���q,��G�ȇuU_�����q�Of[Ϲ���4���^�����T2��<�/4h�sR�s��9��q�שE����	nF$�n�5R=�&�b�U�W!"��ѿ�'��a�E��{���6�{��%�kMh�k%M6�Q�T<8jn2S�".l�������$�R��c*Q�.���b�@G=+���`�ޛ���Y��.r�3�[{v[���Q~	ڨ�CZ�.��:�X�xԾ�4rB%��{�bR��B<�)ߝX�=6b��f��R�&�m�5�+Z1���)I]�Ef�`i��n�Q1�JZ	ԟ>8�a�ⓁF�>|�x���Bb'��|:�n�oR�Q>T`��c���o�E.q��n 7��U�@j���퍑4�f"Pf�Z� �����i&���1�w4��ѣ�������to�6]�ƅe�R8�$��#����Li��$�M(ԇ��c��ݧ2v�Hn�TM�cŧ��.?0qڴ�f%�ݥz���0�.w|˅�U-K"]�s�1!G�`�Z�0��=�}��y=i�����e.y;A�t�t�k��Բ3�Y��m���yQ�pT�J�J��c��d2§%:�Ibx�{����[7�]w!w씇���f��]0=���޹�5O�9�5s_1�_���&�ʎ��v�A���bNlj)!�?�i�e���qtRs��^[!I#Y�8nA�=q=�ziF�n�L���s|"ȕ���F�'�)�x�;��	�S`@U��-��UД���=#�t���d�ሼ?MH���`@5�x���B�pa��}'˵z��k�Щ旵��u:2��l#�!�H�dAa)�eo�`P�*��M�L��)�����P�=F$�o�Vy�Ȼ�Ds(;gF/dJ���I� 4]g�*i��.�rc�"H�Ҙ�9��7t`������%s<��q�s��dop|�J�Us{�#��J���-E+u-S)&?��@�q������Y��s��+_�R��O!7���)�.@��T�<#��[~|��j�ܖZ%����mv�lt �~v��r�Q�A�	�"u|�7��A�q���$�s�g�tg�)�X�H2�����BBrp�AQ<�'�-��|�[����w�5�q@�Ɔ*��������7��=ع���?c� �Ӧ�_�@���vLkr�>�el���w�x:�l�<�tt���~M��?qW���׽�6������j�X*��V����������˼1ټ�D�K=�٣��r��a Lk�aܟ@;g�m5)�-ҁ ��{�,���zÏ�����`&� ��v|&L�@*�Ũ�A���-�MI]d�"�c6"&O!t�����JdH���y2�7��{â�`��< ��hec $'��
�l��(�R��#h�7�wk'�1f�)P`lk�NucOB�ge|w���@���r�5�	��QL���r4����r��)�=q5"W���#4]�fn��L%랠Qm�_���ѦA��PgH�t@�<��ӗ���H��S��G���'���pd�:��	���oE!��CDZ������	��.L"���^>����@��d��M��G��-C�^�kR��Q�#d��cR:���.�B�$��h1�����?�V���Mc��`((u�Y�����6�Q4ik7�?F&P��e�zA���'ϊT���ą�B�Py�j˺&�Spl)�T�i�Z�1F�v�48/¾��{�혉Gw�1>.4V琶|�]R��<O쏨n��g��`���{���l��:UyP�
h	~�~�>���y�X,��8��T���SnR׾m�̉xݹRЧ`�5ǋ��?����F�$��u�dNe�e�H�w ʝ���ρ8�D��X\����'i�
��Q[���@��"��`�B�4ٶJ�D(�Ò<vp_ю&�k���v6�7�D�P���W-�e�P��QS2��F]|I�������v�`O������S���",�I�B�例�t�v������ P��C�7l��t����z��<Hq��]h��$$�K� ����F�ѩ��\�Ƒd��M��7����$���ݡ�a�����eX�(�c7�T��^�v�k���ib9hU�����h){
ga>�U?l8rf��7���P!��𵨜E��|ZG� .���pᡠ�l�E.�K	��k5�M�d��f+��${�*_s��ț�g�/@��JN�/�_���Cx-�"�9r�E4#�d3�������Ӡ^�(W��ޢC��A&����`/���{&u����dv�D 
�tdkOK�O)�S���~SD>G���:H;'��	�Ww�Xݡ�|#?�ie��x��d ��3*3���y�*.�Y!RP,I�/� _�x�T
�~t>�$`��������|�A�QWo'�Vrw�v��W�a�Qҩ��5�	=з�6���O�6�|,)B�SB����f����#nX�b���t��?7��E�n6�[M^l�A%�j8���֮�5�6����Kb5�fr%��b���Ó�oڗv����'	}z�>H�Is׊�|a��붚��3*j�]����,!��%ՠ*�Nc �@����ZY��޶�U=�Î��"����q��u�<�{�#)��[���6�X���1��v<�R*�NU ��]���v��B���uT�ߦ<m?Y�җ�8�y�4L�*�#����H/c�M^�{&�R_x�
��=���&@^�0��`��h��N��Vs���ࡽ�s&%�x濿%@g��{�'���������go�?�B�/_zD���9N@��/G3Ӭ�>s�տ��¾4�u���S,�[����?:�b�d#-���,[M�[��I��=Ζ��Y�%���yc�����aʳʙI@]��a�W��x	M��],:RW���}_���:��ͥ�^��w��^��Z#��^&F���ף�(j��J�!��L�{7���5�E�!�3J��R�fJp3K�f�ϓ�:H{jY���[�=ս�D2�F�K�3��%Ɇbb�����Q��H�6�`�M��v�1t�I%�i�"�mb�	�ؒI���/����Z_"�1��9N2�;�`�ە\��y�e�AN;���JmEb���_��ݖB$
OjJ?P�.n8�r��c=�����ա�L�߷WN{#7��T<����zD���r��Q�����:��\	o�G�t�ٳ��i�ܜw������M:��i���-`�A�t�89\Y����<�#��a������~�|;�n��7���>�i{��f�=\ǎ?a$l�N����Dz7H��}?�'u��y���B��2���_6N�&��bgeZ/����}��:��%��s��ld\6?m��EˬD�~6O7�̔l�΁ɱA���4���#\u�n�`����Š(j���C����7�Ӯ�QT>�0
�;�ݕ�xx;��t�����A|p��~#'���D���#��)žjܷ]�=O���0��0m� ;����1���1c��Qs��n�����9KW����T��߼%�*|�d0�u˗�g76~i�������Ca>�U�V��pa��.l�Q	[3r]<�R=�2v��JO|�U��;���9~7�C�?]C�ݶr|��-�M����)��3i�l�Nb9[�X���;$V*��
n�G�];����nn��/d����:��+� #�_�'�<�)�nf�[]I���6C��ISU���`p���N�b�,G�׈]���l>�����RY0&�zw��1x�Ã��"K�Ѝ�6��7��߁�>�Ic5�:f(Ä~���o�a�n(�u�E���'8��.r�8�'�̺{����Y$�x�$�p9�t,��k�k��i��_U���ʵ�+���G?x�g߆P`6������6���(��k_�Ť��n�:��a��mݣ�V��2�E�9Ns1�����u��ʝd��;��`���DF���+ǈ�IxL? �C��>�|�t�j����Ps�A;�\
�y�!�5f@�႕��-�{XXۯq�f	\�u?.y-�B۴!�h�OedH�ǌ�EQ�j��چr�wpT�Әf�x}2����UO�G7�hd�4uc�R_V��m��,P����4�7�Y��0R��͖�
�~�Z����ȅ�tȈ�<�nN������B�u�����w�l�Q�h�{G�ب��(�mT���?S�y�3�V��J~8N�r��(�Ғ�G<nr�Gy���l r�laY�!��YS��2U`�����6�\p���I�H�$d��P�<��(go�9�֫/$����CN.d�����h�c8\�l"��	�)���4�E�t}F��2}p ��:��]�\�(��@��c�-�Y��n~?Q��O�hږ�(N�9A����R�	��Igo�:�訂�4��;��ӹUs�<i$#^1����$l�!��se+u����1B�zѿ�#gcq��	�S31��4�-e�|����7r7�y��)�� 6��������_W�fwy�
��R�@����j����q�c|W�#������;�t��$-D��J�>��>D�G�`?|�^%�Xf��ϸ��9ُ )�p��g��M��Nҁ�V�4�V*�J���J�]�Ȣ���f� �]H������622n8ݺ�šwObNN��X�\�\�n ��B���S�zj����Wt��_�OM^���H�d����T*�Ղ�(���8�߆+�9G�e;�w��wb�F�,�-����p���{�(��C�%�L=����ʴ�����\��⁵��kT.�&������xEp�.
���LQ�R
�2��ծ����D�����R�~(�M���jxk����=ƣ�@���y�dʧX���I��H6x% pwgG}��y$r��m"#%�&���(w��lK
$��p�:�&e�j�=\C�s�R�#���)�_qO�  �U
�h:H�����>T��=JB�<�P	����Gf�q��Ic��uES1����%���8Z�QQ��k�C�JfJu0ľ�h�뫭�l�ή˭�J�&#i�I/��Ѱ��H_�R��mXI޼�H��vgvK�!D�qxs�bg�/#�C%W��q]a��
^ N�NjMȔu5S�r�P��-f��t���z��vw�����h�m!7���PK��k�j>�g-���(`�c���*N/A��k�������gn0,�Y��Q*93�( ��1��*�L�����6���0�[!�t�V�����C���G�4N����X�Ae7���.���I��S%H ~�5�j�����l
�5��"/�CF@��bQ�X�907�kLc�ϳIU�G�{�F,Om,����-~��3R��X��xU�d�E!f؛�o�8lZZ��k�9�G�҃{0����΢!�=)ƩD���*q/Qz�`�,x��ã܇�pB�J6[������{�M�	��h�$X������gR��-���7�O�?��r �մ��6o6�<��$s�'t�>8U<S���;�7�0�|�/}բ�P&�1"��i���0`��U
�@���%4F��P:|*��ۣL�콨BP��8��Ӯ��7��2���G͑��m��ߙ�M�~(��st�?Y����r�	� ���*��)�0�����v����ŚJ�|����6�x�����I@�A�a�}?k��RRr�ƹ�P|��@o'<x��5sֻō�<v�*�(����v�툝vʧb,�	)��͉3��t��]�d8�������
�5���*Y4u!�$�q:W@�?K����PU[7��'Ҙ�y��L��1��ыNV�|.�'�����	8�օ#cb�Z��D �A��E��t�� ���l����%J��1�_s�Fq�����Ǉ<�֓�K�UB�Yj�i�4r{�)֧�:������n��H�6Ah���LJ�@t�E҆��#�b݋��N���Oj�
�,��� 9�=�x���p3#���'�-w0�qT��ȥͳ���A���V��[p��]
�l�NRk�tP*	��2�3`0����ۃ���"�K�?W�?G�HE������;����i����|�3۳㬲�Q�_�Ӡ�?�I\��Wj���`���K�ȽL.(&�R�)"��:�Dbe� I����8Z�K`�&z�~#�1�G)�9�5�(:��� ��lu>1���M�H�9�_1<J$[����<���)�pfG���4��0I��LRH��M��HuaVHe>fۯ�fie��Ŭ��ڽ�.j�g�a�C�"0�����,騎��i1������?7_�stKq"�5��O*8�3��}�=�JGvW,���۔�G��k���v{1��"���a[�S�����C�G��ֶ�d�ֿ��2�j�	!��?�y�Zv��r^*��gn�9�6����]��^����*���"l�[�'L*
l|Z ���`~x~�I�>�yx���_>)j<s�Bc<�:�m�����4o�v�U�F�ib4�u�1�l����9��g����P.쒟l�G����pZ�ڬ�<��T,On���B~b�W�NE!y�`��>l�:|�}����#�<���	t\��:e�.�.oXo���H(V�r�;�3�8<��N���ԢJ3���OL3�`��Lt�W\�͓I?yI����%�Ϳb&�n�g*����8N��v7��8����,�ngo�Z�,���E��a���i#tU�%�+bUO�s,�:���n�S;_��`���Q���ƏƞzN鬽p�����xJ���4 �v�=�oy�Z��HOR��rҧ�/U:N�\5-�m���N���ɔ���jY ��R;<�
4��~$��I:��`��Q����J}�Oe����ƙK\��ֿ�ѐt�[|.�^��������T�j���/�cn7�z�f��)�!���	F�J�M+��ꡅ���d�~Y�y�xy͇ PS^���%S|=R�/:���,-oa���rU�l�ma�����$P%�!QR鱫Nus�VDn���ÓG�l3�F���E����S�3�cJ�@f���M�7�ƴJ�mq���J_���C��ۅ�F�6�5�x���s�P���/��_k������"�C�xiz쁗�ю)�m�h��7�+���b��j'����%�%^��:c��{2}�&�~V���m��T^v:5�H�}�`6�5a_��v�����;m
a�v0�_?s��B�<r�gg��?i3���u��B�6ӹV$\�
�c��ԐQ���6�*[w���a������!��4b|��G& ջS�wSc��E@��0ȑaw(]�y��@�$���ޅԺ-�MȍrKX�����Abl�D���$�*��]��0}���n�e_8/!�g����-k�rV)�Â\.��AXhX^I��ߒ�+���E��N��P�����7���M���7l^��S�_�0Ù0d� ��L���ުmJ�����l�h`�=
}<���@�����PA[q��
fr?͕8�b[N����\�1�0�Ҝs�ChtA7��l����J����W���h�T&]
@� ���aa;��:�q���^v4w|��*�gH%�[���j�� ,+GU���?z�N���1#��<N�1�ʲ�1%���"p|�۰0��H�L�,�]��IC+�n{Zb�B��JlS�9�q=�{�Ep̩�{V��؜vg7�L���_���s'�1���aP��:2��.Ž�5́��˴l��'q`Ѱ���<�G��2��&���.[�j�4��Fc��Hh�a�R\�j���µexj�еDg��k{��p�.��1XX<�<��ʖQ/�9��QZ���V�3�h ����Wd��.��������6��.�t��}C�]�;l�[�a���<��hu�"њ�g)�
�*��E�f�nx�Z����t�l|��ǆ.��͂8�z8U��kZ\��L���MIP �2jqWm:, ��s�`RO��rbvW����q���'a��YP	�D����XБz��x�_\�j�Ÿجh�_��C�Eƞ]���#�{���|�oM40@*1r�����w0��b�֟�#��uaPmF��n�K�L.�y�I �4�1�<�4B�~9N��g3� ���n��=p&���0������7Ԕ{t��p�VQ^Aܓ��h�S\m�3�P���:{�kqZ�>�f�r|�"=�a1����Rr�A�Z�S��l6n��ɒ�,5Y�~��ʎ�r(�Sam��8�}.j3�����\�gە�E�%�ݣh�O���d���x/���ݒ?�TT��ic<v礭��$��4�#7,�Zڨ2�/�i>UН�����M�T��/�y?�,���G��:�W�D�N��)Q������_��R��f+�:�+�r�Bm̋e,��6���5+1	�'.Ź�z2`DV�9)�5917�� ��n�p��-�K��̴��3G����	n�Й��ȹd���_S�}=6�Y�7&��W�&s������p���v��?&d,�no��!�~E��Q���m���.D��ݿs��dӤId��2/A��������0vfֵ�g��9SX�A�W���M�_�������O�;),fw��Q�,���zMO��'�����"��\t�@�WP�JQ@��F���P��J��iת}���E�ԍ@��L�)���m�RCٽD��T���r�	iao��7_�
��yBխ�B�j�5����'�7��c�d�(������Ĝ��y]����E�"�q�-h�Y}�/Xa>�
��̂*����^�>0�tb*�h��فAVj8�������5yG�����Qz88A.� ��	����� �!��l�(�Y��
a�y�z�?\��\	���@��1�k����|�E�ytW��]�������:��S�0�OI�`7�$p�[��K��f���'؜�0�(�VOx�.�N��aD��0����d��� �a���2�iO�b�<_�zs�;:�,}\3ٚ�S�v7 ���!6"�L��ͯ�N^j`�J��&���V��&�sި%�V���%� {cJP�R)�p�m��m��@<��h�K�0sSm�:��*�7W
CcW�r�E��q��� 8�nPiW:>=�P7e|��
10��y�`��Q�+�^�wN�ݞ��+wxtx�O���1��Y�i*H�S� ��1��a�6��9P*�K
E�c��CU�S��@[���ÙV���7r���}-�e�OVd_�ȴ�HU󌾁��*K��]�m�X��s�)�E�����~��n$<6����f����_nl����v$�n'�.�;s�a��z�O�b*���C��)Vo 5+�c��ktlN�&I>ɹ���t�@(8hHВ*p��x���`�e6���,����ǖA�YB��Lx�œ>ΦO�u?jP��,L-��f��p�ix�����g�Í;��t�5�c��`Rs4<T}\G�<.��+I*�:<Ί��5:���m.���É_`���*��;~y%���M��4|{r�
h�+'��+����� (e"O'�|c w��'�溲�ࣨ�D�$�D;�� ` P�È���M�D���k�Rtӎ�rU��k�u]���1"�Z��/���pT�h��4*�T�0��up�1�^�n�T=}��,'l"������W�ncA#�Lf����S��Sˢ���Q�!y�` \@����콋�CH��8�FVK$��&�	74|U��>v�/�Ta
�6�����ݒ���$��g���b��u%�CjW���r9C��-���s�
/�o���؀Z����,�o<8��遱�f�Qo��0m7fz�*�͋�	َwĮv
����}�isO�:b27��d�q�4����.ئh��3���oE�F���K��/<��8,>��/�.��T<��Eh�pZ|OU2-x�x�f�\]�|���	�
d3�#<�迻M\Х�Ockx�-C�ks�����%tʄ�B�������'Vf��q�@�ǫ~��Q�1�{����r}0�Z�ut�7�	g�7������3u<}�n��͑���	#'^�3���y���~�#�TF��bh7�Ӟ�L(����eB�R�D�"���WG�_7;��?��x������e-�����]g(����>�:j�i�YC�(I�2��_����v~E�\�0|I,u�חńm��>�N�4������1-C$�!��uۓ[U�#2i�S6�c 2��CʧqWCΰ���}D'�"k�v乲�"��a�TVw	өӫ8�4y0���|�4�	$c������:w�y�_����g�X�$f���%� -�T(4N����g@_>G>-�Y�X+P��i\����eXq��Y�T�S���X~C;�b��ОWظ(�]Y�B����?��
���<���~7jOT��#g�,4:'�#�3&{��0پ��m��l۪H��1;Q����(v�#N�����nj�&�Ͻ���9@�ՔIg3F��B�
4�)<�o�B�&�i��Ss���Գ�{�H�
{N�K�6a���� �գw��j��z������ބbV��D����8& �#�9�W�elG��4�_P?Z�!�����i93��#���}�c�U[xa�J�%E�mϹ������K�����2x��s��P�o�?Qj�5@����/�G(��&�Lɣ�!롘�0�?�ד-�ƥ�
�ּ����<g!|������B4.)Y�QK��B��x<�]�����!�ȷ�5�MIi ��� Ȟ#�����%t�=���pE^��}' �[^���]���K�ڥ��1��}^�F?�����Od�6���2�]�ї -!��T4I�+Z����N<�F��n�
��nR3���Dĝ����@M��
cH��7`ꈄ�?��Fꢈ��:n$3(o��2�l)�JQ�ӯ\�SU�[� �ps��8	�0�]M��k�������Qݲp���y�9G�W�:s���͆�+E0����'�Dg��]x��"�]����n�/~܂FZ����|�p<b
ނ�O��z�(�U�V<<���gᲮ�Y��L�"'�sR�F����]��k�q�U1m`1���p�ujYn�1�kmb~�Oޥ�]��}o���u��E޸-	D�����g�T��BF��O��u�*4�n�/�k�MUS�$߱��>֗�uWᵌZl���z���JxM��ʉٓ[pƫ�����]�U�5Qܦ=t�������(Ҍ����@\�R�n��2n����y���5��-�W�lK�o�����G��եŬ�4D�՞�7ݵ�r:G��q7��%��Ę��^�U�6S*�Cf�k�(�9�Z����O�G�m��ȧ��m���_�&���DY�����5R�<���'G|�����5�0<�����Y����-$Ŧ�@�Ţ����>�o%ՙ;����(��ᎏ
H�\�䝹��6�H|y8�
K����lV3Mw͞�i�p�˻ ��'�_�4s���__��^�Y�^|���5=��支�t���"���]�����LU-��Ik�1:%�	~��B��(;��#3�G4j�-k��iHCI> J#{/�D1�!�Lcm��!��d����b̐O���,�`��%�\����s����{ݪzo�n��g��`��04��*���4�R�>-��1�uq!�#�,� ��*,����Ȃ���T+z:8���7@��gT�0�X?"�[��5����x�[m�oO�iW�ρ���#C��G%�^E��StCu]N���p�9�A.��R�B��=��I�m܎cqهlh�+|R~o�!��ez)�D��� �8Xˁg^iCv�CO�ȵrHӤ��P�N�W�X�.O��o�}(�/������?g��Ue�qn	k�]���;������d��z\e$A��ە�+�/�SE4�<��HLs�����R؍�)����w������+xF�R�)p)�dR=u,A���Zb���Xx��Ս�.ޯ"�h�؉�HV�n1T5�ф��2�Eh�*��US��G�_�	)��3�{c��55�y�yE�F�"VO� �4C��kX(.I�<y�S�VA��`�<ݛl��ߺ�?�fT}t6Ж�7`	��Qv���+��n����f����Fw��Q'�4b�B�f=d��,ҵ����/V|<Bn,�ko�u�����0���r�
����$zDB�.Q?����A�1��F����_GUۨo�G6���^�|�0Q��Y:^�a�!�3ѧ���ab�B��f��ٌWf%�e%"*
9��xP}��^H�;5������G�D�:C�h�>����6J�J�D��lF�t����g(�ıb��BZ��P�6i���;{uj�*�U���(!3��N1���O
n�A��n!����� -�$���H��k>(���/���`��Rq?đr��EM���QH��>OĕLI;>$���ʴ��~=��C���ច��� ����*�ܜ6Qi�6��)�#*^d�۠L��t��B��Hn���7����,I�T�!��,̂�������4���,��ĸ
^����	
�·=���dH�*D�XJ
��A�l�q����Ԛi2�g�4��N�X�mY#M�{*�f��iY�.O ��۪����}���}�az5 �����^��e�0|c
6�(�ZM4Vs���k�Q�@�\]-l�#�8'8��`��cp�<�+]��u�<�b��Oߥ-�N�!x<�ǰ�+L�;<��y��&ٸ��w�&,~��4p�aR������b&&ڋP;/��+�X���3I^�=Q��(%pU��C`�����&P��f��Ϗ��?�!�ý�����jB��<Ҋ��h���E5�H��vJ�u"�;�IU�̓�+��w:ЬA
~`Qo��"��"Nt��P���4��v�/�G�j�&^S�E�鼵H�c8'���?ȏ  �W	@'H��μU��1�b�,��bA.��7�ྛ/(��3D�� k���Y�`���e<�����B1!cf��O�),��Hc�F�$����"���RT����m�%��f���W�Փ"�������on���'8N�O� #u.�{:�������b~ �#W��t>I�� �
S�;S"��>�����'.�=��J��d�i��u{ ���uA�g�������N�Ń��5����'���l���e���9��	ֻu����O�_�=�!�*�H3*)��/H��.g�"��A��J�
��~>�����gb�C'+K�fK���3>U���C �r�������ٔ����(���]���T]��Z}�:
��`�rv����Uu�������E���c�8	�'0$�P?"ƢWq냁u�ّ�(�)y�	(KӨ��ǱO��Z���I=�ǝ
┪}ŕ(E��aK�@�|U~�.G��%��>��:EH�������섦���}Ǆ���������C�@(�4%��+����¤��iU��MDI�6��]T;�~B��yG�G/�E^'�a[x\����������/	A&����w8:��/�h~��BH��J3¢�Y�N%_W�oC���O�BiJ�m�W�P��=g|��7��Ъ�Ċ��.���DRʈ���1���8�p�AI���xO�c?g�����E�?W� �EVr�O�m����>G���NB���և7��&#���QB�9*�3�gmL0*g���EÜ����[��2j���,����q۳��d�D�Qr8̏6�u�Dw�{���sy�� ΂�6���w���D�\�zk��5��
,�.�	X��;��&}�K���^�� �gg�Zl�3�?T?щ$?z�:�^�=6���54CX�:m*�a.C<�ʳ}�f�V�f�8�U]�a�`�e��N,�w������KuFAd�(LxI������E��:Rw[����%��1_��[ZJ�38NS��b\�)}�Oa�Cv��<����y���L�0��Ȗ�)��dQ&ې����,�eN�B�4��(Ԧ�@�tړ�,�D՛�2���-Kǥ�tܘ�A
������=��-��Gݫ� �ל���Ї|%�hI���!���֯J��N18��:���U��l���,��,�MK�Az2=2W����J�> 4�ŉ������S��! Cw��g|��&�~@�P�������*�M+��͈Sj��̠+��#X)�i.f�eߌ���*��w�q�����*`L�g����g�eN�ʋ�z�P�h@HӕB���C��K0��%��N~�ӄ~����)�)t�
V�I�eX�oɢ��?m�ɓ@��A���p�����PjXi�i;��{�uL�	�P��e�戀&m\�،�&C+��C��)o��=�Zj��R����&�����i�	�b�m���s�]�f�3hG^���� �k�a����ϞF��Ѥq㝅�r6[��y�ozt��#����zd�ʣ�;�#�E���A:�ݚ}�᪟�M������m�]%����:;�]Y�	������êAJ��d(ɨ!y#|�\��S�V\�����Xͮ]�t�%�ΝC���o��K7��U���)��ө�p�懃g��3k�	�@X�@PF�
��F�tB�K/^I�ۄ�_��kć#�F[�P���t*q�Sw����CV��Ҳ�{���h^��ꜗ?iJ��d@�z|���q��o'��4\�F	�{yx����&T�������v�S��y2
x��=������t��q�
q�t[�g)[���k^h���q@������o;@�	=Z��&��* ���>�����Y�	�V��W�S θN�%v��-"1�_�Q�eR������|8D{�<�. ��	&�q3`�^�����n��UI,�ו~4� <��T�@}W<��'I�����z��M�۞�ZAv�SȾ|��z�Ew`=d�w��%�o���4�!�9�K����6�ʹ�I�p,�� �d ���i<�vG�2ll���v�u��6�\� �@Ęl��o0�F��d�u2Ll<�S`X�-#���-�OI=�N��F����?��yˤ:@���5�o4+;�CaK�>�47lC���s�Za�zb�t�Mب������r<�ɗ@>���ؕd(������M�	{q��YoO�R�Ǳ��OmĈr랠��ɬ�ѕ�ZlJ��#��q�F��iu'�}�5!��W�S���;P��j�eE8�EF��n�ސ�7+ =H�r�@7��BO�z@Gg`��g%Hԣ9�J�⡒qs�
H�Ӊ�G��^žs4��ꡄ��#�mV�<^62��<����U�s�R5bY� ��f�?/���/ �>��4��4I��u((e�y�_nu���$u�!H3f�n);!��XlyLwܚkþ�e�H�����{�!eIݣ�d,�P��,r�J����I�]�w���kbٚs�c��[TS-f�Rc���z!o��4���t�P"y�i*�(�2�Y�4�(Bf� �X	�6�w�����-����ϙ}+��U?�m�b\�x�	<�g���x�k::)�=� \02�$էI���}f����a��,�jТU��&W�|S�U�ᧂҿVҚ[���)���QLa�GGjh,E��y�`y!4<�U��W5���y��I�s��h�O��uL���$ .�^�L�mI��1|)�nR�=��e���t���9����S�7�P=�&|��>����Fm��[)���������I�\��X��+K����+�����&�
��#D�A�<}��ڰm�{�ϥ�ЙgF
C'A�����ՔC;���h^���D�Z�2k*O,*�ҊL��+����1=��P�����ɒ^+l*�.eٸ��U�q��Y��3��:R�7T���E�-�6<I�h�d�[Ԉk�i]:���i2ǁ�s��{2�}5�J?���4_���\u��y#܏-�0��HZƑ��v��V3�ǖ����_��˺Y�-j�j1������U�B0F�]a���p��2t�*���'A�����ߒ W�d+$|���f�^��OKc�*͇�G�V����M�_,����CdB�w���Za�����6�%h(��eN�?N���s�4ҟ����-f� ۲��;%��,@�f�CƬ�My�ޝ��s���!4��y�3�Lg�[�!Δ�P��׿�Nm'���i8,A⠠H��.+��ҟ�ŮG�KD\�a�pv[�,|����րNE��}!�}���hŎD��X�=lO� ��Ƣ�zfG�����HSޣܘ�Mٲ�E�Zg�<I��'D�eǇ,l3/l|��'&�א�:��s;l^(*sX�~�Y&����WC�#���C��{��+U�&9j`;��W�qc��pKC�]9�#ӿ�v;���D
����F$C������߱��K���sT\�ם�p$���5Y?$�ꌷ3�^I�cN˺���Uтl��tl�D�R�#��}e�l�8�X��F@D,�˽0�>�m�JǸև6�W��ښZ��s1�W(��}XY���e�Z���FO�ڈlc_u�g~�O��o��4G��
Q0��f��
}��yG2���97b�vj�}�GDy��$N�iw��=5���
���������!JWӛ��Oɓ��k&3��ػ��'s�y�u}�J���9I��J�\W�Ve ��)Yd�J��,r��Ը`7�,�2�r�R�
����$�*������Hڳ��'E�&�l[]�X�]�[�nT�u�_t��q�"kx����3��t�7�h=f칭.1[��Zƕ/xG|fs�K®�����i_I��ภ\4��V��J��c���@���ss,�V�i���
�5vKF!B�������_��v=1��Z����
�,ځ5 	��.e@}�N]�ܒ�W[�rxaZ=� ��Of�n�=!� �Lc_��4Dgj�/��j�����}:�(��kÌV�	��|,�懂�^ߎ��5D81X3o��p�����;5�U�Pt�KU��O���&����B��0;n�����5n���[#�׻ ����S��6@O?�u�|m8]Y��e�����#�R3�h�'D�t�5��aP�T�2?�U���V��c��Ykf��l5��B�hց?��sU�T����rKE�@�&��ۍQ¾3j�f��7�F�����;����k_g���3�|�s� ����1�l�P���J����]���x��9����}�]o�-L����R/�m8`�DK6����ǂ\�=|��m_{!��!���x�����\)��Ol�0�Ց�R�N/�Z�:z��5*���:���0&3J�?ڋ�@�o��#���>�4̱"G�mƼ/��P(�L6�>+��n���.�Gf�AQ��#�A�^3(7�-����&:-�z����#步=Nv�$3=��2�!db�֗5���N�?8�"��vM!�r��#z|ŵ��a����?
�p�HD�*6i�.�|��%zp��� �f�C����b>�g{�\����B�#�ǋ�GW�p�mB w���)g�	(U�{���s��u)���s��:�4H�>��Ȁ y$��G=�Gn��O��p��ډϕ�Z��oa]�}z~M3	��oUfN@Ã��{�4T4��+�^yk۸�ri�U�G���y/�]U�7����X3%��JsOA0i����'[�9���ޤ4�m۱.w	���� ����Ŧp{�3���y�)G��rxe�w$��x�c���t����[�&�A��i�Q�Qd��?5(.6��u�~����cJ�Դr��S.0$�:��bA��ޙ��%2%n&�Z���F�& �-D��h�kO(nK&N�V������w �6��`-_P�ī�_6�Y�P��b)
��Z��v�e�mպś2����ǙN
ͷT��<�l	r�E�ky��]�a�0moM��]Г�i4���#5�O&I�Fc�nW�9)��=�S�D7L�l��z��	s&�2%��ö�z�����MG�"�E� ��[R�!(�ndTK�ͨ�0|�U�����}و�#r�*�ǯű����m�e��d� �7eW"y�pR�V<ӳ9M���ꩃ�,2��_7V���fK�R�����'pyl2�cƅ;3"�w�'���=��j�d|D�P4�?�B
����+���f����hϔ`������+���-��N�O�A�����$�ݯ���=�~x���5��ZQ�BX��2�����
S�9]7-�F��Q^�!��X*�J��O>߹��:ڂ.��������(�k�H�@�A=��L���%<PU�XWސ%؛rlgd��-�-:4}��*]`؛.-��r�^�H3�����?�=8��a�����J"~O�-�dN�<^6�<G��j��p.���!�I���X����
��7SL��΅e\�M�V0ԭ�J��]���U��/����4Q����v�pஉ��>�� ʙ��붋���G�[��ܽ�&���[�;y�x���%"��H�jf:0dW��[��#F�t�̥*θ�S����>�k&W���=t�G\�T˴�7.4lKY"��]��Qz� ��N!�ȕ��`��t4����U�ZL���>�������ή�dS�� kO�3;D��w���,_P�3h����Mt��v�vO(��t�І�&Ks��_����j@x�Ӂ!T;t~q�r�'#|�̣���0�А�o�>�m��K樶x��	�4c��{tY��T��Z�<@��*�+�s��<䇶��5�pP0<�a�A����^2M�N�3�"e��O��{ѐ�{;��#���q��;��^\yQ\y�nO�>!*@���`��-p��O��?.�����$W������'���5�����ˤ��69>;L
�U�)I��u� W�?���z
������gs�~0;�����q���o��և���e��k��3�;�~�eO;�P�S�h��Y�3�]B`[�9�>q@�����
��x�଄(��fO5��rN�5�������m�I��,	K\<�����j~ϛ�v�IΠ9��z����X�7�K���<Q����cu�p�0�O����t���˃��Q��&��?k}��,v�%�"�����xyfv� �����?o��F�;��&(�$EΎ��x;9�}^*@���9d�}b_7�=a#�FP+�c�'�Ie޵H}:����k�h�W*Ry�\�p�g�
`�n}\x>�K>В������#B�(*�3W�u.U �����+!�&ɑ�$ʹ>�$�e}����9<X-��jyk���ov5�ǡU���x��p���3�b�b����p���˷OwO3��{�,W粚��!�$Ғ�O�޲��T��vQK���o�g�Ī&���@OkP�^�nY[�i�$����dg�e./)L�E�ԟl�hx�4Vv����}|y��-�4$l�Jח� gl<-����T;������� �鿼{�����������..bQ�?|�b�NB㳔�d�xkW��849T;k�삉fA����fL�:	4���&��5$�C��כ�����,*%� h%�ie�ۓ�"��#�.%�a��~���8��if^���ٌp	�!�~gi���wO�oY��2�>6g��P ��jP�խ�=����V�B(�r�yƒt%�rױ��~�=�t�o���(C��ol,4����Xy���a�j<�����9.��S�]A�����B��t`#���5��ģ$O�����S0�H�|`������WEjD��~�W��Z�O1/	�*�/�T���䢂�%Oy�w���Z��q5ZZ{\�+�}W�g���o��`�!2j��VL>JRV?.�!\l���e�H����Oj:T��� 3�tG�.���덓�dvB���!R�i��>�B�4��-�q�:ֿx����UZ
#���$�*(�È9
��4R�(Z�x���xM�Պɮ)!�L�:��ǻ�k��ŋ�lQ����`�0o��	�y iųZ��l��pE*
�o��N(q��I�Æ����܎a�������a��A*��wr�d��K����g��$!N������Ș�I#�v2��`����-�I�즣��_�A��e��3>���+��o��.q�N>6Y~kAm��e"��<39b^���ӸWʁp�D[Z6s��\�#?%����<Q��2~�Y�.U�����?� A������f9+ʄ��F;@Ѭ�tߒ�[���AO�����*����6��4��\xH��3@6�d�����@z�(Y#Zqc�I���DO\���`Bc��8��WцXu�@YV��و�.|�	���ۢJh!J� ������d���Z�~�f��~^f>�f�ܯo�R�.�_G���@�ֱ;ܦٕ�?��ˊ�>!e5���� �<8��qV��ش�Sr�Y\���{�� ��_�l=FY�,�5���[����7�!�|��}<�8"�J�Ĺ�t5敤tq_�4��P�t���:=Dq��	�9z
�lU+\�-���7h~�?���BX;�������]�e�b}|�M����;l _gLj+e$��~�TO�ɇ��~.���=k�k�{��3%�c3Q����g`}��4}:�E�\���Y��
>����[�楫�V��/���cƵ_���&_�MO��i���-i���Gj�W
� Ǳ�����MdJ8��/N�����a*��Z�> �g���uN,N�ᴅ�Ђ�����g��Y�+�fV+X�-�H��?�$vu���I�Zxqe�Hw�P��z��=��x�J����݅�&��d�E�ۘvZx�>�9=��<*�N.��o�O������*�jd�b��6����b��yNūܤ	�<��hߣ'�U��>�wA� v�	{;�҇��v%��F��m�:�����ǝ�!n	��R�����7��j܍i�
cЖ%)�������UX���rY2�C�ن��bE��ᘛ�Y)�ſ=|�����`���pE�����$}s�.�b�Ui�����Vc��r���� ��h�
�ԧw�1Ϗ�Up�ZF�3�lդ=d楀u�8iE˱��a9�c���g��?Dx�RWό7T��~�����r�G��k�a�N��˒���1^ �U�- �w�������t�\�	�zp6#���^����(�ru�d�f�^R~�|u��8q �!�35��>�F��2��������i4J�Q=9�m��[	"�"�z�z*i�C�9�$:���}���5U�V�9?5���1R8]aD��r$`�s�j�����w@U~~�rP��1��5\L�>~�"�����E���lk��tP���X��lrW�p�C�Y�oyP��zJA��n����k���R��k�=��>����:F��cǏ�m�Q��ա𝩚c ����#���pi6����nWwZB��5�*W������U�X��g�哋�'��39*�S��G{������d�Ԟ��s��e�\;�Jbbq�H��3�����%�Ҫ["t�t;�D�R�GoF�߆~,�BJ�E��u���1��e*�7�A�v��xxb�ݡ��IOzjy��n�U�1mhb����7g��l.�3��ix[����֠�ז��a���(Ksv��K��������!�%�K��̞�P���'���D	M&��.�@�	��;��o1��Wg�*���J��4�^�;e��~�0����5!��7mm������)��^7Rǲv��f7s��ֺ�2fx��n<���O�խi8뜒"ݕV3V��j��NIr�H�Q��y�6�+�?9�{N�k��&���,_�-���L��˹i|Ag�L�I2
�DO�<Ūm�x(�����a���{��/�>�m��D�s�H��ƣ��7���aep��La	�?_�EY�h�cCiR�����Ɨ�;�� ��`ۣL�)��t����ʗdB*�*��zr��w�l��V�S���J�+�I�k���"eՍ٪k�H��p{�C1a�kZ��]d����>Z�Tp�:�M��/N��R��ˣ���ʇ�(���m'�(�� .5���_X�~y��&�"Sf��C��J�"�is���#u�c�*�~j��z�B�j�=�jĆx(��L��K�<T]���5���Zxړ��I;c��r�ǁ��S���}�F��翯�٪Nb�	�(4 �hK�!=E"�n5c�����T>�;�W6�=9���F��~e>kO��=b�vek�\v^G�QS��>�����-�u
z�@^��t"$;����@6�'�d�,����^�xCt[s�'�:R�������ً���&b4L��;�̠����'3%��s�A#;oI,6��>�d�A<�^�#����*ɦ!A�#���ʈ����t�N ��(���H�����.�� n
��#p�=�}����u�UzǽJ#Dp!CB�e�i���/z���"D�����^�̂9=�F���Ѩv�5�6��-��X��xu-rg�E��� �_���4���l����S���>�z��R{�L��Bm��>5*�
���|���Ad�#��O��Sh`�f^DN��^�v7
���E(�Z-�c�(��>~�&!gIJ_�A��y�5�g-X�A�����JKC�VN�H�5����r��(v
�2?��!-�����ȩ��(� b��`&���R��wJŮ5d�k{�Sc���@ҕ<����b�� �f�s�w�)�M<z�_k��@��������t_�$�����p�R�c���E��+.:�.�ı��F����r����j��<��>��xh�j��P�������B���@����lFʟoO!���B>y��G���(�2vD׷!]�V6��Mz��);B�8N+���jQ^ދ�@|�B�9�f,��#���~G��`�_���c�,��uɿ�x\W!:�; .K]/!�ah*�EDHL�Xd���"�#�|��a�$���e ӿ%[�o`��-�.wx��+�S�[��a|FC�m�@�����B����מ2��x�v����.�GL�G���qI�f����t�{��iyݡ�����wB��&�h�SON��).�j��j�+K�W�7��v��@�(kD)��1oc���R�yn(d�ܔ���� ����t�������1?N�� (�-�?5��ڠʧ�H�'��̝�숹:&�Lm	�G�%��|��9I��,#y�و.8��Ԧ��omgKC�� ���-ᾪd�dPx]����8��_��B�OI��kȬ�J���5�(���������V���nZb9֥��F�[�w�ۍ����-�T"Fw�~�e��k�OCL�
��У��v���� 1Z�	�Z����ZM S�BV2k��M뭌t��%��G��mv�����U�q��Y�@�i�1fBg�E@�e7�v�+��Gy\�gRv#�̏ ����q�<I
�ژ�f!��8�P2��;+�ҸЪ'b��z��_��]��ʹ�G����`a}D�)�SK_dĽ�	5�
�YH��i��'��Խ���G^��QY[����n-�T��
�r�]-=�*����J�~��x�x�������E���v�RW@%b���2�}�|V�?�	*`To�C�mt�4��~��E�tgt#ܮ��b���sTT��(��m�7�������&Y?��-�z	�����$�:���9U��j*�� v0j]H$�����g[.�d�G,*���7M�}�a(�o�[��\�DG�	_���0��Ǎ);�J�՞�=Z�������ΚM��F	�^`L����<������[��A��>#��ͅI�Wf�#>��Bj����x)�i�_s�ʾof����[���r�<�\�%�j�vu�X8-*�#a١�ۏ�u�
J��rd���8&n��	7��\;X���l����>��:���.��2��o��W��qxTz��[X�t���΀��w�z*{�	���=$0��B�۸�O�0��F�-[��*��3a��Y:ďD}m�Ћ72 Ҝ_Ҋ���t>��K@`�)�ic��e7���%=f?��A�r�B!��m9״��~�p��6�B��a���x3�O��"����T�La��{���O#e�@n��B��ȕPi�d�����A��/tT�<�6�Zw��7�n��Q�%�l�	̦�8��ҥ��V���*�+F��X��
5���,�*���"ւ��Q�(�w>�:�%r�{��c��.��2��(�<�*��B�*IQj)S�x��e s�s�G�.7)8��Ȩ$�ǽ3�2�kB��J陶[X� �_���A�aӎ>�8�r�{��u�~O9L7οy}���`\M0��t��Hۙ�B�!�!�\��&��'�n,I�cvy������^����:#u���'ή�7@������	s����y��~�.>����"��S�u>L%��~�M�%}��C/����)�|���f��AK_�*j�:I� �"�&b�j/��
Zc���H��d!�[8�{�p]� ����(�=y��A�2 I�E�����3�*��{�Uv�NOY���A]���J�r'd@ꩨ�4{�V|ZߢP���Z��-��A�'��b�l5L�	шF(��Ӕ(S;�؆������f� <a̧�"yr��X?W&�>;N�U�V�T��2D�Y/�j_b�M)A��1�k���<Wm��ɳ��@��Q˓9X��Tp��Ǟa�B���Ae26[��U��e�w�����M�9�m�����+�T�O�=g����5�4}ު��a�pLLV:����Ux�vl��0��9�a��((VJe�s��=���@�Ĵ��p�E��]�!nctVQO����Tw�^�Ԃ��%���%\WfZ��_���_��>���%�>��\��
TАR���E��5`q���� ���?mi���H!Z���j��/�;2�y�`��3�@�7n},F�(Ǝ�~�L	 +�^yB3�+U�
�����(_}m:NyK��w�����+V^Q��J�!ywi~��5���������iU�������*���k�#c��e�ۓ��|��gf*6@)���y@O|��=|? �$c��Kx�;�s���������}��H���-*6R��!�b��#^ݸ� th��A3��ѰeJܔ��P�?Ek#<��H�&_�w�򠲡~��nN��1y��ꔕ����&��e�ot�C)XV�$m܎��[|�mi"W#țA��d��J甆wI�R��I���$�m��n�7�e"��O���Y<[�eQ��Ly'� ڊ�<�l,�(9�o��[lF���H�a�zW� -�"����EF,⚏J��������@��ͼ�EN�}ˬ����p��ȋq岱�|!3r;i��cF����?�&[רwT�O�-�}��)d^��a|.IP�2-���eB<�qP(bX�����%Y }��s��=t����P撌�4�-Qب0j�F��s��5QKW����ς�-�.m�$�	FxE�{�S��3$�F��9R�;�2L�[ =���~�$m�x��eVZh-���"QN`Xɱ\R��#��![Z��?�{e�5�M$�(n�۶� ���c�dvc_s3�ˢ�#�l��<��{�Ț��~(���(<JJ���ʃ�Y�m�X암Q��. >�B.���<ɩ�D�dp���O��P�h��hi������yhg�#�!*u��c{��L\Km�$���'/���rXUKt���)�!�0�j�k��@�R�񸎀^��h�%t���X8{'e$H���z
����\��{8��Qu����x�+�����ޗ�?ז �S��'�YUU�JѴ�bxPm�� F�*��){�#Sd4aƋ���O�ؑ/Fk�&:C'�㑦1.�F�j��FAc�'>�>�ӂ�J�Ë�S��$|����p�'tD���Н�u����K�_�|�"���� ,����6O���o]�a7�m�Z��)GӅ�"�8�<x��+��O��~?���>1�g��6�t��dc�1f���Z�@~e#ΫM�|�	/��¹���֙7:��Sw0�����O�_m}9�s�D��N�΍��w�5�X�{�<����r�����H;�52��,l;�h��0	R�Q�W;
����4h.J}�	Qz"|�	��$�P���ǽ�p<Ś�y_=����;[w'[箩�9�V�aPa~aag��%��V�x����z	��?Sf&��B����W8�y1s��5
��W��d]{�e\p�~_O)�-g&�k�W>8��&-����c��쏅ؔȡr�2y8�<.Udt�;M<�[c1����͉�:�<��[�ӂ\�7 �f��������M@0������ٺa:6�t�j4)��"�?���sl��V��|�, P�D.k��̰� g9@x��V���;BT�v��ի�� ��oN�Iϡ}��^'^ ˒��T6����#����`*�������jr��i���PH韊e�v�0n��i(��k����,m���FK�U!���?8B���V� ����dї��"=���0_Eۈ�j��(�a�����ɱ��ۜ����x&\�V�K�:6�����C������{��Ҫ��j���LΜ8g��7����=�P�H��Iu�(��OJ����Kk�t��U��WM�`z2g^�'$�a��`f����*�����W�l\�����F������,.���+Ct����h�=�Ґ�����I@����4j�� P��e��g��E����!�6,�>�cΜ@\�)�V$1<�x�����r�Z<%�HWǣ�濼Gø
UjO���H%6;Ճ�x�}&+����"]�^F4 !+Y��-ԡ���UTn���a%j��v�*͘�Ԛ+vR<���r�q�zq�ƙؔ폲ȥ�<m��5a�*%��׼��p"���]�̀"q�?�&td�#�S�+tý���Y���k�_ri��^.���"cU��`�=-��A��7�T��w�5��C3�=�J��&<[ƃ��.��b��?5:Dy?_��])˜d��O�KD�ΐ2��Y9�{��������b]��0\8��|�9Ѳ���B�Hj�6k/��T�>N�|��VOYG��n�E|�C`��8N����s(O�ivp�X�-3I���W+�|^(��?�&�4�M}��L��V�:F�Q���蜥(�7N�w�ω�p}n1��姻����i��L�տ3��������b�Y�E��r�4�Gݺ>��VrD�|�����^!l�O8�"��B��`8�҆u��_����%�!�a)��l@nG8����$o�e���ׯ�'�a)��`�y`���n.���JԵ�s�Dj|��6�=� -K��Ht�)@�L�*�߅%G�yQ���	mQ�5R����UZ�}@މ�mb0ȋyy�Z̘F�Ao���A�8����~$�t��6�.��u����:��)�����N@��s��G�Q�t�S�'���&>8-�pߴ}Qy�=�b�ݺ��y�|�\n?���:���|����K���L�����o�J��j�f
������WD4��� 6y�A~��F��+���) ؓ�(�`;U���e��my�3��N�:�V5���α�d��n�5�c�l�PX�6(==�3d�}L-}W�T�蜽xt^8�����è:�G �Ve�FZ�zٜ�&o ������Yg��) wo���;�6x��A2�ͳix�gvf�	�3��÷{+�
UN%��ru����N5�ɚ�K���<��NşL,:S�^��3�m�����ı�6sSFPp[3�2YX�9`莦��Y�*�y=�Z*8�D��L�˧1n����vcg%+�E(��d=�ZPA�Mo����P��<PS��"�4G��@&�6�������9��nA��JM{%m�|
T����C���-b�E��_�M���JY��<���ɸT�e����Ӛ����"V�㏚��R���د� �z#���t��l(La�p�b`�W^%�_����o���dXsb��K��v�WN-�0�]G�0o�y��5t��ҹk��|���lE�``|�Z���YA�^a�ʙ�^�`�щ$9{/H��0�_������bV�i���'|���.�2�w=c�d��jJ��z{b�3w�D���AĈ�-	BH�-W�$,�=�!C��@���q�Dη7�A<
2��5W�k��~a�g��@]F�#�;=���'�!�q�G��6�I;��f���h�`��H�/M�]�bώ�L��d8�%3<��̾��E[�b�����V�j͇�F�.u�:�.�J�q�ֽ�N;�͎U,�Y.<��/*Q⺉H���gh���D�3���:���� &}�Da�Lb��]����pې��8��{�w�*����g�ڏNDS@Sύ�&�����aY�J��8)ϕP2 ���#96sʽ(+����S�k�����h�x?�	�Nx�6�m|q	ծx~	�$=2�d�%ǟK̹{�X���Bg-pJܫ!��5_>�_��Y#W�QOx�q�84���n_�Zr;�L�b唍��jn�_2�Ƙ<9���_F� ��:f'�;�	y�HE�@�+K-��G)����Wn�wP9�'�x���8��;�x*��"�D�,3i@Db��|G���cH�c=ʭ��PR�c�h�bDT���?]Z=��'E��F{ּS�ŉ�(`�XO�?O�̈́N0fX\5��N��b�׳���"��«���95��;�HΙ�w��$�T��S�^Oﳫ~%�/�҅#p@�ATM�2��;<%'4hmq�����r�����4�'K��c�K�x�H����_Ț`��b�2QB)V�N)������q�]wl٤O������+佝���� =I�� Ќ��o?���w��R��ݩ#�8�(ϐ�ܟ������3*�h�3g�xf��Y�o5Z4��mFӪ��]���lq�؄@������`.�df������s���t�59%&,�v�.W��$ʏ��ŏ��� �#P�"��Ю�u��N�$�!\V$����U\z_�_���A�a�NB�t�Ӗ^p<���������*�ʒ��R2�,\9lZ�t�W���WJM�i]��/ ����J���S�A�h�%��7ց�,� ؉�҈�ā�?Ib�`�'�.ͯK~�
vT�E�ěi�)Q#�����u^�Ւ���@}�%�?.b^��/�9k��¥����I)ѕ1��_�Y��B ��vA��q�Rd|�UH�G>1)GF?�I��=8����Sթ�D�0�mH��V$�Z�2�okS�~7q��l����U�l�����D͍��6�h+R���ɣ�M5�������U/A��Y���(�o䆶�p��ۛ���F�\B@��	3�}-k�0�O�u��;������鈌،^��z�����f�/��i�Ħq_�d��%9�ӽ��� Ǻ�1~.���h����+�	L�����&R�U�u�'/O�DH��ҫ$yw�K��z���\m�Hs]����<D�כ���B�*<��́DM?�Jl���7�O$Ĉz����}��Q�]�����kD�0dۋo�~c��We�S��kt89�9ALg�^+r�ho��g�<�Y�;�j"�i~�}��P:���H]��vn���v[=��튪Gd(���WLH�Jy[?:��K+�����%-�|���c���/�����!+�<�z�_>p�,{������yư� �[I��,���\@Y) �۵�d"^�#�G��b|����IZ�:�����NzZ�L�-43����%z8"F�_H�0ř�&�, ����P�G���A�dW_���|	�+�5q���c�x�5tZ��L�ں}ǭ���w�8��4�0O�AU6���q�r���G_g(�ƁZ�-�{��׿L�8=�(�]������d�����2�O;n3��C+E�m�2E�H�W��'��+~c����RdJ�h����&O��껣'��eؿ$2O}t�cvr�b�c�p6�Z*����w���6���E�
4�PCX|�6���|*���L!�y�f;	�y��f���k�V��^���\��@W��"��Io�����qIǪ�gT���a�bFw��F��s"��W45{���W�z���tMJ����|\��k�r/��#�X�kD�@jTÄ�D�3nhH-}�/��j�� ����7�X��u�����4P��w5�4����iy���D��rlSе�z*6}:]�S��ȱvf�n�}�;�1q I��O�����Q���H�*R�I8w�>!��[��չ���Eo���(��y�_ȵ�c�,#+�pKT�rK� P�vO����jT�c�v�S�������eJ8X�7<�4��$�fn3G5#0�l0UIC�<�?4l	�o�U����be �+��oZjG��_��6D:�9n����5B���L$�/��g���~+��'{ʤ9���c��6�f�
;v|$�{��j'/f��hc΀��߁�����f�|����x�t @yb��VM���Ѭ�[pR6����[eF^ʮ�$��36;�����|�y�T�*�X��61���;�0��իR���H�yQ*?�e ZT!(r���w~D�c@��ep�"��J�j ��k!���"�h|�W��+Lw
lma�W�}���u��oA@��70W�*mӵRgc��q}��j~
���[V�ш��_~/�T;q.�gփ�]�F>�
��׎�����zKv6F�������h�d�*D[��1��Sw���3pΤy���[���B��!��n�}E��r,A�����*��d�Ͷ�X�`d�6��=~�'P�BB{���Y��W����4�9�_�e$��JG����vzw���O�<<��*��Fr)Me.Mw���`��m�4�a���$�qL�������[�ù�H��/�*E�a�C���^>�L�;-;Ls���)��m8��LiZT~�Կ!��9���M����B�Z��T)<�5�P�,"�g;��=Gy�{�_�h��fP��e�����U��V��Xh��|[VQ�64�B�RC<��*A-�Vѝ�W����<����Y��dc ��ŀ>:���L"�9�n!�� �ƌ;(�x��@/���b� ��`yT�N,�2�N�/-p���y]��x<}�ʜ�~�A�*��,=[��v�t�[h_>BFtj3�L�@�UHO|�l��&Y�9�R9����wi-�/���}5r�<ua��x5c�L��sZ\N��7"������s�7If(�^ӳ��_��w�
J
�Np\���]M����	�ZUM�f�Xn"\�3�\fl5s(n6qfؓh���7A��Y�s��fA��7��;���p�²�؂w"~�����`8G<���wu�Z�\[h�؋�08��J���H��M�҆��q1c�ϓ�40B�t��o�dM�@�V�]��7�:谟	ڤ$itU���Z*����gh�hdܿU��������Z�e�c�hVy������l�3�9��}�S��N@�>g�{��%i9�P<A��o��}Xǜxqo�
�
E%���z��P�`h��L�"G��E���E0�����F��(�~T+�]H�k�8\�� ��	�?�h�|\Z��"M�W4��Z���u�̾41ۚhp���Z?��ӿ &`-]ǃ�;�=�k{��lī]=o%\�h2aȩ�ֻ<�I���i0�4A&t��4&�z�$�Ƕ*�����ϋ�E�'�V��pPg��A�������Q�	��><�F�������Q�ۦ86b)`Y
�,�Cף3�{�x�)Tև���`5`�,o�V1͑4�J"Z�DҢ�1PǍ#0���P��|���f~'��	"�VcI� ���W�@_�wO��)Z�TF��[K����\���Q����yD����d����"׶#gO{�ߎ��=u:��4�&�[�b[�����1�%)ƀg�"8�_Y<�'i`b�OV�Ǳ��|E�o�:�n�>�z������]*���sD�ݪ��zeLS����c/J��*g'F�&6�Ù�����F��� t �%>�;������%`'�&s��<�0,�=w��2�cK�'���\c��Ɔ�>���6zAĨ(�+]Qٱ��l#Ʈ5��8m�$�mw�T�yU�h���tY�xd31h/�Q���z:��ʹ��^�s�ǥ��/(S0�O���S�����ճ��T�:]��9AM�(�l�w�0��	^Y�3ZְJE�oa��������T�j--^�d�C�[���:�i}�
��B������'z���6���:�'㶡�x��?H�M�8��U�(3X"�����h�>"/Ef�	8�A�n�j���#i&���~�X���y�F��
R��9��/mɜ,�X��y������٣٫�o��ʘ��9��qЮk�.����t�9�7k�:���^�h�ux�Kb��X༑.V9�*H2x��V:;�{�`$�q�mo�2P��i`.x�?��*i�9c�X�zB"���B�v��)*���|ϻ�R�aN|�j�肽��fQ/���JP��W&<��'��p�V	^���{�Gqx���R�x�����/ig�x�������L�W��Bul]{_�+��!v\�+!���_�e��V�3u���`]E�	��g�rښ���l��gD�|�a�7�7���cF��y:�M�ւ���qk@ײn�Y3Z�P����j#�:�eN��A�#���̦}�\_{�M�������V�� 於_�����2�tbt��*�ϯ�;4\�e��w�ͽ����݃� s�h�?M��G��J�z�o����ƭ��K7$��H�
���k�T�Y�գ����	[����GMA l�ʟ�4�����$�YQ�BQ[�<�SWʹ���R���|CaI�!����G*��G�1Ѯr@o��A���_*0�kۂ8�zTz0�ND*�\���p4�� �<�/�tOe��������4s�]O���܆9��& N[��l&�\�	*��l��K�A���VB��Gzf�@T�@��mJ��S��	}��	�8#w������e]ٜ��Nsu/�=�����U>ByNN�k���I`��K�D�������̟�vH�,?�+�k���B�+!9�j꼈�B;j.�8a�ӵ�̠YHHKiO�8�˗�E�ȕ��J
+����0&:�N܃�(�6D��6��
7t�y]Nw�6��j�����u��=ܘ>h��z�c{��K!��XWOx��#�.����֥#�F���;�jm�6�@p̨Ч��]�u'�� |��@uɈ�wY���_��M@[j�'y����L�D4�N æ������)t7��Z��&�2:F����1��d�$�$�C� ]��}Ǆ���������c��8/Q�?�=c�Z+�\�;��}_y�����N4�?�>H<�����)�z�` o
�p���6��k��)�$�=�?)���[��+)�FNO�B��q��V�c�
V��Ѱ�4��}�W>�;|]<�%��3�ZaЯA�ZyH�����������7��@�5�w)��˓iZk���ס��~{�9rp���h��wM���(!�f W!�b��1ө������ٯ7�y�B��Q\(������C��r��z업`�+���D�/�.&~?WA�
� ${2\j��� ��i\�eí�I�(Y���c�	��Z�*Z,������D�����W�2�f��4��}dvLǵ���<'ƻ9+�����[7"�� � �J%z��L���@=�P<}��Tnޅx���̐�j����w����M9;g�(�\�i��kN�Oݢϓ@P�ȁ7@.�e�=���ԓ�R�?[�B�!Դ(��p�����.k*TF;��M�\��#&��#����/�� QWm���O3��lq�7M�a����Bp�\����G­J����^�­V\��\}×}�Y6b:�h���FC̸�-1v��湌̛�)���JݓJ�|q�A���Z�~�Χĺs#̕��T��ډ�������;�M$�*��G�g?�� ���?mT�%�Ui>�5Q{τ�����#�l�fd�6�@mQ�z7��|38UH�1�I2b��ǡ�4��R��r���o�YtD�l�4�%ױ��Q�F �c\F�������'�z�z81�OW,��j/'���'�Ϯ�� [��O+-	��BW�����r�r�?I~|������d����C���>.��m��'�r�[0UJ8��n:���O|9u-P��C/v9_l����	ʶ�đ��u.}Jj i[�M$��P��KW�������ru6��a�9�K�������&"?ȧ�t��9n�����?�����K��ʬ�/Cw:ތ�����B�e��+*<Tc�����-J��I~�����	"��yʞ�{�(T�L�{4�'�\�W�{��ѵ|.R���@t丕�#{s�n#L�`r���'G�D��~�����	t$���g#ɂ,ʷpJ�=N�q��U�5�ƞQa{��&�9���_r��ޮs�{�1a�?��8J �Kr��?E�ٍoƺI�2�q�=yc�lw
�*���9�j�	�>t/:��Q�0nn������,���)�4�͕[�0�Vr��X����33���7�|�K@��w�c(fJ�`�丁�ĥ@M{�<�l2_{�W�φ�=������J��R��ż��8������~�7����D]R2�B�"~]��q����s�}_X�zs� �U�"�4�m�T�vV�KY��i�?}ʎUJ����䫛��#f�t��te�(D���=ɿ�u�0�����s�����6G,��DҲ}��$���c��ˊ8t��6]���� ��gZ���ٕ5		�������"BU�I
x��	��¦�I�r"��c���E`�����F%&�F |��z� �@-�d��{��@��*����T;� �vd ��e�EA� ���,{�h!��E9�!������L�E��|�H��]}�,��5^�x�8������L8�ap�.�4l�V9)
_�y}���П�'N+�Qf4��E�A��գ5:NW(��}��d̗n��T��d����ֱ�2�V�V���ē��u̪����d�k����+|Yܚ�Q�X�'��Iv�G��z��a�f�M�]I��N?3�=u��5�C��Y<<��7���s)�����Dl�Z@���=�sv~�dU�sԘ��V��%�헲YC^`��X�w�Sz���]�G��l2h�`LL '%A2���{N�w�������3rK!�u���ql×bܟ���$�]��~36�#P��e��Wn!�E�E�j67��V|ZPcU�\mV�g��`�F_�[O�O���5ud|qD1�+%�H�����Fj�͡Px�RI��X��-�9뮰Ë1���JbR�>Y�g����dHK܄C���-CiM�:����r�X{/d��4݂���0�A8e�e��:_�{:�/�l䏶��۰+�p�W�:H�S~h�P0;��F[���}7�)*)�B}�[��}Sfr�t�S��͝�p�� );&@���#$��㤭�e��y��pr��W纅v9h�6!�ndvZ�NH9�s@�v����[u����T������Ku/�	�r�RI9V�؟��moU|[-x���D�O�>eBe��e$��tMi`w�FK��/-ه�9��o4&T��2r�T#F��M�|�6C�����NL��)I�������'a�w3}�%�=K�&;���?�S����cO���Q��<z�:��E�T�e���l�P�z~�	��;L�z�]�`�͉�'�i{�x}�M)��0sN_��qOg�B�˩��p�Fj���ʿ�ǽԳ�DGPĺ5;8Y�L�g"��j�&W�9aۂ	��kR6�5���<V ��5��ň�XHe�fV���̹�w����͠^̕ش��o�);��E ��Ї�s����}��d�Z��7o�m����%t�9�l~*NL5�8��ط%aIg�+_����}�Wn׈��:�NOb������'հ��J��+�!AS�ӕ��\�p�:�K��R�wO)���{�R����K�p�ñ̪�g��i��ws�9�!�h0}ǣ7��$q��>/*����7����L��T�R?���40m�N�^���l���~e� zI�$�e��qT�J���ϰ��4�D����Z��s�|��菋ETH��.iw߹j%�øN̰}�1j6�&ރ !D��<B��.���v�����:���v{�kҊ��COa�L�\����\&S.�b���]�D�_���\��"}:��ai�ݪ�I�����L<�G����]?<S��w��1�`\��Q'�Y�;�o���ӝ���C ��M�((�s���w.�0D��f�8��;Bc�S_���f���JlS����ʢ~}� �R�2;�*.i�*x�ɪ���ܑ�л�z�RRk?jr	�x-�W����djG��r8d~(�!�'TǶ.�'0K�y���XZ�e�T>�ߖmy,��=��OLϿ�B,6X���z�c��M�f��ֆ���O�}��av�;_lE�)�(�~�A"~~A��X�&<��O��P#/����P�y��}�;x��u�_Coz�xX��l���y$e��ƺ�:0|��cO���L}�)������^4=��N���0�?)p���hwۏ�G�45�Qf86VJ�����m�\��j���T���F_X�q��ޯ-���\E�>-�\^fk�;���>VD��Pyx4�c�n
���؝����sP����R��:t����M>��!��{��
�TG~Cߠj}z?=(��ף�1 ����\��w�ŔYyb[�
�**%c�3,�Vf9�k�G�c��0-" }�=@@�~��lF�7t"ʫug��Bb�� ����ϔ�(��D/>�Ið�C`Q��C�d|!t.�e��ȅ*=��
��&X�F��.�N�*��2�+��A"��3福?��~�SAhЊ�����?����[@x���
P�
��-ݫ��N����7�x�Ŋ���9�\��kծ�����l�<���9t#M�[ANZ�4,�ΣT��~�=8͎�f���NύHE‮#nM*u�T��jG��K*���$S��b���pi	�rs�	���2���NZ���H�E������[���ia���с7��39�8+�:4���y��3�k��BOp�#v�	��~5˲U�62K7P��ڕh`�xځ�Q�����g�A�%�,7~8��L��>���>��M�:J��g�I�!�m����r��i$���(&���:~ć�9*BJ)?����1WY.�+���5#x����>J��:I��n,m��u^4���쥆&}����Ԭ�m����}Q�^N�-�����HTM9u	����֌2�\ ��X�N.�@�aT ��6�zD�0������k�����h ��F͠k{}泊��i�# V����#�H}��"��pQ���W���/�a3B+x��(Ъ��πV�ޔ�:�IH�Wio��b8��T�Uk�TY�;Z��ԢN0�h�-�8H���u����BT�m��p|٪K����O�b��g�N�t3���+�pkp�9�Z<"^i&3���A���#d}�P�k�@�$���UaG,���~���ѓ����1�(z�E_�L��[Ζ�5� ����н��[o_�����06�"l�}���- YؾU�W��j��P�?���l���_�Ki��\��1d�a��"�U�A�`-$����[0��fܨj�2�N�"����u�o��qZ�3M|�9����bK�؞L���L��a�-\_P��#̭����*��-�.`�K��+�8��h���&{�oX��h�nA|Q���K�h04���Nr8D�d��VyoԶt�ҭ��4
�A����jLIߟ���S,+�q�@a#l�Uxc-�S)�X���*�1���7�B)���Ϩ�?"R,���O�(����]����.���~�re<�s�K!�t�Ȣ�sQm����j�j���h)ՈX~!Htf��-����z�S�?�XQ��#���Q���p�]��a����>���'V4���0�@DL*����0�}���NJi����ř?�C���>��6�,���/c���:L�(T[���Ub�,2�w�]?)^ء��N���i�+�h����[��Wb�)�:g;��X�WrU�}~���e"��o��*8���"�4��PR��<{��8M�~?X*i�ө!�78���j{o~�E�,Ю+��3���C,4 [8��[�e;����nN�:�N|��{����1�h��� � Ul��Yx+9DP�dgڑ�?'XZ<U���ʵni�zuY}&��OW��r��n�n �B�m$"*��]��_B!``��0"��6b��	�I~qy���ۄ�����tط�	o���'�N}a�_:߼&n���}56$�h�)8�N|S���)�@Sv�hDpL4;/���䠝���%MΖ�`����4M"L+��%)�oT�n.P1A���l�d��2���QhW���q����p_�˫�w���`� ��V����2�Kt-��Q7fv��,�A8�߀�۶��Q_�X9'!��vέdK����[B��� ���,��5�������V�;�1yS���#1uXwg�o��� ��4j�RA�K*�N���a��-\ �,��*|�L�|�Y��X3�_H<�k;#t�o5��/(��dG�+���8����@C�e�V�ߙO�J��`#8��A��d�Ql��io�Z�BW�~�fīwH�3~G���w����A�cD�/���៍B2�2s#�W��7���(�&aX��!<d28q����B�^O*�!�m��g��)�4� �x�ǝ�F�1~�؎b�#F�L���8
\���^Uӝ�b���f������_U!H�����o���+1W�/����V�� �3���)�{+s�E��u����3�WG�A��l�)��*	�S�<�Oc�E��\�\�B����_��V��Ϩu�K8;i����̿W�\
�B&3n����u�n����(��U�M�r0���־j ÞR1�u`�C[ܕʥ��Љ���?����r���=���n&x���I� �5f�d�>v���E]S�(�P���OÆa���Px���}}�9�'�r���C���*�:fa��S9���C�5a���;ފ�S��7����=N�Y�M{2�TR}�8b���=�h�l�lDs�G�(�(�v��ǥ7��=My�Ox��*QZ�]�q��0�MZ�r�)a��s�s!�f@ϒ����b/n\����q�1l�d��_/�v����16�գD�uV�p^�fѩ�N�B�L{p�h7��v�7�*���oc ����yQ�aJ��q	ߎ=�F��#E~!٘��^�������s�d�y�f�";#��U��]ʡ�5X@������d2������F��9UPM6�F_��>�85����h��u�o��bP0�x��7׀�#��?��B[c��%\C���n.��l�e.� ��l`�M�w�����,h�á��4��#��{��ұ��ԧ�Z���ЭE�{��}��eg�'���-��Lv�-E���g�^��jq�e�]$q���79�K7��Cj����e����z��/sxT}{�.7�:�-����0�rN3�s�ݒPM\�c呻�a%)
�f6��<�n��S�b���29p6���+�>c,���x�Bd��!^��T��m�@�J��w�'�ɾ�ȟ$Ug��>@z��S�,-$�@� �E�[*uZ�1�yß�%S�E<�OϾ�����S�\�oo'�ȑ�>n˓��{`��ki��h	?���O����p���������d�TЯ��F)Q�i�wm:��9��������!FI
���ǻ��9��v�B�[��5ՠ>���C�٠N�ҕ���e%���㜰����'(t��+p��h��9��*�߄����}D慨lp�@��ښ��O�������;��@n���dX�?un[eɃ[Q������D��X~+�������̘�B�^r��Ǭ� �# t�������R"�)t,��{tT�>�g1���������^I<6��rl�Ǽ�
?�Usr�c�'<��R�C���G W�b9�1�Sab) )�[��JsPUj�3w����;R�Ӌ�d ��p	4��W���Z�v
��]��A�:g�($��@�5W�R�5P�m��:�R8����ȇN�?����zS���O9�/G������i�e��k�c�ه�����&S0O�0�&�'i~�0�(�\ֳx�� ���x���A�^��䃦�>��	zw��������Z����z�԰�9��[��T#|;�=:c�����xf��V��w�E�4y1��S�\���^�� �0�B\�^��pbM�|˅g�@/:Ny�W$D�>��WYH�-�����	���Xd@��]���r�ǙN;�iE��:lь�.wCDO(����˫��[�����t�ѵ/��GL�������o���{���yk1&a�tD�[
N
HF��O��nXzi*�����S�ڌ�F�sզ��|��������M���������H'H�<T׷�0��6�ԇܺ�I[ap�cB�>����y��1����ٲ��$��2������$��NI�,4u2_���F7�#�:1L��BY��oW�G����P�i� �(�-Z&0��K ��ހ22��3S��}[P�(��u�Ox���~�:X�B�M����$�J�����BX���6I��ܯN
��F6�E�ϨM��uCʵ�&��}�;7�r8:
k�#�s�i1n"�̛�gՃ��ͷ�
�$��Y"Zڶ��,�S)��cU�x��r�s#�mm=��v�%�c��`�c�jOн��,w2�gc%޼�7(P&�c�z�����~���B�B2-H�Ѩ��?\q'�x�2�
��r��ue����T�[�0X��8��ǰ�����ҺA�߉�v&#�L��S���j�C�zK����_� z�ꉵJ2\�����tgf�p����i/LT�a����yi�C���<�D+�\A����F	!z/>l��5:Ǝ�`�Q{H�ك#T�ΈҨ;�U�[A�uO'j�}X5A��yx��� �^ᤸ I�^�pT8�l�w3�Ń#I�w�.L*]US��}��vL�1���#ߛ��+m���3E���@z�"*v�vPj��i_&��������h|���q0+2t��5qmkZH�;5���_��La��hG�F�&�[�q	?�ZM�܃+�'�&pjoB���[Umz'�5Ο��:���VZ�M��5�k�O0nҘ���`�Z�"^�R�l��7�*���Ȉ��M�'|T��Գt����EgC��%�@�;��D��D�Q֥���Q���+�N7D@�#{�x�jZo8O����C�.B�����ϗ�������0��}�Ӻ��G�w�٘I��7�XE�2%#g��f4�B¡γ�[��B�xJK���:����z�X�Z4iŴi����ʽ�B^�ү��9��(8'�,�k���k�[� ��IXNɻ+ŤV]�m���a��eO��˵H���K�U��u��#\��٣���8��>c�2e\�]�G(l��N�X@���C��bcM�����_�<$e�&H<�ww5R1��O�kE��TK��*�`A��|l�Awqs.<?�/)}���5H�ՙ�M�5��g�e���v F)�2�z�`�2�<~�8�w��5�N���/�,�iǼ��A!;q�����rϛh��v�7,�Q8;ҿr�x�e{��{e[nB����N�s��N�jdi�v��F0c+D0c-Vs�|,�$����%��e� ���k���ǖ��=r�8�(a[��)&��]�YAJ�3�����s���CX厈&��B�j*n��QZ��m��@hϜ~Z|�QT�Us���~)���I`5wjׄ��>�t�s=L����r`�	˃�&@ƽenpF��ւj���̀�֢���l��]a�[��d�œ��[�#�9Ɯ�D{����ƽ���h�x�)�W�����N��֪w� ]�q�3!H7y'�̊�M�ޖ޶��KF���+~�G���XR5��Q-���[���1�\9�2h�%��AMz]�}n��x���"�3��X��o� �du�{c�A�M��ᩇޖ3k
k��:wc{�
ގ���N�3��"�L���m��fP�1i�W�y� OR:���^��;��A��4DX�k(��Y[��@�W�_���W4�>�����UeU3+5��ո�'��K���>"�;�8=L�up���j���Sδ�]v�4��q	�j����e]F8���M&�
����q�L��\��χ��>���N,{P�1��l�	�h0�gyHʟRUM�x��n�4��=�\�M��$�\�%atd,5&�yڋ]e!�>?	)-�RʦO�DD2�˓�|m��7�K{>���»�wp<@�q⋈�����0|�%Y��ib;��ޣ��������m��x4��D-UT9�1ʓ���*��N�j�4�����P�!s"�A�^����s�̢��Gwmb�����{���b�ى�p�d�X}^He��O�c����.rT�#ٗ΄��lU��A���nSU�{�{���	ڃ��D(q}�/��]Q$BL�;fe:��I1�)�yE�hL�\(A��b�]���
-�W����l ���4EO���	�֐��<7y�'�K4���s8�\�r�RYƳP0�)TQȄ�w���2��C�g��]u��t���~�i.\D����\l�_�lK?�����f�`P([y��j�'�6�&5\�,C��
����=3/k^�}��ŧ�8"�3�!H�-���2~��W������^�UR�%@R�yk�c	�P�bm�~���9u{BdB�9�J~��������͘���,RQ��X����:���Z(>yo"F���5}��MG\%�Ͱ��T��u�"q�	�����]�y~��z�����~30�_D�����I 4��䅤4����-��u�._�f9����Me��]A��9-�*��!�UW���̏���xFZϣ�A���a7���O��i�A��!@!V���noGzFW��ۤj-���3���{��`a�i��7j��� ����&�/ ٕfW{�7���1_�p㔯*W��H�Pg,|q��G�.ܜ[u��eU`3~��6�W%ż/��`Rx��1��Xg�����bk��[�MH��;��UUO�M�~ľ���Ra�;o]��S�j�<8U4H9'ΎH���`7���N���Q̔~Ǌ�1h�:-�M���7I���v�U�rU��t������c"3-^~�k��'U~�j��b_�>�_�N��v��A���m���ZXEEP�������֚h�x��&��sdxr���]m��XA�M��n�~������\��Q ���3�Y�O��k�?Va!���4�ŊWQ��(�W���=��K���Հ�r��*�1��F�0������-�܊X������yn���Ϻؙ3,��޵�ל�ae���'r�>/
0�n��.�Òwp�zۥY��QG�h�/n�9~z�hR�S&��)��;e��8�k�۞�8n(GwoqHRc�A�~��B����w��Y���K�{�0�Ns���	(��?�]R=�ԧ��)V��rq-�����+��2��RQ߲�b�h,��ª�z`iG�[�m�~ �>��4��`��+��e����@;wͮ8�r&q
���7� ���X.ݼ]ߪO����z��O=��i���>��,�o`���������N�u��F���~���a���}=f8��h��[_"���7���2�Sp�8C���\iuqP���9��1I'��/����#x��M�O�|~:~J�fX��Fz����u7-���<<x�2y����e���b��cNc<�9�x2	2�w�6��6��\��X��b��|�X'Y�G��{<�:��F�_n�Ǟ/�~Ɩ�'J��1�Է��E��hA.�T
���~�a���U!b�!^�!^xC�+��AO���ٽ��*�h-�o�aîT�G����	�I�($�/�>��\!L��K�n��\��O��&�b��|�-�
�"���<
����s� �a�־l(�L}�MVL }4�X*5� 뢒��(�
'�n,��L�� <Q�S�i9��y��a�Ő� 2��ٌ�%�X����x��Y�w���*	�58kC�Z�q��s�0�X+z�7����\@KR�?�BQ��1��g~�](9t����cd�G�O;0��c��+2R��Tv*��v:�"�&��˩�4h�lx)���wSP���ɲ���<WfLز�'�*��	l}�t��������|8�zX3�)m��e1��F��T3�2��A����4��-�mKV桬��zu�ǋ����4]T���.���O麵� �YFh�\!/u~�����m��+�)��&�5�<�bO~��&���O	����:4��ҹ�!�q?���� �9��xh�d��=x&1Z���kh�	���Ǣ�k[�-��,�jd��>9N�@uז���(�bj��6ZYM��B���#�e	�(�ځ����5�y� O�q=�ADnJD̗�Ɓ�/W(c��[����N�4҈.��T����7I*��_�]�i�W���x��K|�u�4��q��T����u�Ȥ�)�e3�㝗A�3[�1��fjf��A��JoR-_�?$N'>��e3L3�:$��%���9�|�ߞ�K�3�)�NrG���Q��.��x86�u�f�-�`�Zփ�#Ր;��J`���/�7ɎcO:V)��⢦�],s���@��.�b�'*�&=ɤ�~&/�ۓH�ys�(v���ػ�j�2��� ��|#��0�����f�4\#���*�HV}�16��s2����8���;�o25��Lz�)�˗t�%<�3�h�6��"�i���gdLW~W�RGf�lihP30)���1�^�	�i.ݸ��@��T����6�?ǽ\��!W�P�4�{j ��U��X���0��9�K÷����a��,�F��물�1����E�H�rv�����~��]mLbN0�%ya)�}�<��FJ/\�{2.�GHp�,	��vA~P��1�{m
��Ц�����H�)��Z(�?_y��S�ArD�����=oo6q�F-�c�Z����/ߪ����}Y�*���>Y��*q6U"t'�^��0�}��ư��
t��n�Fa�;3]�JP���"��XA��b@��,d������n�W�GS�l*�0���MFw�e��p�q�xO�M���7��PXlJX3�PK�0&��@*)�'��uO_���}]۞�e}Ɛ��(~���������B���[^@,�4U��h�nF�W�b	��i����Ȃ�΅�sT��`E�c�51:��ɧ �5"�ilZ��>!�ù
�Y��ɞ}��n/-�5�^x��5�R� +m6��D�/`��G
�/-ܩ����.̡D���ˍ�Bn�B�m5R�N��mW������y�B�aT������k�G��|�'[1�9q��:C�0`�z~:L�n<h�t+$֐�`uMb�Y^��S�j�~��["�mc��#i��<��"r�,���}�<�6q��,���n�B!�>��h^M�Ol��<3�9�@g�1��#�] Z��r*����z	^���!�L"�n�ң��g�����z�1,+T�ݰ����䧣��A��l��PJ
a0OWh����CI�E0���v�Hecw�����6p|� h%�M�6S0|���Ò�)N��U�\O(���bR�@`��p��cN@|t�]�L���M��t�r��b�3�u���"�Q�`��J�J��+fv�ќVr(ʧ�m�Mi�
��e����f �ݨ�$�b�U�ekx���,�⺝�>1�,�1��m���|�w��݈�6���u��EB����^4�P?ƅJ�f�h},�b/1j���]��(N�"�"e�,>AP�]��e艤��x�/�O����Y������_ �I\Q�1�����;P~��{��@��2p9}���h�XU_��~T�����F-��US��ゼ�����͔���QQ�ieppċ<ӳ��Ɛ��wŕ��Ӝ���Y2O^����Qp�g��2'	]�Z0�qORF�#�&��ZE]�t	��S�[��n؀|r��;�8���NR���"! (�=Hn%��=��V���:����Rmmd�\.��HK�\���w���a���g�7��/�����
tK~�м��$]�
�{v	Q���v*�V_^�.�Oo����Y�JqPR�Қ�PLVD�z��� �N�%��8�W�O7a �K��baa̕��iigB�F�ŇZ�F-/���Ġ���y�������n�Y1�����0~C���=��9�̅pk
v�Ҕ�b�d�j(�؛�ZN`J����zy7/�r���a���ne�^���0�Q�%�i1!dB0�E�qL�G���]?��Q�?"���࿏�c���s	��m����5AM�,��M�ݤՕ�T�ښ������A��
����^xy��?-�	�8��;�r��k�6�VTs�=tf�Z��KY����&��8�2?�����V?��M���ֈ��L�byB�+ 5��R�g�{�dk?-��`�����^���})|���j���r7 Ad�<C�l;Q�"�@�{ي��bxd��Y(-i�L�:�_+������,�r%��ioń=���� 7��i�N�;7��+`���k��b�\�D?xzjYM�%^��gV�!<R�?����;;.��o���0b�
)�v�րx���fv~dZ���1��ݨB��Y��Y���:]�
+�<b`��j������*��.2���Q��e�f�͉��dm����p������BEGJ�al��oQ���A�K�����DWː8$C3]�ʩF�wџ=�� �Y����b)B�F�wc�X�����dca�S�˺�������:&���3��K��t���(Z��2�	��[��WjW�B2�{�bI$&��?ug�ñ��]���!܆=p�c�ȟP$|���s2f��M����#���P6(��$���%$De|��(dX���S.�e�cw��
�#<�#����A�K��J%�mEs�f5}��2{�ƹ�`Sx�M��;p����1���|�X�m#ՉN�<�\�w�����Tzϲ;�[DG�9�Jq��A��ǰ!]&�^�63��i�S�) �	g*.������L{���?ӓ_�3:��$	��_2�!���r}�z^�(8ocEA�<��R�n�  ]�+���de��ڏ�W���Y=r/�<��������(f��tR$,� �΂R��H��]2�9��疅���f�/���9�AJM�@���e���
��銺��z���޼"TcAy4r��KC�K�]u?9�qy�}�?��-�����,H��o��!��x��� ��#��՛���%r���%R@�+�d-�~��vz���2}�2*bt�"�$�PkO�Җ�::ygp�:��&�20Q�yDm����!��T`���X���\�L�p�I�������s��E�W�z?<Àa'*.}�h^��h�(�kM�H�4v�X�^��X��W*w��*j:���슥%O����p��OSf��/�U(;�Ь���᭓�J��ܨ��y����X�	�J�1�{�����AN�@��K7�;=��m�U���U��bw�ƙqa��#�+���g��!JvY�Y�&4��K9T���[`�k��C���˺���yÞ�]� �j�_9;'��Vd75l��2��X��?G�w?K	���sd�=>����
�u]�N�����43',�@�u�*���:c�4]���K���AAr��o�;�R׻�~�f��շӻm3NU���]������ ��v*�\n���P�F_�(�x��+��M��i%̱`�b�(r����Yc&~�JF�c Q���f���w��g�#��)��g�'�jwU&BQ�Q���U&7@P�v@����ͲǨʇ�~_�*��-ɯ��"�/񻡌��O@:�;�h��CK�iU�?6�LEջ��\�]W�aQ䠺����6���.���Q�S�fЌr�kz$SC�!���(V¸k_l{�]ܫ�=7hJ�a���Sl~3�5�!���h�
�𗬎�%��C�C�L�#�J��D�cnص��ud�����*�^�^���w�V�:�j�5���P�'�>|��v]U�Q_Ͱ�D�(�ى'R�ԱY�W��N����1�²
�Jm"�h�`@x��CR�<}os!����>����Myin�*j�T73kt�!���'}'�)2��0q�d�_{'��UMz '��e�,ԯ�"!�D�vI���ȍ�5��T�m.�+�������I���=�|Ȗ��S�8e^�\	����rN�*X2C���N�B�y�#URH�|�1.e�џ&��D����hnd����MgMH���^<�'{�e��ё�M��tlN��eB�x+nFZ#�?��f��h�����V�}l��_(��3�Y�`W0Q��$R�;��d^$�漈��6�t7��������_�Ρ���MlL�A-븸�ۣW�>.��Z����xD6���qjp�jC��.����.���K���B$��Z�h-_\8� �9`c��Ц
j�+ul�3��1q/��®����da`ێ����Jˈ��U��U�\���K#��mhXp<��������r��љ�taC���2y�(��2!��3��x;�*������R�}u^Bl�(�2R�� +��5SJ�k摕Hƛ�����%�֧��LY~_�+L� v�%���}(�Ȫ�Om�!�2޲Y�H^x�wB��E��i:l�����6ZS7w�ts��#^���w��������V;,�T�Ԏ'�/��0IQ!R�B�ƒں�ֹ�"���3�>h�:_r�r���6�>�NFL7�5HK��)04�Ͽ��J�rmѯj��n��"b��<Ldg�F��s/~]h"Ʌ�\���]�|2�'���*��I(�>������LD��Cǜ
�ħ#(�\Լ�!�i���[�����=C��k�t�P�#�Q�L���:��9�'_*���H��qG�k-��PB�ץ���ȌD�e&�u���M�rĈ�=�1���4QAӕ�p����~0�P	���'+��D�S.bE�lS9h5��*�� �����'�`8�۬"���v>�(�3_d#q�E{���=�|��D֫٤��j�/I�����-�:��˙�Y٦�r
Ǝ�v��y;i*8|�P��vEf:�tgZYe�|zAB�L������F@p����ёC��G��1Fn&a0�Ð|��bzO�c�L"qx��.H Pw	{O	8�ьT!��x��Z���$��٬�ėW#Qg�n��=��T&ܳ?H���b���qM9Z��7E}��^��Di5�"�D��r�����]嶂
���g�|#�Y����3ҍ��@�_�),5``�r8�	�Zd�����L�Mɯ���+ln�l���9��fr����L����tb�Sz���)+#/�-=��`����{��i����!C�5����Z�OS`��DHʡ���ñ�@9C�i���A�1긋�#��n?��F���:`1��|
Qzl���J��v��,.�*����T��߳����K��q3�T;�JYUԞiVa
�&����&^p�sUU�Z�>�Vj�d��l�( U�D�5��?RI��b�c8'A7udm� 6�!L���?F��a����j�52��6}�b��p��ۅ�]�k�-����O8��d�TƺC���jw�(xǄ��mFb�:����( ̈�*y�|P�K�5)6Ơd���A~|*�D�?"��$U5L,`'v�[��%��*���ޙ�-��;LRPЯIJ��NGDP���R�~�%���.�o@�@<��u[�:��x���Ƴ6ޠ�[�,=�z�̹+��
�8�鳩w�plB�
d�����/�P�܌#-$�Ej�,�3��ש[��
��� �F��-�@&�	��l��kLV�nd�N��WI�?6�
����=s`e�d���*��m}/�J��i�h0l�Σ�tx����&�okP^�أ�� vh	8(
�22F���"�X�V(+��н���(�댑p��_�M�	��>I^� �R�X��7�&c��f,����V�!]�
�������3��� QPl���鞋�ʖ�>��X������n�_��g!~�,���,�؋֢��&6]+vZ���9_B d��x����h��'xF����G:1��R�i�/�5pX�.������m���-��������C:��U�x�<�&�?!?`O�q@�qfG����{�zɿ�Τ@g��`�m�ֳyu[�XҙD��� K���x�GU�������Z��"'��?mb�{�]5�y�vo��ۀ�5D����h�rY�@A�=z��Wg��#y�U���+;2;�@�.���C�.Ni�C�����ˡ5r�Nnm:n��ݞGnBg������֌�`�Z�9�Å��b?���u�p�� �\C�,�[ʕ,v�p6�1Q��A��/�ge9O����6��Ǆ{��3��T+������9��Ɗ"8jˑ�[�]��K�3�B����� |��u�$����]1���r_�r�)�0�M�W��r@ﶷl|�6�5n*��Ѽ^�ռ���o�0�4KHQHї7�p�
�`�S�V�g��F��7>�;k~��J�o���_$����{9(�A� �%1%n�E=�#�i�m#�[<��:?�l��T�zYh������a��n��,�Y��"��T�Z~�⡴�mGQ6����,�U�dp�Wɥմ,���4@��~	����7XI�IaP�H�E���>�i9�qa=����U������j�e����l�/&�x��I��P��jt�P�}��ٓ{�׵ '�y�P�&�U%]��-S��4��Ȝ��L�#��+�r$q_�4>O�!H(��.�y��w!:���3;�D�:\�|���6п?�K�OdSPu'B�*�P�u��K��E��P`��k*x��hJ:i'Z��T�=S V��kG�>M'�M�%!TO���|y���S<�r��)$�6
�����=Vp�b��Ա
�t�������3��/	��L8D̮#"*�21�JBؕ��B*J�k4��� �ɀ"o`;X��[Y���G�dm�D!��S�Kb��'P�g���4�!ڊ��d6D�$��i��'����u���H�5�3�ܯ;�6�6ǲ�^��\�����T�����B��)�:>)O`�K���o)B��B�����8�d�n7gJ[zƻOJ��9���OX}��qAJ�=<�/��s��xԗߢR��y��a�`d������L��oR� ݎ(Ĉ�L*1�\�aI�m�1�r�~[YE�B�R!�)xz\����O;˯�������=�lj(j2��vk3���|�I�Cݖ�d�� L��L��:b�d�43\}l�]T:��p
Yd7���w�ͺ0F�,�e]�&�UVT3i翁O���ɮ7��H����*��I�K��Ot� L�Va�p��	ԏ�80�)9"����������v��Fa�Y�U��g�� [�+ʽt�gb�6����w��$T���{��C{��Ґ�����y<�.J��<�=�}^�@�٠*�jSl�Z�Wc[��^ï�����J���k�Ƭ�����!� 2<0��Q���<��6��!ف!� O�햒
vI�E=�=c۰ПNJ޽E�BK�%.vN�?9�zkܩ�p+�� �<4nm��ʔ&�N�?z5s�r�˺'��>ܮ�P�`v/�2Q�3@��p�1u�F�D�#�Zr~F Qujc����}���׍��e<���++i����[}|�5C��-���E�FɵPx��s� ���4�ɫfd�E���Ud�c��lDN�DH��~�1N�N��Cr�f�w��f=�~Q���2���)���9�h�?�)��o14�)��5�搹#�n�&���}�kUO� ���	Y���Y�o�[�{/��N�(�\O0FG��������`o�> �
s��L��{��9KhO����m!AK�r%�B�b,L�"�Xr4/m�g*����I�6j��u��=%>��;���J�Xm-�}��.�ta%A��$T�3�_߷YIb�-	McO�=�xl�q�a'�l2co){�^�/�p�KWg�X�#�p�@͖~f�q^ϛ3����[�~*$�t�U���$:�P�0��m��Hqzx��y�#���y�J$�K���I|oYѳY���T��ԉC���^�Y֞�^t^����[_���჉>�!� ��@�j��(HV-h�@�0?�4^�:t��<����J8�����'���,��N��2� ӱ�b��_u��>eB
����7�-�h��!a���-��DG�~�J���G�Q'�$�E����s���Ɖ�<N{��PϦd�;nP��WNM�1��A�"�������g�%!���W�-���%�2��|�'I����#J:�}�i)��&9sm�x�91�����	^��O�F��=X	pQ���C�R'�"�����C>�۟�U���L��4�Ӱ���v$��8��E��5Q��H�������şy���Gɜ�^�.i	g�x �N�U�**�LC�'�����#�<~��@�[c��	K�c
����٧�U���6&���vw]�:�x9y��</���Vw��ǧ'	}�7R5��X�*�9s�(�yV;7V.�^��� #nmW����Y�~u�����h$�J�M~�J�e���hA c'i�p�T�珯b�;m��[L&9 c�^�2�N����mbf�!�
#D�&��Hm ��Kg� T�ާT��7C�_��`]�;]<=��z
7�y�i�8�Z���i�P�)"Ze-�D*���]���Gn�����Ic&C�r/���]���|d��ƾ�\�A sfO�?ֳ�8���϶63���R�8�����f��y9�H�T�lF��FK���@4F� �]eƺ$!�� ?24�x�b�V��π�����f���U�7q��hS;�"�!�D�r{��Bޱ�e��b|E���'_���׶��l2/}�~ʗl��h�m-mD��-��j���~Df���})�hj��*����/��se�� �-1������<��ᓷ����Eo�c�K-/�瓎���� $T?M��"��.�*�d1�gWfْ�>����ą��yq�G����EH��!���?��3!x�d�JW�w�yğ3I!��Z/x�� �~/Bh��J�<�q�s0����1岆a]5�gk��qO��]-�BP<}�d,Q#���&�-����e�\q|��bK�������.LD�x7���-!�sIU���Q�ս��1��VZ�P`B
��=�o;AS�5������	m�%�%�qTy~:��fp v�Ԭ�RvK1F�l}����xv���Vܢ�齱8���e�]^7 O�:��>�y��d��ԧ����0��tU��,�����A$�N{�%y�>��sUM( ⼖A�6�q}�d�M72�0#�Q7�9��vHOIޟ�9d(]��!mimh�V��8E���$ٵY�b�J�[�ȃf��>r��9,���D	U'A������ئ��J����^>��]X+�I�K7��	�B
}i�-�\�<ȼw��*������Uu�Y-����LL����������WN/JrP;kגd����5M?��✒��/D��s�a@�[����^@�oh,�X���v�g�v����2H<q��~p�����w��ne6|̻��/1_IA6~O�b��M"�2e�c��is0������aێIA�<�C���n����� �(�����_�^ܤP�	ʮ6���buzW�JC{�guz撱� Ѫ:K=鈨A�H�Bp�~g�� %O�!�rv�WK���i;{�u��$�kG�|�YC;Ǧ��`8f�uB_B!�r-�<��F!Q��,|Jd)�*��T?$�f��&���ՙB��xbqc�ײ���G����Yü�.Ϲ�|���0S!�!4�ÆJ0֙qzp[����d�<�Ji×����߽�~�Ʋ�/�_�(ʱ05�D�m���׊6>f�������.t�z?��(99qĲ����K�ؓ�������Q-d���JZ�S�S��nK�}�!��`�E���@�{�՝x�'e���ń�7 ��B��B�Wgw��4X�E>�A�,�z���#�
����R>O6�,B�ܴfv��``��?���3�j�0��H	���-�$
< �KU�M�諑$T*�ч3�ѯA�^�����3����^�Z��~��1ɻv��Ku*)+�\ߍyԂL����K��ᗀ���f;S���j��;�W�TQQs��j����n�ˠǀ<���>\R!�
v�O�|��{&fF���0�+�j��E��^����Q]��I-�����g<�>�W�b�s��a�O�[�pzd��]���P�	�׹^�i9#CXF��F�#�7P�w���	���bBF1��!+����j�M^���������p,���f���Jѿ�99��u�Tի