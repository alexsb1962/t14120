��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:��������uA��@��y���<����xDET>��W�����C%�=U����3v���hj��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	{>�nP?/��[
��g%���0�r��M�6�ť4�s�M<y�Ò�����z�u�`/A���F?視���ksO����%��'N��=O�<�Ș�{b�)�g���:or�W 2�՝j7�`��^��w;@��P��C��Iv�&w��ɨNw�����.J�-�o/��$^�h�@S-knS?�-�67Ļ>��Yė��3���5pU3	���HD�?Y��Z���=���N��'w�A
�Cg�׾�pN�X��lH+�-.���VYѰB� �KHk�"�%��$C4U���?dP�>�Gf�{Y�HK�+Ԇ�qS���8<�u/'�H����V��о��Ă�v|k�~�*)�t�'sQ&��*���@�-M)JG7�358vVnB���`��)ی�%�P/��s/XzN(��vshO�"��}C١;�A�bh�j�2����*����lrE+�魂�MM����c��P����U�r���i@��}ke,�Wʘ�5��=`�q���l{������O��rcxW/M~�9d֞�w	�"��`�-�s�ԙ���`�N�*J�2D���lx2<s�=����BA������$&��%���2��J�~���p� �!��;Kf�Nb0;�v6��O;^���|P��i0���C��i�*�]n�9�j�J ��~Ԕ��lm�b�4�����U.��	.�|А�m:|d��7v�(��^C�w	�V�ĝ�σ% ��BIv���}�4��3�ζ#vm3��)#tp�Xc27jm�y�.
� ��ޔ�����-1�E���~q��=7L�������*�b��+�Y7f���C�
S�@�?Na�& M���^�������'>5_ͬ
y
FKab�����L����ü���:ʤfS=�Q���	�Z�m���	����N���0�t�`A�t�g@���!!��(e��|�ӌ�,��)�o/������Z��ju(~��MǗ���^� ǲ�xe�`�S-�S�g�`f�	.�����w,�"�^�WqD_�m	�(4���)��ʼ2�RJ^��T��C�4t�Jn2�����QV�|̗gXE�.����&�W�dQ%6�֔...��$=��Xe�r~�󳙽swxN�����(��NBk,�,�<��T�֓P����M��n��Bx?h,g�,{!����E�g,�kM�|lh��+�q�stv�{��ח��YkTV�{�[k��)� @������@:I�t6��i�gh)ٸf:.Hx���q,�20���R����}���N���j9��B��������V�Z��1�3��=|������R�.z?ޘMp ]�<`��v�cfwd%}MAjE�P���4���%"�F"1&:ʤ ��f��C�7��36uy��В")M�TY�|ely��@�ML�,S����T��O,-%vmv��yY�X�2�kt���RV�@ �h��)������)���/�?�#E׏�p.Wc�Q��8�VY�{«b��ݝ-o�6T���ґ��摣'%5W�s��Y��*��M���G�F�����uO���x)�����H��7�VGt��c��= ��߭�7���%���"TCc�Nv�r�\��`�3���m't�A8Nt�n+.����fO9� =:l_<���y��ӣ.�NXݵ=Y"ǃ��L"-���PC���0
k*�~Y������!� -�N)+���{�����]R��7n�
d���>Y�&��;[ ��2����$G�^cH&�i�1�6�K�c��NA���	�NN%����k%	�)��T�����K&�b�l	êڴC�c�7���&e7�ɀ�~5�eV�-Pg���c98���F����n�Å��F��ps�g�C��X��c�\0{
3S�C9���C�f*h|9�ϡ�^��
������G��@��`�R��Q��&]��&^�j� ��\���i��|4#�hrОS !�E�-�s��}�����u&�Hƨ^Q;������I���������ηZ��}}cN�J#�����v zɓ
��$X��F�L��,עn�긢d��&sOʲH�aD��&��<t�_����0� ��2�����=D�Ҿ�oT��8�gK���'�9���� �ϧ/mwY+�G��,Q���r"g���V��G!�Y= �Y^��e���EK�ͮ������b�9\���]Z~O]T�f�'�!u7�u�-���ל�B̬%�y�O19����=1C�?Ն%-�%
����}8��TOב����M?��\t�<7��4�W��o��@�O}:��+�	�b��˜>�ɀh7�z=A��׭'��˶�1��븓uju.� 6���ś� S)}VbwF���o���ެ<�ͨ��q)�f�`�>\=��$N�=@,�<5%//�ݮN=ռ>�6�<�ͺ��������ݥ�>]gZ�0�z�Z'T����U�L�r�|� ��x�Y�QA�L��2�:�27����Eu����0%/W�����vQ��$��f<>�{� {�C�fz��C�Zxs#0#ˌ�-N��ʳl���Q��v��M~�GϨ�����¾х�t��bE_	�ϻf�&��{��q�Ӝv��Z���f+_���V�����A��н��9���z7�W@�si���Wuƃg���������u�?�(��`�Q�o#%AU�:M�NQ����X}cG�iS<�d[P���T�L7m��h���G8�I���ax�ZO`nH��V����G�zt8�?U�=����,֏�x$�� ��\vz��	vz��@�h�2���=kgM�-��~��*�`=�:�*f��Ә��?V9D��(�M�7���w�~V�%��.�Q����L��M�"V/2)b���e~��n�/�&�'�E��?^�c�1��)+2\BHjo\��v��?�7�Y܍4�NcU�����%{�I��t���������MR��D�}D|~�g�1��Sii�S���s������7��AS��"uyIJ�cύ��
��]�9�f@�1pR~s��#x�;F�į�yIj9G�!'���OyKV@���,�4�{	��̾��c��`S_�G�0�*�DV�t?�_��r(z�G�$����M���d�F�t<gmy�Hw\&
�M�6k��YT�.Qf�!�~�������Tk7��p)�&ic��p��o�%C[�g�UQp�7Ȝ�c�DC4�7pv���z�i�MN�k���roՖN�����Bl�ٮ��!����k��=��C7C�g��x7
�U�}���mƿs瓘P�l���E/�\F���h�% �3���=��_�B
���N1?떊��#����yZ�\v5�p�?_��v�����󤋼D��9�)W$�~����O�d:�o;-�۳�6�9<jH��1b���h��H퉤m�0�C-E-�ة�0��i)�K|�վ
�@�t��D,9���{~%�	P@s]�]�Rk���^�峾qUb¡�8&���D(��u,)f�}uʹi�*)խ�3fת����SH>*�B��2%2��6R�q�ΝG�̈_����*U��W�6,9�!�UU]�le��V��K��a�H4����}���#n(�ڣ�P�;.�"�Z[����D��
����w�'�S�o���J��q���8�C��[u�Ak��J�*��f�*��9AW��c�;ܑ��B ����U�vL�����l�{A�4!U~Z�&��n1eHM4��R���`����LiK++��K�?��H�� ���A��п9���_��qZ��햜����D���t�0 �*<�*Ds�\�`�H��$� #\�^^2,l�M�̂���|��<#I*Sˠ@��,��o쬖�$�~b���$/�g>h�d�=>|.}o����N�(,S�Z�E�~�ۈVy�4"��ڷ��5H����P��#����<
���[�?��Z�J��DKA�R��)�|��qSR���09I_]�v\�>��������=�<�2n޵H�LO/���F+%�V�27����$#��9�N��U?��#�CsQa����w
t%6N�4�p��G�@�9s�@�N��Etg�{e6�АY׭�ϱ�ߚo>�AIm�O��Ke�4O��������GL3?�F�	�g�6R8pC���ٝ��W7���w��2iP��?��E��1h��rpL;f�cg��A̋�L��"GW��Ҥ����K������S�
�Z�3co�Qr��,+hB�8Y�:O�Y$9��-:A`|��F����&A���^ۺ�9y��ڱ�b������22{�(�����|�����L4�Y{v^"\���'�G$�P�*�5�3&�)^�%�Q?d�-�;Y"�r0E���ޕ;/��ֺ�Y�zH'�� ,�ަ����KF���{(�t�5F#�������J���<\����kM��n4)w�O2�9��4��u_�p ��f3>>b	�E�LJg��� r�[���-��w�1ӑ<�/n~�Z��O�]/,��IP(��:һ��AFZ`x�9�dA���&C�D���y�o�`n	1��U5NB�ZᵤȣƗ{�[+�4�]�QP����è��E�Ń��E������R�m�~�-y���+�Cѹ��B�>�UőN
�"8m�b	��6�E�������e�@�W��u�7��H!c�:m	�iO�7�8��+��h8��T�� ;z5�-�R���:+�c/��VQ���ʪ����{/<��Ŋ<�1�C	aq-'*Psd���9H�t�N=@|�z,m>Y"����HC��^��ʓ���i�rή�="X�n����[7�yN3�(�&/���n��h����hK@�FSb�!)Qߝ2���8I��������51��ܲ�b�*#�S��M�),�9ŗ��&ǘH�SG�V�H6��^��w$��j�Te``l7㒴�T���~/E���m�_@C&9U��!ؕ�p��yd6�����fPY�p�q���kﴵ�t1a&$�]���ʊ�\�VeP�F?.�� ����pv�b(LO������B�r >c�%1��"30�g��_I���������3R_k3���q�r��9�m�č�!����ko�*�'q�W�f�Fͧ��"��k����}�{�"�6�F�Q��v��|
wt1�̭�4�MW<�1#�%��3���P��I8YB��`YZ�R�	æ8䕕.�qӗ�N����բS;ϷP��=������$��6����-T���PR�֚���^����o�|�,R���Sr~XO��%xk�ke�["V7`^�����F���K�B�H"v�/��;�qّg|H��=��wUF*���*�O��Z��.�쟡��ZON�e��	aۭv��l�D<���|I��2	���*�56�����)es�I�< �ͅ������o�Z>�r�4��(&D	�{˘���]=��,��e�:HRu��?����Mh۷�m;1j�i�R5�x�^a$ -�����,��COx�il����{�eWٷ��!c>Ʒ9laeO�c�Xc���5S�=y�9b�Y��ѐ�7T2ݲ�R�n�6k���3F%�9VsKջ�V_��W����?%��Y���wF�8����鬱e�Q�,yӡT�Ás{���#�������B�q�����N�o��$K<&��!,���Oip{�����J:)[�cJ��n������+�4�i �Wy��?Y���nG2b����S} �0z6�w(D���g��V2�h��r��+�,ІJ=�����4��sE8�dRI�����t6y��bٰE��B�ou�,/Xb3M��G3*����d)��eB����V�
���DS/OY�ǹ�)�/@�$���5�Yz�L�1�ԧ�.�8V��l�i�:���j�϶�S�E`�����X ߧ�����a����@
���.�Bp�Jjj��e�wgE$t"דl�� >����0 <�q/��=T���A����{�:V"�&�{�~֡h��u;������H���&��ė3�E`i8P�B_��A���A-_��"�t��� fy�{L(�gជd��o7g��#=\�D�L�MJ�C꒺/����
C��4]���o��_(3U�4 t���<kQT'��g��dp��t�#��MgU�yPu���n3U�\~���}b��e\���wx� �i\o=�$'�ɀ#��ނnIJ5��q�x��c6�)�'ZFa�]
.|:�&��Y<�ΰ��+VV�3��7�R-�wη%$��4A7S�Я^��a�CE�����o#���G�Miʨ�z�����t��,�}��7��3�D���M��%cʟ5�1 іh�"TZ�\
0	$�󥨨8�җ�?"�ɦ.فX凵5��U%�v�������8p�=֕*�蠯�F�&l7��:n�����/�M�v�4�)����wk6��R#`�G#F��@۾��w17���!J��1r��6_I
���Xl�T�$���Ƃ�Z�Y*<PAM'�@X3�!QG�<_)T<�A�L��2{�H�ݾ�)�ԟu����]�����+ĉ�t&�/?�?����xp�l~*����Jb��*O��^'c��|�{_�|Z	N�L��?g\ �e���cε9��(�������i��R��x\Km�:�%Ō��r<�}�{%��?�hUA��a܍7(
U_��6A:A:k ¹����#ӭ�$��Uc��b�Q��G����M�uy񾋣8��d�B^�����}�z���s�<'T-ʫgn�n\���뵂&z֓�mk�tR��J&r}��*���G�5��h2�5ijG�#�������U��R��VH�G3�\�uŞ�rYX� .�[U冨6�?ئ�{�퇪�p!�ZZ0��4ב��(�����zB��b�&|~�H�ǵ�6"㫾���6�;d��ʻ��k'D�r�� �^,-��b�^!��Z��7ɏ�w	ueMc��#S��.��fS1�F��e�B�j���[+���m�F��)���ƚ?���k䨄?����bU-��A(Y�Q�ǐCy�����?��D��$�EiZ8�	�"F�ڜ��rH#P's4ާ�y:���(�MX�)[L�T��'l�[��`@@�.M��W����Z Xڄ_g5vց(�)M
�E�բ�8P.�4��������F���~�o��i��"Aʱ?��Y���o1�§T&�߳ymt�Y��\1<nr->cq����0Y?�A�	,��<jW�ܥ��!\�#2k�v��8185�8�FL@h#q�����+�[���MX'�� ���H �2��U��pf�c�.P�����qZ�\q���(%���MK�t��?�ʅeY>Zw��ӹ��F��>SF��z}�qL��W�`"��^8�j� ��c
~T����Ԟ��_xԋ��&����,�2�'o�k���0�����Np�w��Y�/��}e�)Cm��y��c�o��@����um.����P��X
���̉�dj�i��,!S�a���?�0��n����2�(<�2-������1���x����:&�a�9e;S��m&J���gL�%'�e-"}�E�H�d�Yd������,$��3ٺr�e�E�������)*B6tz�TѬs�R��%��~�L���f��(��C�/r3�ɳ��?H<���k,��U	�:^�ot�{�˷iO�]D����P�! �4>R��@��dp�O@/w�6|>"W|�a3ۂ��� �T�v?�}�DX�-�T����-1r�o�Ԟ��g�K�VI��d*<=�o�UUVb�g�l�f=`KR[H�6��o��U�ω�����_:�*��؟�w�Wޙ���{�pZ�*T���ymj|o8�N�u#��ޅ�ڤ��i��<�cnmn�d�[��V,#_�u�bV����2,�&
>_l�\�}�V�wOrVv�������++�.���٣��9���V6gMG!d4���6�LLB���� I��-��0�!��aN�`��;��b]�֗�6�amJȨxs	T�r���X�g��K*2R"45���q�?ϥ�g9z����λ�����r��I�o��̶3�C.1G����h���NÉ��e�JZ��R��d>������B,¾������1y@6�r��Z����}�����:�8 �� �TŰ�M#'e�#�$S�,�E�kjm�����:.2��)]�Բ*Q�Mq�� ��c��j��F{�-�7����;ٸ��) �X:�"���N;�������
�lD�8���<�a��.��<�"�+	9�,���V�(��+��Mt�ʘ��t��|A�Y�A�fL��/A�FC?\`��W^�M~%6U���0m3�{��r��E�7�i�Y�.&f�:0�5���S�#�� @��IA�Q������nF0�	~i�E�A��`�iʌ�����T%�DXfY�Ux\�x�a	��w�<�Oo��y��f��[� �מ eb�[����A��Y��,譆�c�!»�ӕU�\��u�����^Q�8���xaD#9�����#�E��W�N�yY�q�z��Z=�'۷P��V+ Y������^�gN��q
�p���4Y���������:���+^����P��y%�M�4!4��^��A�d�#���r<��s�k������:!���Č2u�b��"�z�c��8��E�����/Y&[C��"�� � �W�^�e��L�AF~-w�4b���;��ٹ?����i�S���1p��<�8�8�.y�ɬ`��Y9�
��9��\y���U ��G�h��ig|�HQ��!�����N��X��t;S:��h��u��\�����l\���!�_s_<�#��4����Y�JK��9�l���Aޑ���"������:P��&!���0�$ah9<��=ɮQQ�%8�8q��2�U�=_���Hԡ���E➺��D#;����K�7�u̓f�G��2=������>��Ե�Y�K��&�7i��@��˻V8�Q�%���x�`���'o?���:I�F��c�Z�Q\��3-�����ʊ޳��N�J��%j��k�o��1_4��UZ�ɩ��A���"o�T�̿ϡ;fl�8ח	���!���L�w�c�?W4F�*�|ã.�A�筓�.=:B���(���S��ӅP��l�d��w��� n��Үj�a�liZ�+��3@�ά�4��}�1��<|�"?�L���'�\�ȟl�7?�-M�1Yo�_*��u8�_�LR5tT���B� 8UTdeC_��ڞX�:td���Q;�Y?������[ #ֱi�q�!?�v� �H��+�i��
s��bfd��`�Ԗ��|Ƣnf�e�lY����\��w��q(0�N��-���ݦ�%x��k�z�?�g�N��!�5[��uZ$�0�Nm���j8a���o�ߡ���-,��J�~Ʌ��!����!g�\B�㟐�ŭ�ۙ�u
z�;��1���w��B�VTZ;�%Ϸ��\'�k!X,,�;G������y��� ϐs��� ����Y~����#H�b�}����ݘ4�6��=)�b?_Q�E�K���;����H��΁˼��K����@ٳh����̗�W���CvR�M�s����[Q�|��/��_TT(��%�7�ݷ�8�n먟����)��C��G����MUˠ��C`�MCOQ�\����KKQ��ӽ���%�lI�������,�Q(�e2Ƌ�"}.h\>q��������?�r�e/����45Yѥ��0o)�|���X��|�L�����	���w��q�����Q�[��B�q3�"�;�5�	l�"a��!���?(GS�x']��v�l�"�_�l�[]�%5���/>�G�~LS���}/���)p��
��O/⻱��F��s��J5MY��pR��E�d�J �W�{��v*�Q+xV���²��&T��&)���	;�^7�j3sv�Zr�+��ZP�Ik���	�� ��$��U��[��������ݲH��9?�@�C���p ��#*Z;Z�N]Q~�PáIf��r5UR���Z#l�r|Ol	"ӦN���bW�1�c�k���y}d��r��ڹ��t���4$�&�>s"�Q#��5P}�N2ɐkf�o����0�ϣn"y�q���C5`!iJ�Rޚ��j��n��)��9h�`�LcY벰��7����33�:M/��&�R�c�9p��-}�}S�7`hѴF���=��T?��/g37ڨ��e`"�n!|��i�*�i-X�<�R�Է .���0-Lؙ��g�ܕ��h:+$ o���4�~'�	j�4�>�1h�3�Q@�?�<U��V_YÅ	f��qж6#Ț,V[�{af8�7f�s�J�E<qԅ���@N� ��\��#e��4��ʗ�����y���5p�X ������������ ���9O��IT4��%���q�?}v�H���ňt�Id�9	A��,�g���l�,��R]��,���أ�y�sУ��'�Ҽ�R~�d�7`;�M�vG��f����6S�r �[W�UZ�[Pf*��ݓ�'�Ĝ>�-5��L�<G�K����T���䂻	�E�έ0�u�	C�`d�Ġ�.�0��((3b�@l���k���:�f�]��լ?���'�K��n���n*�z����r>E,�Z�dR�� �����I��#L�-��.��s6�8���ҹ�V O-?��?]X��M����9�����Q��
錁��Ne3Яo���*i�k�{�ۅ���O�,�}���Uվ�u'UXw~H��=3_,�wY����8�y#�y�m%��xi�Z��w�X��C�7��;g�҄��"	�4�c��h8m��z�SªH�첦�����"��c��'� \�KRj\a ��,��O|�[��깨6���A���R�Z#�Jji]�ޫ�2M."9M���L��{*<��l�Y>�s���W�#��]���fB&�D��e��sPг�����3�o����M CAW":m��V��o �H�t,J��%��ʓr<Ɔ%��rt�<����1���]Os�x�d�}����@�t����F-�>,% ���3��(��0�/�NIg�\Tj���uM�0:��Tp��j'@�,�7���(�p_�:����N��~�_�O��mEW�0��� ��61n�F�l�E7舖�e+E׳�x3HZC����6ʿWld	�
��v{r�C��G�y�
|��'��_l��!�9��'�����F+fX��E]�h)��l	L��-;�Jo�n$B(k����S*��/+nzt�����Ո�~��#���;V|���]q�U�q��0�^c��̔�-Q΋�TTB�(@���; ��	��k�Ϙ�-�R����-$����e��Y�^���ƅ������$��
���*�0�S/*��n���9ޒ{W[�#=��f"��.:`�!�����J0p�L�/B�W��	�2�"3�.�`x:R��MR#9�O�z�B$l�U�C��жj��K���ޣX�.}���g��G����cN�J�4�Z��N��@���䴛[����p̩�u�W����{��-HH�x?���;�K�a��Ӕ��we~<�i}�`��-��^��� 6��V�xʌ�a��c�ג��d�ER�	�h��O�O�$�L6JƳ3JU��b�ߒ��t�! ��D�,��Vʪo�����8���< �S$��E��)�-�UxI��˰��7!~�ed�w�y�F�7J�u��a�]��S����qCa���6�Wx�z�sظ���%M�_L��|�|!��{�XW���-��g7Ѣ~O ��KiĬ0aUBN�.���d�;�2M�bb���Ǧ��xQ;т�6�q'Q�{pf���F���n��i�:���sz%o=8�9L�̼ާ �b?�,t�Yxk%�Sܓ�O�����e�>�&����h�J���m�F��k����pM������Y�VtK����W��Q ���.�,�����(;�@����HTu��5:�gK�Nf%(�n�&5�O"	������I�E�cҔ��;愿v$CkY�N3U¨�`�HR��F5U��Ow�z�w��U�\4fQ6��5?�؂�\�z�P3��L�L�5v^�&|��V�z��dp>�{5���I%�t@~2@۫�����)������k���kLǂlDh����:	�l�~q�2�[ndΩI`(��6����͑ޥ�����k�?�yb��L�.����O����]��P���GPV#������7���5��Cm��
yh>�sU���U4=��@�G3����	�|��%�,�G{nb�����>��� �lb5�gL�𗶞�s�nk�|&^�t�b$E�������A.����iX�x����d��rG�]ؙ)=V�2�y!�,��Z��[����6/���� h�聬��v�h"y �a�1t�,<پ����Vne�W�vzn�EG	I����(@ko2�J�.��5|<�q��Ь��Y�WAj~��]�cS~�˙K;9�.k���ni�� EEw��%Z�{��ip�K�@<��?6%;�R�{�y��v����#��DJ������h��p�V�|	�LټTA/��J��Vza�:Z����gV����y��&���)^:z1�������c��n�����ݧ�R%�-�|�7�2�F�n"��V#V��'�1x��y
�g}�#�?�\�Xǒ��.�Y�}v��$� #@���va6��ee( �
�,��P�����;�1���gc����Z}D���xHj.�'+Q�NE��m���V�Z��������][z�c��D�Lɿ+>@�6U���՗��{��M����:L����Ld=��vwhS������G����!>ڎ�z�(x�wwU�Q�X�D�k�,�7�y��;rp�9����}},��G�Oo�<UV��nFop��&5�Ü��Nnz�lB#���]Ҽ͂�ͼ�� ���3U��!1��dX���W�����\��!���	(�'�.{�>ҋ�ԩѰ.?O��"i�	���l�nw��UڛЁg_�:E����� ht�^������v��W;�?��V7P��Iwܰ�:��)c�Kv۟�f�x���tl)28��J`Ov)��/ϞC ��H_�|����+aS	��u�0o:��fF�f'<�H7��j=�P�C��Tj�Hl�|O_��`���&��w%ib���QB�o�����nb���NgU�q/�9
��ȹ7�0QpyO0l��w,Td���gByֆǩ�ФXQF��{�>��Z��!f�p���I���(����|�㘇������|��@�����e���W���\��I�s.C�D������+�(?,�U���4L�<��Gf�+gh�Z����f}x�v��qL���F�\Y-#����{�I'�6f�n�P#IQ+���wU��*'K�g�>� ˃�wo}~�
:|l�g�J���F7�wBmȫ����_�xc]=M� �pj�g������4���v&PJ��@u!{ �`�5�ҋ�K�[�۾��`h�r6E�`��`=*�P�>Agg.0z���a��#涥��N�j
_V'^�L����1��č�z��D��>R.eP�A���\8�ԁRw��BS�B�qJ� ����D=����ϣm���`W���;�f��E=�Ǭ[$bg ��3�U�:æ��Sޚo�Ѽѝ�o��H������0���?}ܤ��U�v鑲�q6e�*�+^]��3�}�w*e��-N��v��r����N�������ɺD�Z]�~S���8�J�2���QT�f�2c>q�@�%��͚��eS%_�b�bb�:��3?ܾ���Ĉy�X3X5����%�3�7���v^��(N�G����kc�����1���T���<�zed�q�>��H�R�p��f	�'�%י���ӟyb�%=��:!���|@a<H=^5��f�k߂�[�\�����ݫ,~ōV����=YR\R����?@�O�֯����{M�(/��T-��\_�6�tX���i�CF-�@�"��7^��h�"qP�t����_�;�r�̢vҬu�G���7�����vp3�k	��6%awn�xѶ�s.�"E1�pM2�QVA��F�b�g�Yf���>	���&�Lt��v����C���̕��%��Uk'_n��uou��j&0K�0���:��Y�����NB����Xاa�g��+&uC"�3>��5�L�o7��'��X3;��A�N�3<U�Yo>[��Q�?�y�w4׃��LrǢ��܅�AzϷh���\ҟ�	o���H�Y��	Mt��0��u�L���-ܨ�q>�\�T�69�綧 �ϰ�������v��'�n�HJ�t�P	D��Gώ�'�<%�1�
��?r�2j�?*�B��s�p�?����T�,��ˎ�����s�[�+�(|D��ᑥ]���[�
'Z��M������[�ѡ,��Lm��M��XvU�:EPA"���0�~Q�O�맺H�!P�o�|�v$-��H��c('O�@�:Z�SS�;1����l�>��Y3_���i���m��G���I7QT�U?��vI����m���i���t��e<a���o�������q����W��`�ل����" ��-�� I�v�h|[$3x��Y~�w�~���kj�Ʒzv4z;q�pM�t�I���m��=���_�a�c�Q���8ֻ�g��8��b��Y@�Eq��{̤F�^��+��O׀��9��������C~�3nn�y�����Q!����6"�l�B ��>k�P3g[���b��C�;��L�G+}���:���E�!�&d�h�`-ʕ$p��3�c��]��V�9-�Q���OC.\t2�~¨!C5�|�F�r��\������th�I��+Ż>+��?�l0V`��
P����?�
B
&2S͜S��c٘C�@`��)��Ba6�>YZ���p�L[+A���f�2�6d��1:8�̔
y.��8�0ݴ;l �4�X����&���&ba�,���b+����lf�G�y�3>M��|1�����n�k��eo��+��QԐ�`�������/��-S��A��
5�6�Hd&��ό��`#��J�|-�R�+ُ��'b�����T��w��n���x������׻���/�%����E~�PL֢�͚R�d���ܷ��Y4pjs��#��P�+�@m۽���B�?0T@iZ{b�T�z�$_�G�0�U(�n/�I�k����*��s�Cl[�m�mO �����} "�f�壗`�+�`��q'BY���46�*��
u��GG�^HPbW�Æ�23��r��ۥ�7��j�#R��>�<>�p��[�/<��3�`O�\t����\��kk���a7�H�E��8�-hF��1�p��t��V�Y��F����$
�TkK�P���ć:73�.Kr�mˉ>�J���Ҫ~V8��z�K����J�W{���aƑ��Dʥ/��o���y�������������]��k���.o�hWh��y��V�TVT/F�Hu����G�.�Mm��������/�#;��^�v�B��F%*���y"x�n��%%fA�v�&Zf~�H�O���`����]O~R�
*���1�Lg���*��#��������Y�W���H��"k�v�K�H�N2WttA��-�w�L���;�0�)j��>��[h�]N���>��?�
Z7?�Y	L�lW2㓆2D�=�yO&�As���y���$���D�3��2�l�	Ʀ����Y�zE@���%�Cn:���ۉ���û���nP�Q�����zW�y꟫^*��R����EN�?������'�w+4�������/ ܓ�l��c�{I��9I�oEŉ�2��LS3]$�*\�2�H���b�(�Gm<���(օ��5�7"��q�x����#���*3�o��	�P��7�}˻��F��> �#7�%f�򾰢�z��F��̩Rl��)H�ȥ�D��d��E�+
���B����|���b�*ڟ�ь�0Uي�3�2�'0*yt
cX:�[~�W4�>����Z9�
�g�}tv�; �y������2O����Ewi�9�ey�gT�e��%s1ޯ=�g�4T����A��c��������*n�M�N�l���y=� ;pY��Rt�d&�Ff���I�Ij��QA���/�<psɢ���m���J����ނ���S���BkH��rOB!�=���Dэ��(/W��	!�h�0��%���|`��?s���	�8Fj%�;��q�H0�Q���Cv�ñh��E���͟%�Wk�2����v��q�t�𠒆�0�J�ͼt�|���B4D�OWEdQ��a�(9Qr��&}�Z�se��4�,NH�+_�)z��O>�z���^�/�g�SR%�ȧܔ,X05�Ⱦ���6:�;}-�����QI���j�?U�rFt)̫En�\T�@���m��|WĖ� +��8��r+�v���6�k�U?n4F<<�@�cq����My��1�е����	ÄN�X`)I�!�z�	1�Si�GRntg�J�������(/a B*��C��
!�;R��?b�~|fpi��=T�[��«(;|I��;�n�4l��)pCY�*�>�숞4m .?�@�M�J;DҘ|
�y��Y��N��f~�*A��DR��#����>>j��P��<��K�=��H0������GZ4]a�B��g�H
r8:D'F�!�$B6_��Ғ�"�}�C;�ȿw�0�g�������bр�W
��,DOy���$�{�/°y�a�և�?hN ���AC�xU=prok�k�͍�5"��>�c���>O9���@'x`{��gs֘���gc�tc��ڗ��'͟�n=8I>`��"�lXyz���4��U�=���#fO$!��o�N�A��r�%�.�!����Y�8��R�2>F��RQ����*-`��~�tJt��L��N����+ؔ´�L\�ϴA9� �4;ĸ /X+���ƹʴd]ng�����E@���W�H�oIN�Fe������G_Z��
t�2B��jm���A��B��6�솊���{��[�Ko��*͊�h��i+�AAAEa�6����c�e)�F�EfE�	}�\t��� (ɬ�J���r�5�� .��=�x&���z���.�p�{��D�C��D�o���Cp�層�;�{�����HT֗���VA��w��ʠdތm��j�u2��~V�=���9��=���R��SNܞ�I~Ws���MY���"�,���������kz�h�\�(�+c����P��ĝ捿�k��'����ͣ�7����z���0]�5Էq!� �J�M�	�'�퍀�C_o�xoAN�k>�wA;�յ�Uf��Zt;V���g�}�/V�y��U��Sf��ԫH--ۛ��?�}�����jۀ�3R�!BÊ��K�>FMm����R�p�v1�EP+f=�J�C�L�w�|��_�\�U��/�7mC;��i����ه��[�V����
Wf�`���[�\�)I��d���;y��l[S!�
+x�M��N)n�и���/�$��l�^dީ�	�ɪ9��Ù:D�G���ԅ����6 ���$~,��gO>z���x��{m.�IF߯b�(�`�꫹�*Q�vobr���$����6n�V卞�e�9n���������Y����r�C���R�d����CY������03����i�2C�Qx�η��7V$��D�u{�����:j�����<3G�x��WLǂ5?�*U��S�i������a�%�GإɊd��2�R>2EM>����5̮��R��=p��j����3f������\��P�Dk� O�7C��lX)��q啸��e�5�g)b����Ӧc�9����mڲP���5�@	+���z6�1|�{tҵ#Q���B�~�yӥX[f!F�9��_ya�!J-���FG�do��Ṋ�g�@"ur~����f0l����A�D���nV5�[��C�|�%�מh��p�,Ue�d_���c�'#�F�a
�ڈ�6����8k<*��
��J��8�\��T�fS26�ޱx�PGQ�2�[A أ�b˩�	�� ͉�����~��X�SȥQ���Ӽ�|����N��Cmn�i��f��h�Voi6S��B+�B.���.�p�9n��^��M�d63� S�6�@��q�杧I��!���.KÓr~3��_&H��F� �u-ĵ���`�������
�99�j��d��x�N�>�[P���u��b	�YH��
X��`�P��;�W$����γk���B7v�2Iw�00���J�������Z�����y�2�2��m�^�b:�0���؟�����V; ����D�W�baƖ�Y�  ���9yD�L����ʼ25�I��!���Iq tU��v>�g,T>�J$�����4�(���!��Q��G���~H��#ipz��<k�h�"Y^hB VR�n�!E�a��@{�S��+��K$��Z>[�Es/:~ |:�ώi����+#Z>���~RM�
���_ڷ$3Et������KP��Mm����1�]*��m��!�;t)���\G\&=�kt)�.�&�`ë���*�u�Eͯ�]P:��}k���m���Ѩ4�(+1W�;�{�?5�{b����ڢE�7��Q)�j��4�'�g�]��H��x9�A���"���`a��=D�S�JB
.�IZ/3ԅ:V��d̍2l�R\�R:́-��$�P+��D�`(+�>��A?c_�]b!͑͋��)�.����­��ED���x�M��;Y>���M��YM�����bn�v�(m@y���&��ȉ�3(fA��hf�����&����u��B�c�7uE�G�+iVP���mQ�zY����/j}��ҕ�O�����9�'��^�D=h^#��1�ꑡ쾥��.�`c6�R�Њ��{c�e����o�,�E��Oha�B=n>��kT���x�އG)=T!u>��)�z��B�"CrO5p���J��>���o���	:����#5���R�#�O���WO��D#�����b&:8Z�I; E��p*Ы�\��� ����%U`��Q.M�L#��[�*���,M�N0B<x_26b���-�a)�f�?��ҧ^2`C��&1?j
��E��E�P1�,�K�����'�n~��o�W_�
��-� g�hI~�x?Wq//*��F{�[����%�tX�ţ|N��) W]Z��	�{[����?�TK�ԯk�mJ�1P-��Ρ��w����o���Q|(�Byd���cI� �_.&����ZHw��H=Q�9l���</	*�"���5����w��6o��P�E�d��+Qb�x�zt���.�a�Q��1m��BK�"P�G��Ʋ}��6gצ<������պ���"]�k���?G����w�V�Oʆ0��k���ׂ1��l��s�V7C;�����\�Z]�&נ�!N��Lߛ�)[���s;s�
$|&1�s��[MjK�I��It�>���
qV($9��@d�J��Z�'��Dz�f��|�4wX҃6nҖo��,�'&>I-�\"~H��b�/fx����r������ilN���d�N�s����c��:,3+f��C[�(��+��W?肬�ڼ6�g�O�5�Vd�o'�L0#67�sM������1���US�j�
0P��2N���l�cm����Ց��ހ�#��Y+��?�\ݔ;'���1rͭ�6@�h������u�BG�A��D
���Hn<�G7�� ��%1���Ὕ�'T,-��S�<=�h�V ��ӻ�I����;ݼ<����ߗ~v���e�I1(����/��&�u��4Og�`rH������*XES�Ӗw��6�ѓ�!�3"Tqu��!nRI��?�Y��
���THͿH�����=q�ܶ�� ����@�:���$2�+��X�!��k]��J��>O�jY�~�R8ގ�pFݲ�����l*�Q���;�l)�%����� 	햀�v�,V=K�~2��r"=5�X��;l�`�c1}�1�K" �2���-��b��7���1�5j��O IC�fi��lH��Ԉ�Q��p������������I�SG)�xZ1m�u&hSm����!T��s���F���zޫa#�Q(���j
*__�l��� n�o	��/���|˜��h�W.��|�M(:����S�<��钯?���YZ��}*d(�_�:Џ��A�w��s���e��ƔE��s�v��h�Qࡊ�X�<h8��\��_��	=I���Jש�|i��Y	ҍ��UQy����Pt���w�M��q�V÷O�K\�O���-�Mz1�0h&�_w�%�Y���Ov�}q�GVq0W-���C�F��?b t��"�W0�J�yӺ������3R�e�P�VZ�Ɛ��n��0�H�!H>�md��f]���:=j�[��L����tH��k��	2	ֲ�U�v��c�ma�Z���ԗң�i��6ـ�z�I,�;���Ɩ�~�?�v g�]�:shσ��-àIhE����M�&��-J�O�z`Yp��_��1��}H�m��폫��� =[�~��I׈g����T]�m�+�,;�]y���KMGFz�%`	|���k 2J�k��_�Mr����g7 �b�%���}��fC\)�JY�\u��K��Lj��K�����r�*��-��!�@���w\�p�%.�DJ��0Kp�C�kyE�R�|��
��I�\�D�t��٨�%\WWk��XL��i��c��.�dM'�a���|�uE	� �Q���]L���|��w�H�9M%?��\�c�*|�r�R���<A�(�yf�v1:C�(����,,O	YC�L%�k�5>�Ñ���XU��������LOۈ�j�bֈ���L��#&4o��i��k9]��Ym���fO�t�ԬpV�N� c}1GI
�*�9�0��k�9d�B�}�G;T����jV A��%��@(HX�����)�3M��T}�&�f�X׹W��;�G���.
R��l�&�ut?�{�7FM+�;Fs��F�3G�_FԸ�ΰf$ܬ���b�ؾ��b����g�4ɰ^T!}�i'Q.[�Ef��a��u�mH))`������f<�IP�gY�*�B�9^>��m@����>2*G��;E$e�G�����|1�2PZ����H1�a�s?�

/%֛��dw����f�!J�˔�oQ]i�)�����1xO�c���	;@���h'DKQ�eZ�#�fy��5�мQt�n<��~���������|Z�W+0(4s$?j��-��62Lm�K>PV�#��ȣ�Jd뇪����um��f���*N=�ZI�6R�Ӂ��y�@A�h�FL��C>�~�!�	11�q�r4u5���7�P��h�0!?Ј�V~���z�l��B�_JBr����z�.�i�xsv�����@.�Hg���"엣2&ҭ��|F��G���kLYs;����k��� KjU�8#�u]X%��尻דL�%.�!U���y��)�Ȅ�I������]l�QKF�d�{�\c����
 �Y���R�Nt2��,�T�T>��ˤ���9�v
����
�~��t#�V���-�>K�E0���΅�C��me5������LK���8�9w�
��q>x�ӠRC�p��������̿]���p�-���VEjC,ژ�����a���|��E�h��z)Y���?�� Z3�>�;ޥ,]�ӎ[�����]R�o4C؊R�0�o��2�⒥R�a}Ĺ�o)2��������j�)v�3�O�!��JfX��s�)r�wR �����TZ]�i���(a��;h?eng���G�:?ś�y%
W�^�"�nKJQ�!V�o��$`�}�Do����͠G����)�?�&G�C��t��,]z?'E�O��q3f&�v�p�dZ;p(�P�(i������U߼:8�Q��7��\&r���-�:f�W�K����{���a�Ci���d&J�Ol�5(:6�d�E�e N潱b ��[_p�'��O��i�)"]I6%�'1ӓ��J� ���odRgz�B/W}Bqs� ܅s7��qw�i���Jr��_����V3�?��3ٰe~`S�(����<�F�|q{+�0A2n�kx�t���RX����a-��V1���r��z>LӨ��S8�B������zx�'!򫢧�Q�F �� <XpE*�'N 㖨��s۹���Y�j\����u/���+��y��k�:�׾�%X�Vqד��^����J���k?i�@��M��o+��)[��Q��Q�/�����9�qv9)w"E5��o2��5�T�]�bH
M!@V#=;�wmr�H��'�"��C�,iz�e�Jz��.Q x6ث���')��?�0'8����c�2�g�N�G�8�weq��nd�Q~ք�_Fڸb�PW'���"��|f�c_�I�J�⓲��"#���{�/�^��U��ռ��&�W��	m��N�}�=K�.�1v�6����|��b�	T�u8�F9����V�4�dKBh|������q�P�x�R��Y��6�pb��_K�"��5/���SJ�c���:���L��C��A-�"gh��u��t
���]I������X�M~O}$��/�Ŧ��հЕ&�c��shK�/qI��Z:4'�Yɮ�jJT��t��}D�9(B���Q�35��Ͳj[���]��;b��V�r��[��I�t�ֆ�u�˿��?��1�ܑ�r����ɘ��%MUf� ,2�>�<K`�9�Ii��O�6ja)��x_�Ɉ��0�U��#Ф�n2��߷dl܇G�FڦJ=s.g%Я6���̠K����Z��6�a]��o�P�f<����a��Rd���.�����[C���	���'A&LY%�sHQQ4�l��� ����)�=��l��"�b��l,����|iq�K�*i���1���k ��Eb&��y��H�Ї'ZS�;>����~�x�������Gu�T�]�|f�w���30h( ����z���զ�/:��ɡT9�4��'����1Ì���A J��]W�O�������z�l�Ĉ���t]�}�����pF�b����(؁e48� ��VH�xYAݢ	PHU�iW_	�������Zm�:�T��Y�݅ç�����A�}:Y�� �FBT�:2t���4Х��,�4�{��O�%J�����a��D髓9��>'Uh������O�ͧY���ƇT��H�c̖3��!�ͤ�ɠ��Sm'%r�L;;��,���XܓY���Q��df�X����=q�gT�i���\G���~e,[f_8<|����ZwN��/��5Ib �T,*���{E��	�̣�v��6��w��A��/�E��=:�b�Y���頿�j��.��E8T��k�Y�a�ۭ��� p�߃d�U/S᮴)��Y{=������v�>w���t��	?���t�L�þ�
�?��M���r�c�S�[�Z���e\�5��@�r��$'���W���72�[h_�ۼC2���0�=��R�]e��0aP|��B���Lޞ�{�Ϫ�Y��牒'���bH�O��hGNSF�U]���<�ci�
�'I��ޕ��B��s�M�"��t�<U7Tvy�s���Ѩn�� �� �i�VT��,Ћ'�ijC���>�h�w�v8�[Keɲ7;,���'���8���~aT21I:�a�D�ǔDY-�٩���C4KJvTf��BvϡmV.l#0����rjca�||�k;e��P�����wM�m��2p�$�@P��n^io���p�j�j��s�l0�O��hE�a�^�r�!踴g�@ؔ����mo!~�^�ny� �/�/�<�rY���w]�%_�39K�L�\�����ܾ"-�
��-��(���}qW����E���0���pd�l�;��6�͗��#��~���7��F�J���R�NJ~t�9���T�l�RN°�ˌfJ�4j�-	�2n�O��!���M;�<�.��]�±�/H��E-�-�y挙��0D�K��lD��s8z�~����SE���bR4��т;��4�����X5���(�<�%�P�j|�,�҄-]Z4k��1�*��ίu�7)M�
ِ�b��z֞���
�p���K�*
���_�ʑ������"�>�{����M:�%~
I���<��]S�� `��1
hȧ�
3 J���t��dc�x�٤���b����B�B�|Neٟ�ݟ���s��-�t�qp�c�dN������&;ЃX�Z�J
E�*<bx�vNv82�f�S�x��	��n\�Q�a�MH�3�����.��X�!&L<�\8��� 9���XAԣ�J���;_6{*�١7���7�b����<H"~��fzy��<_�bG��7�G?�j~]9G*O8�6Q��f�u�@f�>F�p��\�b�6V�7�i����+N\݁�������!���$��@F�2V���uMt(�o@GB��q���I�/*b�6��S*\���s���v�,æ	��s3J;�L�HVw,/��K1�	�>����~E�k ���i)E�ﵑ!+�wSG�Z�gj��R��^��>�S���5E}j�(���g�&j�ten/|�/��o��^xd �����&$-S�"����`8m���ɹ�.����+8��{Ԡuvl�d��؛�=;W�z�`rǃm�<��~W�u�V�d�Z���Om�<j��C��D%U1I�ߊ3���c2O%3*�T��I�q'��JI�%��u���Ȥ2_���Ûͻ.L��ӄ 7.��,�a�HT_���&��:��V�XC�`�*)

҇��D��x����%�q�%�����
��T	9{�K�����.ϕ�m�C�Wc ]*�m3�,)�w�p���e��2��R�C[
1��H5�]7?��bY�X��ie���S��'ѐV�!����tō�	�L��*?�D�z�V2��8)Q_�d���ό�SkI�_%���D1`$�ǥ2^��SD��]���퉝�Qwǡ+y,M�_�,l�b�e|���������/��br�Y����LLbi:����F�X�s��~�9@y�{X_�m���H5�s�|u	;��C<�<�M�*>�ɵ~ �-�O ѻ�3XS���9�Mj9xBZޑ�Az�T�B8�Q����4�',�
g|�]_BX��
j}�r�8�{ڰ�3�����-���7.
a��i��2M���,L�&�W�ɋ�Z���5�D$F�ڐ�K�.����0}���>�QX�9�E��m��s> 7�>��� �6ʴY��#�7�q�$D�|Ci1��Q�%��<�(�/��Z�h�O~��v�%���2���-θ�����:P<��ٔ��k�~��W�=U��ԴF�~���/~�1�73L���_@��h(�;����[^۹��q3��wro�>QC~�1�Y��)����]� W��-��te�&��(����	�m5��W�"5ߕ�!�k�y-�~�r몹��\_cOYr,�AGQ��
*�S�)Vv#YV�K�/8��IJ0(p���Ǚ\o�r���i���&���9�4#�1�p�ֹ�(�xb�:�E�"�@(h�U�X�ӕ;X�^�z*J�|�Yl��B�,/}��d��2D�k6s���[��r T�X֝U�*��*���J�
�Ք���W$ �m5�V���..�p��;5����3����'�!5�`���p=Y�6\_�,�A�[ H+%��F�g�1�C���"0��+>x�I��RU�48+<.��9�߲H�W����M��@���z�b�y���y�����/	�8þm�MT���Tq�����ٝ����LÇg���}j�mxB?�����\J��}�F����"u�#��,�|Z&��AnM�j�����BD�MT�P�wq��D>�T�ڿ�Kz�e�j;T������7�5Q�NӤ�Y�<�y3�1�7��a^�e'���d𑴹�sz� R+����L!(��\���~�+�(�,���PL�nz��QY1Q���Ĳ��J�᷇�t*Ǩ}Q�41tb~�ȥ{�̱#�Ad	�c�X�v���2Q��{@�Θ���rJ9s�P�T�!�=��#�m��jbp�]�k����Y�AǮ�u�+P�D���t���tkk㕨oO*�l��^N�f�}�`a�nP�6q�z�A5��Ue�����3�-�%���3-��Ӻ�3nQ(t��y>j�]V�_wҚ%���t]ۘ��ȧze[ڷ-�#ߖIo�q߇�~��VW�Qzg�pe٘Bh �S��O���jLk�2{���aʿ@��%T:�qĘ�|".���[ʷ}Ф��,���8=;<�
�(��Z�Ėa�?!r���0��`�Y�@ރ�g}eRg��ֻ��ۨ��:~	��'����:��\�3G�J�W����Q EL���ԟ�@��8��51��"M.�#Z�"�g%���FG}�ɢ|�E�;��w�r�7�[a�*�lK��yx�lǖ%9A���u:�8f�nc_���6�j{�+;a��n�Sl�q�y=�x'x���O��BJ�ҟ9�w f���h�K*{k����F�n���-*H����W�:	�̉W�Mw�bViD��q�{���묫�k��l��$��[=!��ٟ'���5�˩Lm�x_��L}A`���>�о
>IY�;c]�l�ʺ`��ݪX��$b�.A�C�Q�^��*����މ�gw��f��ɐy1��q:�JN�G5����㹥Zp.Y� ��®m���6�W�?Nߺ&�1Q:��=^�eM4��Y�%1����v�m��S׎Iц�+����klџ��