��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*���o�!��=e��O�	BIλ������sI4l��N��z~��������bW���v^���Z<R\=r�R�(�Ԩ��i*�VD7��A�����#0ٴg{��]��z�Rx� >��%[�Q���J�&��u7W��7��LP�NΏ����Y��D ֤˗�2 r���݈�G�O]���O ���mE��:l�};�� g�P;��G���a������{Q�K�ʃ��Z�˱ԟ�A�Ƌ�3w��/��e�P��sN�GƳ&*=�'k��Ȭ�PW���!�@��j�Ey}P.����=n�ãU���ٙ^�B���cA�H�h#V�i7t��4��`��ژ	۽�d�[c�x���P���e	����S��d(���4@Q�����+���c���!��'����58J���#�e|͒j��D�m��s8�7��Mw�V,�Ə�mmu���a"(V�*���J����mwP��r�	#�D�H�:�aL82��*D��hҺ���ָ���W0��k��fi.�.����h���;��f� 0���\pKh��+�;"/"K]8���P�BTí��̈f4�¤���q��0�aM�� ܃�l��J`~�nyc>�<G��E�ǎ ur4�ݒ�˶q_�G��+�{�tmi0�E4��q��7���)�C�Y< >��)��l �c/�~.~#��}[�X!���A�c�h*�z��RD�,���Lk�f-<�TG��i(�i��Fv )]B���<}Ձ�	��&&7i�?�6ޚg�����U�vrV�-�N�����d��TLl?�*
ql��{/16~GЫav�,����/���2�V8�Х��]�I����C.%VM%����AD�X;�8SP�_��!� M��q�$-	��d�)�5x*� ��Oheb��n����9=����Җ�gD�?����K��󗔱`���쭕u&a�d��2�N)����T�$~�� nR@���L��|�[	�C��/��r0�Q0�Cc�D��6�b޺
����'F�����\���̆vy��d����E�rp^Ҋ��0��/U�J:�����er�~��I��R^��R��[�n�	\�:�Em�3�����n��������׍�����G6GZ�0` ���_@�x����^I��#�^I�|dq��Ww9��Q��2E��E������vo�zf���FF��6�ސPt��dw^�Ě�8|�±��:(C��	���Hޜ�]�B�כ���#��w�R��0�%���]��JUZQ:�n6��t�OS���
�ke���)Kt�8��K��ůyVIs����o`t����'����I3Jۛ[��Z���4�vG�:�u���_`W/#�.uLiE�6��$� w�\%q�5(+�i0q�.i����>Ӵ��=loV�Z�*�+�m�ڂ�mU��"�(~L$��x{�e���)�H�%��>{E)�n+�,鶤�QЙ�fy[��`EN�?��b�9�i��n�����w��@�9�+�.����c��
�ֽoeK*0������]3H͕�kl���ˣ�w/�d���!�5]�ˬ�)7<�y=N�t���3�ʼ����Y���Ǵ���&&O�;Œ��b*v�,r�1j��H���C�PV�Ĕg�nps��L�DtJ`G:"o=ܘ!V�j,i%�
�l�!v���b5n����A)�~/v�a�m���;Uk�R|L�7�6�թ�UDK�cB�H�Ȯ��Y����	�f�I�D��畓����H˺yKz<0��f�s�?����f�~���F=a'����9ؒ1 ���̘�s��y)��6P�;��m�DIx:|��ˏ��HD�82�s��R
+Ե��~�Y??ڟ8^��=��H��3R bf��0;9v��S�;̧;�@QO2��"ζ� w3��L՟�Z����	rvG����i�W���V����+q`�R� �`ޗ˜9��WNK'��Ȫ��s�A�C�*p��l���M�u�n�
��O��w�\������y^jt�_Nmy����1�o�r8<r��ޣ��6�S9��R�7��-��|�h�O�5m)f���v���&�o��褏����Z���?H��3��h5�IU�@�i����#Y�5��^�*,���
�Yu�M�H�Kǌ�Z�t�|�^�+2!�(Y6���*�ޣ�,V��^�YmZ���P���h����ȼc�,=4uC9QO�~X[���<��병�Ҕ}׫�iOS����I`�=AA��>�jF�Ѝqi��U�����q��ȶU��K)(�|�/w���:5����+��FE|�Z(kK&m>���*�$b�'���;.�nV��<�x�Ǡ(H�q0��n��E(RZ����i���3����T�|�O��$��R�ϵs$�����`�RhN���ٶ�+U��v�|�s������R��$���e�)��D�[�0�n)/3�{4��w�[d�l�eD���Q�6טP�qW�ey�&���NټX��R�U�Agl��&�'�3�
%��0����u�5��I�"�W�
�_�ȃ������C���Yb`'����r;�����1�F��hZ_=�_ib�͸���xy;��3���[��ࡶө��9�*�� �̉.��A������+�C~c��"MC�H[�����S�Z]7�j��x{%��Y�/����\o�,T8?%�(5l��-_ٚ"��
�[��u�f �X��VR|`a3�K���z�xiI��*.�Z�G���2@��o;�,��#7�w��z�_��I�Y��G�c��|�=�����z�|��T2�ǳK1���t��rb���M�:>���S����&x����9���eē�x��QU�d�5��1|����ȺP���̱���b���"_2�.ukk�[A���Zw��I#�%�4X���0>)/�(c��L��� ;���h�0![Q��;����e�>IJ�e�D��'�Շ���Q��S�Q��S���p��B�7v�/�ᕍ=��r���r?!?
dIR�쭟�a��\�Ū>G����������(�O}wA��ߛȉhF@����-��g��ERڢ���@S��D�!{z��&�T~#W��u�v�jIW����KW_� k1e���3RoVb0����[���)�^���3*]��(�0��َ�T�
.��gi:��#��S��NG� ����{��K1���<�JIȵ��ӓU	Dut��w$J,.����w��R}�YqW�gJywZH��-�]{A�7|�)�O�6�E3^�c"���(^ce�S)�fw�L/��H��Ȕh#��{�i�ȭ�^Q"*���������'}j�b�@2��Vw�Ӱt=��|M�5����S6�˝�	���/?�:]ۜ�ty8�4����Ix#��{��)�Fz$�:�Ȍך�	��FH(�$EHG�$���c>%`���	f3pk�f�#��W����yl`t�DM�.d�3�M�+�o�	�H��*g ۚ���RZ1��i=ȵ��$J*(��9pT֥(�L�%����9���U�{��%�sO_?V^�\fg�v0/� �S�́H�qd�9��
���
�g�CG4��*(
��Tp�N؃��1�/]8�'�d����濙�" ^"Z�R����J=��Fp�QS�z�2��>�D��n%_2}CC�oӋ鐬�b��	k�d=q�^N*�0�U������]�F�( ��;��J��ԅ�2�yI���O_�ʔX�{DJ8Γ?^��bU���4E�>��+2�!U\���5>�"7-�fY��Q�K��1��㞘f�����e���l<>ue�;��`.eD���B�t(�N[c�k�=���N��3�T��T�v��q���g��Ѓ�����?�#���1�nEg�e@i9Xfg@�yX����}�����^~.,>P��r�k[��2��EwH����������I�_L��/Op����zR_q���8���Ⴙ&o��W꫁�G�t�]��G{��%%���\2���;c��M��m�[�[xLp�LjI�u��ʊ h7j>��kf`k��s0�N����|��d��{?��k%��s�.n�lb2�ox�� jU4%&���Yy�x�̡(zu�z_RA�{ׯȇ���v�N�i�G�b-�+|���5�OFꝕ����k�0�D���� k�Jf��!���Pȋ��0��tC���ǜύl�Hܿ&�������ʙx�8�tl��ā���� W�}y `휼[#O9���Y�þE���9��=��F���6J�IZ[o&�̙Q���Tm8Q�R�8v\:���4��ϫ���07�Z����q �,�hXi��;vJf�4`ɽHx`Gw����2���}.��IC���۶�������B�.?�
��j�==�6糵 ��ɇ�'S��]W0k�o��D�]��B-r*!�����p�v-�ν���C�A��8.��{Ć��d����oI������{5��l�J�z)f!�ZL �O�si�%|�Ί*H2�E�����*w��|��0�8-O��%WaKB���b���.��W�/�������e�,�~^"G@���1�賓��n�c��|h�8�YKr;Z�*>�$v_��T_!i�y��k�mw(������(Vfp�E*� �}#t�PY�z� O�-�O�8���n��Q��H��7e����<*Т�m��H�Qw�u����B"rX����h�6�sBb4�Eg_m����Q�ե!���a�����ݣ��`)&�J�r~M���V"=�|�f����c�\7�'�Me%&�H�T�����<�����0�S()��s�Ƴ&Z}�
����B��ߖ3�[�<�1]�gr٧�s���mD���EkK�Bx�RT�ll�	��@���FA��1��)}�8��j��C�t@��-���z�.���9ݭ���Юy���(����+����A��1Es+��ɀ^�筰=�!b,.�kC���*�Ɓ���&�CWJ�D��h��'E�a?��c!�a����vs"�den�?�ȵs���؛���		��='z�73�ݍ����e��}��!�M�E}rW"D��&Pi�|y�P�p�t��02>
T4�x�9:?7��`;fau<������7e<V�E� �u�%x����*�T�T���8C{*^��;N�~��e��,�s�W$���jC���;{�-�K�F��W
}����!�4�O�"-�!B�Xd��%.� ��j��~&�z�5�KA6����/\�WM�^W�/���T�r�/���ۃ_��5ǳ� �o�p�4�|=�%�|�-� �lQ��-����t���l�l���WL�	�;���l /8�r����1�d@~�E*�~�ǆF:PZ�ҢWI��G���a5@&P���D�{���Q���A�{�G+�w�ɉIu�z�)�xI	��B�S�CK��¸s��Y��j��#���]���J��K嘍�D�B�oV5)�o��Ļ������6���E�j�<+��{�����z��9���Q��wN�����%Kׇi�g�F�~�L�k�"-E�fn܇�ff]<�Fl�U��1��d.,�/�e277�.���wO�mب�^�F�<�;O0�e5�{,b5u3��O�g�4U��N�8ы}rг}�U��2u���<�)ƫU�$�5I���9p�
�O��ٶ���O~4ցqc�A���Cr���87x�r�#����X��H���|��oh<��m���ђA��*���f0��U�3Fi�nKx��`�o!V{R�<�lF�<�( 3[5����p�w�
��
�d�F�c:��sY\'0�p�d^p^�ȋ7c�>Qm�R�]������[���m�#_������}���?����vY�gS��">�p9�J<��N�m)�
�>�Y�
���.˩�&hg3K	���$�& b�΁3%����|j���=���H�'����Ꭓ6jJX�[���
7�Ze���;���U���/b�PA�Dc�֘u�'}L��Zل���J�?��(a�\b�K"]��=�����wK?1yTTo�XJ�ĩ�$k�Bb���;��@�����v$�~A��e��:�Q����]�W.��:���3O����wo�~F��\_�^J����ç��]�l<����iT(�V�1'�R�/�3��t1m��yGqT�`Q��;6'l��P�,9eA��W����cT.�Gm@�m�Q٨kx��sX���y��"M���M|Eq��8�a�*A#�uN��i�/6�E�d����a�>��3: �(.�fʢQ�����s�)vY�C$e	k�zF�d��Ί�#��^LQ�]+0	�2�����!S:���_
�:/9�=�<! 3e#sȢ^�e�~���8�{7��x��"���:�0�	 ��NtKx�E(� �Odd���k-O�X:X໳Z�l��q=�U�\�Hl��?��F�vqآOi}`j���?z� jl���RN���I��U�U5�0F���7Y�(�vm	�-�"���0�e���(#:�$ُ�* �.��'T��w�t���'2�P?t��a�L�א%V|���[�����]�R����4���#V�BA��P�����r/W�`�K]-xҽL�"�g�j��������P�B�p��_�dT��j���t�ΦaZ6׳��#�R܆��}/�V2�����6��д�*X4ÎQ������8�ħ�<�L��zG�%~I�Ҝ��r��#&����^��M��u����M�("�����Nj���j<x�~.U�<�7:=���"[���eB_�`�ע|�l����w���R�H#Wp�' �`-����i=[��c���nos�U[�g�A>�8�ncUV���.>10��9���l�"�i4�O9�]��C��_y��*����*�{�-�Cz&%q���W����Ϋ���	�j-篗b�i-,����!��#��q$7�q�W�����[�_�*�?Zd�7�8Է*\Ûr�P�`)C��=j������sY�.�eYX��3�*���k�.<����J(}Z� .��m�Y<�*�+��[U��x!mY� ��c��7
n��:g1��FQT�Sb
ξ̡(�,d����C����i�;��m��T�����}AUK4z�:<��G�nSA��UPUE<����ߴW��<u�&M�N��wiE^�<>���z��-�����B�}��67E�_�{e2�^U�K�����xq�o�1ˆ�J�\U>�I��B��QP��u��ůP9y$ϏRm���(�)`����A�v�*��¯d{(kY�|��J%�H��Cd%i�Ɩ� �=$�O��R��<��f��d��b,�e�e���y������n[����y"C0Y� �o�L����!��5[V
1�xB��s>�XX�,��,��Bx�<�dkiK�^��_�ctQ�u\���%��f����V�N�K}z�p� X�����twǤa�B��v�/�`���]�s��	�F�������b����O5�Z�{���gs4-Nu�0�X�������@k-@��Ξc��ݮ1�.��=p�Uk�D�0�h19�k���!���f:�Δ�!#��׆�ɲ��] i�����1}�����5&����]�;�r�������.V.m��M�\��(PD��V���O]S p��(
�8��ڇ�0���[�9YY�8�y�;}9�l>{3��fy����;nM+!�	����YH��`q��f.�$~i�Mϒ��|2��z�Ζy7��|�gF�$�X�Ҽ.)����AFߠ_��O�&p�������`|�>�ZF������c����Iɿ�k\5�6m��̺���{�#ErSЂ�{Չ��Pz{�?%~ #(hRAl�*���S���e �4{J���"�3�5':h�-Aҳ\�ӄ�(#��Z���}4d;�^�IP���!w�u������N7.��*Wi���'���~����t������ۑ���Di{F�d^�\�@ɱ��9!�ד�G
n��ݱ�z�vq�b�����ys[5�.��ٍ#��M��q�5��\�8�la����(��<lR�|�W�]+zJ�³���z��$7���
�R*����^-f�L�n�~�N��ZIB�V.So�c��}ɯh{�+��^�����#ٻ�T(s9�j�r�.B����-OwD��8�Z/��%�!V��[fn���W��/��!v���iP�-0���p�i��8I�K/o�T����rF�RK.�f�g����rc������pQL�\���>F�����E'��!�B���RO'Wf�����j mW_h���]�@}��� ���Y��>T
.Ne����<�7�>4&�|7�ϝ�S��D��d?~`��T�P�����_���r�LJ�O�p�G�4�m�@��M����AV{���Vy�@�Z����%Yed!��O(�����*�=��}�Jy_���w�TP������~a�4�Ε��9�(�ɐ:��3�V?�S[�ݲ������-B�}�C^��� >�i2���皆	�Ǜu���>��QN��3��2�5^���C��r�a�{�g�̸�i@b���U`>��9T�
)�����f&���-� �@]�Q������Y�k�WG�#�-����R>��׀V$��n;�{>|mf��G����_߇ًEo�1��o˺�	iY��u����	fN[x�luM��d��k��+���3��y���7;�u�C=�������V��[@�b�A��@o�!��=�P�����,��XG��#�x���(r������)��<�Jb�eNv��3��$��=��`�t$�VLM⓮_i�����g�ds��1J36����I��SPA��S���.f���f%��������eQ���`��W�Dq ����O��R�ŝ><�d��f(L*{*ڽ���s��Oh��|�&�=:o��� T��kS.	GUU�(��t�'�#�v=�N�>��1C�:��t"���W,��I�%c���`[w5�jh9(�s��.��q}ߛ����Qjub4��R��\L���I�]��Q����"pl=���Rg�Κ�SaA��'����.w���Y��ԭ��G�lF�0����F��ʼ�l�����^9t�/���bt�����{�hJ�(�i�9c�0uh������HT�q��[��*3饎���f���D$�����;�g��r顙� �P�9�����+K��qߵ����P�K=��W�O��`�]�cw��d�I��d���v�֍���#���ɽ1?p<t��
��>v��qȦ�B��]p��'��]�EQ���'��G��$�0�;��ľ��$�L����q(�ِ�=��u�[TT�j9�7Hg ��]x��'V�o�uμ���sJ���g#�@#�Ƀ��-)iR���k�����
tt��Pb� �=h����hDŗ`�/��[�Mj��d�Vqʀ�'��K�M�=�57��Fe"N�$.c���8�g��� �u�!Y�Bɘ��3����+���6�Dl+��+��u�/�<�JɡV�/�/U�Z���s��BYPԨ��bNLi��Ј(�Y��T�ROԟ�LRw�����*Hl�U+����ғV	7�\ި�
�牭��^<G���A�e��gf	O�~��zy�1��a����!wa�Q0ŤK�(�C�F�D">:�áv,	�����t�zs�[2�Ԗ�?���� w﫛,�C"�!�jz����~��GLv�u����t�-.������u�q��d��n�4Ps�s|���n���5$6��n�ʖ������:`}�C(�w7�F��6�7�ˮ"A]��2=l�M���7j��Ӭ�=���IP{�ڵ7
�9�i���eO�p(�K�����吻��)
��_���~�s��;U⵨M�|���*wڻ^'�9��܆��'M7P�Ƒ�p�w�8�F�
� �s�^C*�zC���h�9W���A4�����)��\��a�����zm��x[|k;���;�,<y(k��,��}�=���b��y�
o�R���>��;�h_�~��(+I�0O��i�?�N����� ��F��������K��Qf(:7���e�W1W��1��DҠs��v�-�U��� |�ܘ��
�"���
d���4II���l59�
��<�H�Qǚ����8*���	����
J+�7�/�a�1��O ��%�G8=�����$����Ii '���FW�۶4�$Ȅ_�vfs��@�����Ot���T$���F�Ԑ^���y������Ò��s�:�[����q�9�Gѝ5%���Cɍa�C�|�:ϼW������Jћ�p����g�t����rD��2�Xղ��T�F_&��5Ӯ��w��^+�3�ZU�}8Jm�rbOa����A�P�gt(+�E{�T���~Q�^��@@hC[������%N��U�G�uQ�e�H��#�v���G�)�2Bڨ?H`���_^fع��L�	}#n��>O��Ǉ ��3�i��B��c	D�ǚ�vp=i�)H�>�GG�)7ExJ���Ɛ�>�v�#]�:(�7��E��H�$�v�Li�x��?�jT���%��ѹCfF�R:�S2M�[�B��'%���ٝc��*W^6�}ܷ��l���Z� � ����<��*�B<�T������'4�״M׎(;�H"? ��8-����S��<���:���d2b�͍V�3��G�C<��Ŏ�sl\ͫ'���=@��x�~�S�I���7e��@��Ap�u)8K~e�����t�:�w|'�0_	`���x�R2�yu�l"&(3�F�4Wl���,�ѿ��p�6�������}nf�Y��ܾ )'�o�|≍+�VAr��/�:RxL_�<���F۩�]�%��_��pņ�
�Zv���}C�(5:��2H��Am���,�������׹B"�;�i��ܸ���\*~(��h����u���򂙡"Ӧ��å�ּ%�Y�2�HF���@<Ѭ�Zk;�AVVVE�؄�+��̈5���$�/�w������;��Ѕ&����H#G+�(�D�"o,ȯRW��+u^�rAI����j�oD��]Kx���^v���%�z��I���W�w�X0�nA��T_�Fcؐ*Щ���H���0��y(2Lt�����D�b��k,XN���>�b*�2�;DN��ɬ���p�x&#\E���ks��4g���R�)v���d2*ƴC��K@{^U3�t��)D_�삇�u�[��ה�	�Vz����d�ص	N�Y(\������]¤;5�������� e��͝?j���hn׊dz�5�_�Y}��	-�H��Y�4<�Cw�B��5>��j��b�k��6!K��|����~p�_��z�#��/ޭ�m:��t���8a��Ƭ��=%K��Jg�m�7n�d�&q����_H(	�oB�R���<4`X�V�Y_���A�g�,@�����#�f�ۻrF X>�?�Fڢ�rN5���]����BJ��'��߽�;�vyDn`�1+JD;9tX���OU�T�^��S�[���'����P,�>�m�Ic��R�~�/�m��ނ�-}���3ǂu�s1�yO���U�p�"4��'�%��Y����G=�	�;�o��F�����X�X'��� �wm��WWy?8�m�5��OD��O�������M�{
��dN˙f����	3�K�	i�*~�#LK�����t�G����aڛ1���4t_LW�+*������
u g��=� �s]�����$+?���*1�����+B��Oa����6��9=��A����&�bA$xʯX'@3�k�g��X>��I79V�134D��'��u0����A�� E�	�9�� G���q���|`��`i�_�(�V�~ּ��!��*�Z���:��u�� �����)+�W�,���i��w����L&���tًC�,��<�����G�K��~�TQ��bF�q̞�[����/@!�S4ONq�����4,�{��zJs�x�:�ƴ����ܤ����6 9��?�_vr�٣�� 8Y�2:-���rs����%�h�q�	l{��0( [_.��$s����8�۝����JAqH�i��N&F�����%�谈�������ϓ���<�����x��J����������5u�vp���rά��J�� � �\hӁi�߼]c�^߉|�]8��*ϭ�Ai����ݏ�ۻ��d��J��2�h��TGL}N���=���2�A��1C��P� Q(�oK�Z�tPaP\�u�Ћ���
m\ф��?1��� 7�d��c�	�v:^�Z�M.u:����D�j[<s���a���0_2J�\�(���Y|e�G�n {�#���c������a:�M2l���M�F�H�ZМ�p���fMr������p�.܎��1ilX���^ �'%9�4�bi(O��	��?��FT�c;�w������O��z����p�>��`����g�$�l;�r>�;���!
���K��J2�JK��o!܊��^ i��J;��08d�x���[���P�V��BQ>L�ް�vow��S]�q�Ka�R�\%T7��l��6���"�*dH�61~e,F{�R�U���gt�����\
f��Ѝz�"I�A���Z�(�<4��̵��H)5g��,ЄPe���i�\:� ���bb<�Xu����i�㌯Pʏ|���ϓ��xi�֦8�-�2�W3����S}�[��3Ƭ��3��߭��ȑ/�_fG���#���@V�'O6c)����+�B�G���5ǓM�(�E�!�p|Y���ɱ�~a�����:뺃:�G�{����|�WI��0��7��,�WlO������/V��ߩm𦓸�*s�+�*�w�P�r���,�����:��-O���oY@���I�[�<�5��!on⓽��j;uqJ����T�dߢ_�4-���0�s�3�����$��l��x]9�'�6Q>r*�^�8��3)씸Ö�f��	�a�)���<����Mp�p'hSr5�T�b��kǰ�����l��ŷ8��<��+�������'�\_��tf ����]u����Xz��W�jLD��BqO\r��х��T ���M�����^%+�>g�8���?|�.2����x��h&}�[�8�rɦ�uߕ���-R����{�+��螩�l����!G����tS��#�����ҧ5[���t����5��x�ډά�J̗�8jAK�GŠ0J�7���!��YA�[	#GA� 
'D�3=��H`���i�������5w?���;�6�j�H|k��� �-tzbͩ�Z]��I'��i�������8+pn(S<��������w1]�fR�l/5H��0��K�|w�9񗔕<�?B���A� `�0��sZ�W�	q{3�B��?�8�dP���5�s��NJ��&3��+���y�Z��v��|���̂�χn}~��
��q�a�H-V0�{� ��3@ǲ���^d���-�OY)��YRT9O�]\8#:g����J�t��]΀�o���^�|�����u`�A8h�OG�LB��\��rk�\z��`ղc)�y���P�mh��_��3�����8�X ����N����]�:0w�S��5��c/}{3$�/�(���a�Tˢ����.�ך����KM��"�?Ս���OW%uu�v�
�z5�.���ԡ齝�W�-�;/�3��\��9s8�+2���)r��!4�$E�w�4��OV�	Dó����;�V1��������S���-���Tp�����^����l�ܤ��ܰ������{m��]G�1��|3�7)��� �mxD{���x�����H���N���d}��i��xߛ�Q�(�L:Ju����`�3T�1J��&��<���q9�h�~�U��i�v|)_fMg�a���0��[�
uk^���.�"���ǒwo}3K\�s�:�H��(���1�Wn�.a���X �u��������$̴�+�LOJ|����Z0���Mj��l�Yy `b�?�A)�~4��~�A�q2M&4�L���s=\Q����DI~)������5u#"� �dʍ ڣ�D�L�b���,�tW�;(��޹����9NNy�k�2�;;���4�6�Dȑ۸�m��89��V}��4x$�C����RyWv�O�FBmk�p<b��wJo���ZA �}���/�#���$O����� 9-����EAI�:�E�ߴ�M<��E �_��Mk��K�-�l_F�K��;�]�w��M$��Y�W�L\��Na�$b��p��Y���t�
��0
�%�%	�r!n	GD�U�9Cz�@���i=�X�gv��q����M���	i��'2�v�0�q�؁�R3���`=��QDb᧕g@M��|�sQ�Z�U��eՉ�\E;R��[�vxFV���5�~|��/}.C�f�4sEw���O�by�s?nE��k��[���=[N�m��+���Ν�J��; ux(�-��>�F���r�te��GL&��m�aa2��������/k&C��v%�n�~$� Mν}9��*G���W@(�Y���x8�_�.	Eh���qbk��`kԨ��s-�y9%�������m>ڒZ�x{*�p��'�Yɭ�0e�$zȵ�@��m�{�W�!0���G�UR0�j��(w�(��PCl�B�۷�$�MQ�8��P*��
�wG쮒���n���%N~ĥ/^9� p�hx�jPK�y��Lp!&:�z�����*W�<��5�Z'cG��[�32�oP'��N�'��G4�J��ߡ�$����c�m��t���90�'�u�k������:˸��4t�ɜ�^0Ȇ������O^8�rs���|i�%�	�ۊ����*���{�b�6�E�D��0	=���y@9ҋ��5�7!p�/g̖1�wv���U�"�v�Y��@�(iG�h_��|�I��.6�W�9���Њ5k+�/`?|V	 M~�u�J��Qvt��Ks�>��5�Y1^������_�\���m��&�e</I\J�r�}ѡ��0�h�x��p��t`��\x�@��ryɃ�c������z耹ʢ�yo�vC��|�EM{x���L_�6�'1���h�"L6H(�s_H�%z���1��Xy�W1[3���3���X�O��������\YP�؂��%-L����Cg�d/�v}!4�:����ަ
x�٫")��I��fswG��ͩ�4%�-���A?0�Rȏ������M�j%�Ɉ^j7n�n�q_�Wv4`9�f=�DP�D���/2f�ӎ�'nL���i�U6H<���}�'�1����Y�-���Rbfb4��L�^��=e�Ĥ8���apc�NƓK��]G��g��*�ؾ9}̧��� ���9�kv�^�2;�'����wҞC�?]�&B�}�+� Wg�v	��c0�*�$ni>%�]"��L��q־�NT���
.!�7F�<m�1�h�$��� ��!�Ԭ���o;S��G۪�`�f,�t��@tA��ch�6 l6�u���;x���P)�1]��O~��:k2�b9�{^^s��֕Tě��K��~zѩ�I���y�܌Q�����Qy����XB2;U��BO��.Z#M7ơ��uA*9���M���C+j���6�X��lE���q����I˥�����<k��ѡE�<$�tg���!�˱m��+�F�yXr�݂���D{4�,��c;OQ1��~ɯ�C7�7�E8��"�̧��ƭ~�y�]��zw&���lO�h�^##�p�V��f/:(�!����ΰ�_�>�Vg�i;��7�b��[�*d�:�ɀUpYrv�o>E��%H�S,�����C[����Z�pK��Z��Ē�F��M�L�����	��Bޝ���8��UH���̞�F�\���t-?���� �'�/��Zj���]gj���q��sW-��x�o�L��3F�8�/-��@g��'�D[��z,OJ~Z���zW���[��?�HĀQ��ҙ?O�f�4�����F����Yǖ�O��-m�ۼ>�8�`������ c���;X�B�Bt/AyCx:�ɥ��nL����ʢ��	�~/��-(��5�Ʀ���&4��Ya�V��Mv��G닾K!EpO���ҋ��Ҽa�̺+p�!�Fn�t.���R���Ȗs},$��G�lo[ψ����o�O�h�f//.Zr�3��>{�{j��o���ދ��P�� ��W�{kή�s�l�j�q�g��H��A��/�R-�b��|����ä��v+�:��
�_P�&;9���n�!�^4�S^� ̨f7�ؓ���0Q8hy�z�������h}���v��D����Pm�	^�եJH��dx1&C�{|6�|�.���։z8���}�{������K(M�K�L��L�{���[{���|$hl�vx�[4��ĿS��2v�����o+W��/��א����kk�eU��1��X֊(��y��J�dS~[l�}.�����;F���*�?�m�.�o� �3�����y�b���{)�.�Ė�΃�a"��HR��ŗ�G������a��b��DS�C�������m�ef�r-��𬵒Qg�}O��|<��FR��\tD��6לk"o\*aG ����D�rL}0r�~�ճc�'aT���\c�w��<�ҝ����e���s2�k;��|�¯�3���]��ֈ,��=�ߛv�{�JT~���_2��s*��e.\��B|M]w����K|�	L�kh�˵�Aim}T�$O���9�c,��B�hrZ���UT]~��b�Xޗ6��N<i�mP��3��t� >͊0d�2B!T��m,��}n7	K��71�~Ӟ����*�4�ѨfXeЦ��r��~ަ@\�D%{��o�HTs�Z���7�#8m�e�h�/z&W�j��#߮���/�tg��
;�ssP�$�%�0���Ǔ�/�Ԛ��BnϋvĮd!%��J�M�2v�,�ّ�����g��.�a��ceb����8�-ޣI֍�m�F-�5�f>�@�8��e�A�h�&���a�ۦ��2�<�c�d���r�-����чg_]��m	�gL�	o�5�n��+&�'�?�h�L�e���W�x%��L5�ԓ��ږ�ZZ��KRp":�jQ��wGѽ`As�⸰>\�'����d��>�!֧D����х,n'�n�ڴ;��@.fW?g���Tm���|�ͺ��9�l,�!l�Qv�zp�D�S6����	V�����ͥ�� 1�'L�ӷԖ��	,H�C7�����d�-�P�~��U����G�:��(��
\߷.�6��r�f緂��P�X�jK� �|2=�
�&�1^�����8G����$y�#͇[f`�ӌ\��D0�<�c�^���N8yW�$Y	@nG����j�WM� #Vv�^�s���J��fe�7Wٲ8ב�^уi��)�w.H��z��0�C���/D�6�m)�����w�� �-����@���L��<�~��ngn+��>=��;�$��w���K�]4uy��`OⷫA�q��<�v;o�G�h.�p��+f��uH'�#��U��Z���������g<��1�`,�{~D^��VRC�u�᪑�ꐡ;gM��Me[�	�I#\v�kzu��u��g��h�Ņ��~�	fB��C!^���t��m줇~���q��c:�e���ƛX[ _��T�8'�T�Y@�:�~�SҟпI����-WL���\Q�jۖm���9����F�~�>�z�����2�p߸������r��}���@؈]}U���"m�)0R������Q�Q6�\�?���uX����|�lj�^�~e�%AL��6o=�n��/�['����,��ም�uPM��������C����g�b|*�2�����gX���E_��x��P�\�
�nɃ�>��	��*�Y$8N����r����L�V��~����N�i���/�������pn�Y�wirMge��[������K[���T��Om����M�Hk= �

}J�h��d �v����u�L�5�Le���P�)��]tJ\�/a}A��uȅ��	�#�r3������"�P�ۮEU~�[���X޸U����� �/ҕ�¨og�#�nW��U��GH|����ɉ���q_�Dиi;��W��G!�fD�����!Vk�+�	o������(���g������������N��W���	"���A�}K�<D0BUc3�4�	D�gBb������5X���0X@�y㶅7��},�ߩ�2��%ɵ�'�=�f=	}��$W��%�]�#A2ld���� 
?ش��W'��@~�NM&������	���^���ϔb!�cۈ/E�)��`����w���L}5K��@vq�OL��w�d
ݻR9.pG_�4�ú.�5PO���H��Ƨi��[�}2�.��^��9$�J��s��z�C}�%3���4�`f�uG�Ğ�#�_��Ox?��3"G$sR6��8��.-��_<��u+%�=� ���]�Ԑ�Ť�&^�P�:zH!M)���p/پ?�, \�+�q��eG,p�Z����υ�[s1}�Jn��W�o���5r�boY�q�*�u�o,�Ţb	=�q���������M�踳J�DƂk�v�n[����á8=�J��Ⱦy�xs���tha3����=:����{7��Byp��d!�fv�(�6��������<|�S٦�!�x��P2K+�|�\�������W�BTY�K~kʽ�f p��g�Ť�C�IF-͉n-ߏ�#R��6�b`F��.p��X�F��ʏ�Sx-�́����i(�$�o�u,����T��`��d��Vم��yX��P�����n����Z��*R�S�'��jd�`��-M�#��L4���3-��t�*m��B�C� `���Hxu��;��W�����}b�K�;�ԥ��:�i�'Rg�����ˏ/�<�^0�O]d�fa[A��M�&	��O�}��=�΋
���4��6�(��p�����CM#�a�o�N�$�W�f���@r��&(��{r�Ҙ��f�E��ϼ���@S}� �-�s�����#����)�ڂ3�?kn)�"�8:I��wM*$aB��KV�W�
�j��̕q��1��n��lĥ�0�2����Ͻ���k��$�LT�DA������ا�dg��\�= <��K�P� b���n�+6�
|����Y�7E(Xh��-��¤^��.��6�^��!q�Fx��:��LGR�)��8_�KF�4�9��G�$�7�rE<���NOjn��Vܧ�O2��� 4Z���j�j);9Y`��r27h���:k�w/C��!�p8�L[Ґ�F,1�����N�����cq7��`{�Fe98S��@~u�"'����=���`��'r�2򺶛ࣆFj�6�"]�c9̃�b�n5��y��#n8 ̈�����A�LaQ��?)�+V�;"B����4���ec{��>��;��Zg���^-
�5�ơ���m�J�o�q_H�!a¸���h�$J@�dQ�/7�đ�v`�w��� )�"8/�~ʿ
SW�1T:,���'��� �c	�4���m�#�g��n���τ:�]*��J�#L���H)�k0qD�D���d���ob���z����>�{�(�~S�z�]*�� ���=/d��݀�u{�t�E?3U�x�_�3��2�����f���eoj��TM�n��]fx@yP9��j(�i��Nk`;$�E3��BU!�䪒��=�ơ�{�&�.I��\�*5���v$)myE�F�m8Q�~�T :?DHn ݣZhn��T�Az��m =��J�I�Vx������׫��Ƈ�q	q6|Xy?I�ziJڍ@��T�!�g����e FXp��Ku잣N�Z�0���I&2,���g,o@б�-�O�y�2���ZG�������<�U0�XY�+��)/,&̯��t�&�,;hZ�N	0�����P��!A�k��������̸�"���(c�g��!Nh�I�jkW�Npƍ��wq�����ց~>d�t^f�%�����	BDnX���O ��c�$�P�ڹҌ�n+w���~ׄ�Q���va98ِ9×rT2sK^�"8�5-�ÓR��'UV:~3���_��}�gE h;��ӡ��Rk�d^�X�#�.BO�rU@�;�y��cAT��G�U_{��
�j����)o�s�
�J�*����y9�?G0��|�i�a�%�Fn����Ζ��-���E��J;"����>�NXer�����P�ݏ�_�1��X%4��J�!6�ע�jP�_�/��M��i>/ŇE����dK�4A*���w������Js$t_�.�	K3�5�Yk�%+�;?4�w���v$�K���1�H���y7��C$[f�����Rl�+l\��ݣ��K!"$+���8��(d��*��e+�GE	�i �rj���:����)�[�EK���V�VF�Ѭ`�ȣ��~[Fsj!�kK��\*`�M�����9��"7��?c9�13�$�o�T���;�l)�+u�X��'>��a2ɚ��@�e�Ԭ�!Y��))�ޮ�j
�q��{K���<�5C���F�#��+�\��̲&��V���l�<Sy���쬈`�����/�i����4��L'K����q����J?��t��u߾ÕE�!c�z���>�Vd���ZϮ�)?�V'����@[{⽈��N�՝cn ����k��w� �k-+o>2��X�e���R�f�'����t��NP��D�3�N����wBx!��<���w��� �,���Mf�)�w�\Y5�i��6����i�N��P���'�Y?����a��g�E;i3����D�R���>41���ݠ�V���}q��*�;��yS����{�(DCm��a	E'Ю��'�-K������I	��_!V2�$��PS���;��T,�H˼C�&K������ c�aǒ�Gaj�:V�֣��r�o��"�Y��6>�?0,T%���/W:�O֏��o&V�L;�W6��W�UΏ�:�r�:Ѿ0�\�&��N�ҢN�iW<U�Ǘ�^jk�e8ͧ�aΈ���hD�պ$����%G�0"͌��`;D �f[�γ�4��������$�v��AF�&���>^bn;�(������j�8E������=��iV��θ���d�KX�M8I�A�=���K��9 �D��V���6#��q����-���ݓn *�Ψ�_�/˩�c,6�.31����8�̭ڵ6���e�o�e�����:�T:���Hl�vXsej�`��eUe%�5�UeWQ��[���z��R��z��7��#���4�QG��qņ����}ؘ�����8w<�zܬu�`Q��<��Ǝ��8&9�][5y5sC&S�<�s��o��8��Y�����f��kֹ�%'��9�К��}F.�7!ڻ�h%hRM��c��N5ݞ��9\�z�o򖝁�\�	}�w�*p������ە'�mK����b����y�)u^c�j`�ȷv3*R�6�q-w5����~��p�fN�=i|����<���T�@��E�{����$��n�{`{�u�)�Y#�0<�n�HI�&������--;���j�FK@eW)R�����|�J�b����3�Lx�@X�B6��N�x��xj���|$MK���r�Nn���SO΃�1��/���361,9�4T�g$'N��s��A���#��~؊fud�^��Y���*��&��AQ��)�pi�U�p�����iu#j�ɿN!�sJK���&ّ|]&��d����x#U��V�Zt�5�@;�����;s��m	����U�����0�7�E���M��I.��%����1i�񝱿Y
�K�����(e4��O�XߎN�h�jƙ�\R����T�F���o�Y���%5���Z���N7��2���[ r�H+b` d���m��p����J�a�b������i�x̪�gw���Kh���i_Wg�cq/���b� ��f�hZf�xzd�v.8fH�L�ʩz���!��˴�|"y���
��[��Q$	G���&��� �朽��=_ԅ�:5X���������D6�v yᮛ�OK�u�.T��Ng�5�)�ZQ��J�룕��e���@K�%�y�xT��[t�|��}�>-GIHC�����n����8�h�BM����b���qŇq��O��j��EV~����ץp��'ۗ�v�}˩
u�p�����X��������c67��iC�������T� C�RO �S�������쌚_�@�16��s�%\�&����!45������2W�o�B��+x�b�&��J<@�}���#�	Y��׾��X�PO���o	~��y��n���,�K]%zR������^�� (A<~G��ۜ⊰�C��J�C[
H��Lj��U� Y���t�N�?��$5k�]��_��/B:����>_|��V��Gf(����k\�A�qU��?\�e2�s'J�Iz�Ɉ��#��9�}��|n 	j�R9�+��Z�'�b>�{&To�:Q`�z6�S0�鉲���GS-s\�&by�ms~H�T�z�S�����i�h�G@*[�>)��@ڼ�(�_:�x/��Q�h���M8W6�J4Jq	��߸�R�(�:tr���a'yP^���٭N�]֘����5�)�j�����!�ux��u+RR��P���|��⩃&r�@���9v��L�2&d����5o֍l4�U����j��+U�u��-eWC$�L&E8�����3T�<�����&㸫bq{�DA��0���Xekl}<}w�i�0[HD��2�	��u��������y�tpOΑݗ�7�YX��dU��`d�ŭm�a�|�<�!Y?9�F�����n$;LxG��r�(K�\�<�@H@A"J)�5&*�r���8��J�3�ݞ��ڴ��AML���E�8J�K�ӣ��ASt���B�����}a �D�D���ǒ���L�`bx�.��{�v����w�ڴ�?'����z���3�}���(�ݵ�Ñ!������ڼ>���Hd==�(�`��p�u�����}��~�`z{�]j =Ǝ����q�KO��r���Yԗ~��ML1������p(�K��=~,N��Wy��g�Ob#Uy�kp|ֿ��<U�6�l�`�*}o,��S;�[�z��3
���������_Z�/؋�T���Ê�ꠍXR:�\}��k<(����&���-�-ZXYف�7��|�6_��������z-wDd���2b���%��O��%�������q��&�{)�	�ђ-�Fnl�V�G�Z~	2��4��b1�л�e���,�BJ��З�.]Ӈ��Kɸ姠N����q� �i$�U�S&9ę�-��8�W,󜐞��� �qύ�K�=d�4k��lA	:N�|�����-Ҋ����mx��y]���WC��6x�:KO��UǨ�9J�E���Q)m��� �}y�����9����]���
�:�ͷ@����]J����	T�՟����{6ˀH��*$�ȇ�<@�
��_��X��z6�L߽N9�2Gcz'���azZ6���PY!�mǣ��,�/3��	 �]X�	8k��J�މ.�.��s�9�
_7뭚�r���븥NfTMEz�X�*semr�1��=�����by%5�z��� p{�cV���T�ی����O�@���t��A��A%۔�^�� �b��Z��u'��;�K7h����\�}8�_��(2!<�ĥwr���f�ф�&�g�#)������5�U�N�;�f�R�>��d^O���U!%.�Ah���PG�hfo�
.���??�t�)Bq�{�ԥ�1�/��V��;��J���e�T�yw}Gl���
Ӄ�%m�����f�&�~i�eƥ��P��x\�����۹S�ޏ�,�p�7�~�>;z��))3$��Q)�d[,5�<�}�*��K���h#ܨS9��̘�6����3ݷU�q��V*����>Q����B
�g�1�N������>��!�kC'��@G�t�k��;��u�/_Y��x�{M�1���^|7
O�U#1K�O)@��
�i�g�9�����a*ܺP��6Ŷ��g�xX��b̌�]�J_��V��Y�I� 䟻�⁹{E��o�����ǩrvK����!1��~�/9�]@�um}5;ְ-Ađ�.��~�����;����iN�K>0����S�$�>�$���Ѥ�ZaK*�F���w�!�˫sF���/�Q::$�v:�<��(�Zju�鋘��=p��`f}��%9��W<	/�+"�6�V��)lba�.r?[O쏥�X�-�B��ԤWQ�S�5�e���<��~nG���jG����[z�xm�A�	��=����+���ce�C�y ����X����:�7����/��!}'����jIFs~]()�����={��NHarU��%u�_Ɵ��ݴ�'�d�t���9#X^�]7f� '�_��;�xV��Nǰ��� ���]R�����ٰր�Xx_^�i,Ta��%��*��z[���r�AJZz�������w�p�
���|�	�|ᘠy�y%5/�cƃ���B���S�*vE�m�	�g�i�G�HE|��yJ g7'��rǋz����?����Fq�1EUP����{�n4�0ʄ͵�7B~����S�M?��@2Q�����}..Un�x�+4��V�#������a��Fܦh/EP?�_��"#�ɳ��zm{|W0�(,��3�.����lv����:�!�x��s|o��k)��p�7k�I�'�&�\e]��ٺe=�_��W�����wqe�a 7$�*�;���4{�k��Ȍ���� �b��B?G�oB�q�X(X��������/Q�VU����F��m6�zvd��f�x�4�ؚG-�[�裏ډ������Ԧ�%pI0^~�S:%A��Q�)~i����q���͌z&�r.����[��A���ߕ�{�p���$�Q��O�G�V��7h��v��ʯ�d"e�)����v{A���,4��"\k����G;��v�9�!�V@ĕ���H�0K�	��B!��@Z�<Eh7����;1�=׽�1{7wmT�A��i;�9���idGCrTȝ'B6m�-���|��/)ַ�cV��=�mP�o�b�5'����5
���i�{%���p����yH.:��/^�ŉ�����5Ps�H^�k�9:��I��ZBL�c�r����ɑ��d�1�y;�Č�.FG����`���@XՏ�{\�:�w> ��K��yO���w�����V !��~�O~����&���Q�/7�! =�P�� �� �,tYA�f�����P��/����� ��D��q@0hqstڻEU�D�
塼7���l��X�\)��=C��&JeX��&!���緁�<�����{����2�G(���&�9ޱ\^��ˏB��Q@*� Qt����JO�� |���-�w�z��{ࢩ1h
�V�_�ߐ���12��W����h�߬���-!-��f�dAqf�˔�%�t@-���x�*��6�&����2�0�B�4^M�Ë�T �XI��?`	� � z�v*�zjb���B�������yU�Zt�:�����RSP��eKs73O��̵�R'_�u?eDsw�$h9���#A�u�	��F�ܛ��ߗ���k�L��y�z�����+X97H�� �Y�c�#���������
����x{g+	�8�T�_� �#��+���<����^&F�*o���w���ꕋ���LK��xb��=[ӟY�1�(Db�������=Y�����+��DE��Y�Ч:3}�:�FT�JJXA���r�Ѓ�
mr�40❰j����O`���a}���J_�g��pyѓ���3�ZR��q��yS(����D���:K��s���[_F��YR/^�C�/,�\��N2��E���H�^��%��p�
T�z����l=P��Rdy�Pf�óu0#D]���#�-衉��5+|�g��QjJL��8��7$Ɋ��D+ƒ�t�A2�RM\��KI�{���p#yZ��Joe �ǆq�_�X�A�D*-�)YQG��˯��r�5��J��\U-�1�rL�[���~�'K+��0_��F���S3| ��֩@d��jޗy�*���_Q����mn!#.}�+��V���������(ّ���U��8��m�6�\���X���Ҽu%2�������g|�4h'j�jZ"�^	Zr��������{�v�Fx�f�����eTq�������0��C�R2��0}�x���3D�	]X�*�cS�)�Nt�7O]�A�� ��#d<\B��)�P�V�@���q�ma����ETG��!�5�♒0&����M��#�e៮���t���|�%Ж�#���=�n�(���Y���{pēIrX���,g[LNU�^��g�}���d��x�I�/��R�[���H�������a~E8�i��ԀQ)]��~C�����bE��n�U��Zf��ͺdq�μ~�R��x</��C��=s�e `��F�*VQa�v���&�ȃ=RZ絯�X.�R��f^t�ƭ��`	���$��ٰ7H�`Pg�J�-��8N���ą�6q@x<N@t��D�?v�i�'F4�4���ǒذ�����*�"=p��S��v�:.l[�a�sk�+��m����п���ԇ�(.@�MT�kN�+JS�5qFCPPSZ�j36�T�MZe.ɦ�(|�O���.g:|;�{X�{Yt�05&�a�b���xۊO�Օ#�a馿x˲ˉ�Fc���<Qx�[�V`��T�P-It ?���7���ԗz�5 k�����Q��cx�=y�;O\�6�������6�s\��Ϊ�=�7>�y�o��l�in��f���ބ�E\��I��G�!ј깈��Exf|���E0�9��ak�� Q%��C@��.v��º�f�E�D?{D� n ��u>�f��o7��b��Vo$�:����'(p,Xh#���FB����$����x>�ҝ��5�̀�)�_��������h~�7���I�\��<7�v��`L�g�޸� J�yRZ`рePb�ƌf�e�h���Ӌ"