��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~`P��(~K(���Ɔ���4!l<k�SC��h�%�8��wl
 Ѧ�>@��mY0q���/'��f�x`h�j�����:�n����B��3����ֹ�W�x6�<-d�����h��*W5�ZR���C(<�����Q�T<~�+8�4�<�}z��9v\��TrWk�Ym� ޾[8l]���wc� �lZڌ2C�����3(dH�҅'�w�]��]��W���"k�T;+|�$`�J��l�H�xa���JB�8qb�mr�d,��=y$ѯ[��zPJ[��
*��L݀�}�Pԙl3H���Î���UE5�B�h��[���i�ی��|{Լ�؉d�M��g�����TkBm@)-X8���ܗz	.�Ϫ:���:^11��|r�X�䶵��{�	�MT
��P���츅�W�ɝA+N��L�@�X�.�l5�W���~������!�����/D�G^a2%�,tɻ�Т��@��9oJ{[�L���+,�3��0ٚ#|�AĬ��͑��p2����krsv'vˬ�e���|��F�^P!�]K]O�`�K���ˠn!r�gD�aMI��2$�n&��I��E�]�:4
�1*���a�Հ��aq.��F�vlv&�$g��E�J���]J�c���횊�z���&�$�	a�<ԋ�V�bRab*��
"_u�o�à0x�K|~�o��;��v�)�"���a���Hj���{��v�;\��6�G�f�@b~O�iRa#!�I�ZuNW�4@�~�z X��t(Jl8��#���v�r�p�>���e5M�����������կ�&b��4�J��z�3����Xƻ�C$Wǝ��7F*�!⽽;���h��j�Vx�l���b��*�6e��<�
�e*nD������^�Q�O"�����H\�k��K\�����в�5�E�5E�T�֪ρ��_ ��LAs�,��	G��4��(g
�����G���cv�,:�n�c�u�|$o�4�P}i�I��v�(�B�ԡ��X������V�|s�e,���p4����U��'�UGB��Α[@���{�̈́S0o}��`4<��t0ӷv�r�E�Q:��i)̹P�\`O[IP�s:ۇ�����_�� ;�	��U���s��o�����)D}�U����߽�F�r\ι���|�2�6�ZsD�����a~�Yg�A<��#�G�[�?8�M6ܿDQ�\Xy��5��Q�džI���ȟf]���:�N�o=�^3�$ :9@��zs��F�������$nI�_���&bVὉ��t=�E�3�q�طA��\��yx�nk���쀹��W��9?�������o��tC)�w�*���H�� n֟s7Qp'R7�Z�mk���6�8��I&�����V��nѦzd��	�a���`�ĵɿ��F�ZE�o`��#���g���D�2pL(Q��[�o^�o��`�=�L��7��Kі�+�Q���TX�I(�LȌ��
6g�z��
��彦:p�Q\�)#jd�)g�9]�hm�u��Z����Q^v�~O����+��\F�a(����5,�zU�n{��%O����x��?��}��ޮ���eJ�m�7sU��R������!���{�nC���L	B�2D��b��&�Y�����mNY��M#H?�JsT�k3�Z+��"h	v.�%`2�N��9�E3�8�}\��V�On��;o���ۢ��ad�F���23"+�9ߨ�i_�^*�R���l�^��nYȀ,�OQ�+]�J*wC���M�h�����%���bDG�n��j���w=�풙ْ��Yr]I�����O6OJ��p�\)K�.I;�/i��u�
����d��[?�qLu�������<�&��Q&q58�B�,7d����;�wK9š�#9:_Gx0>�ni/�e^9��Ϩ�2|l(��q�{�s���jm��+l��x���0�5��03	��m�P�~�h�#�]<P|��ɨ�3����LӮ��ֵ�<NO�(�yΚ�y�]7%*��"��$3s�b�6��F�A	����
ձ���餇C�-%��[؝�fU�D2����l���cA�]�lΒ��{�y���OGOG��nm�5�ON�[@���R���>Z���~�����ym8$���T�w�3X���=9�����x�W#ɛ��ŋL����ہ��&:����n׼���"}x3��mwt��������� �!������A�R4c
�HIW�~�m��a�.Q���@]"w Լ�	��x�$l���0�M��y�L���~6�ش��s�0Vꋔ��t�1I�e����NCǵd��o�T�B)������$�&���г|�&e�jϓ��P��E��#`e�a�J��o�`��~r<�*)��Vk$St�H��G�I4��;I�����S�鼑r���C�'��z����%�c)�������k�c�H�xk��	�˂!����LLa/��"��tz�|��!\���EqY�����'J	0�̽�_R#)*���&�籢4wz/po�"_�b������Mky�����#�?3,��@�n`T��]q	vv��[g����Y4��@��C�37�, �y�a��� L7H#,����:�|�z�'�?-�#I�x=�&�%�Ƨ��{�d��)N��1��@����y�S)�Bx�Sל��*U������';��Ę��v�i��	����:�����4�(*�r�%�kђ�Yc�Ů/�x�	~�s��h�J���m��0Qي����<4O�LD�6�;��Cp��"/�9*������rc�=�7�N �UQ"j�5-�����h�֔���JoȢlo������1L��/�� �]?ં�� �
r�~`���^�r���t$?x�$����9�<,2g�{��s�aK:��t[�ɚ���b�lu*}?�̨f^� 0��ǽvE��wJ����T���X�VKu�9����Z�;7%��h���R��W�Rr�4���g8&/�(R;��"��{��h �R�"�}�>|� �]�S̟X|l��^�P�@��>j꓀�Ԇ`��)�,<d��� A�)�O|jA)Q����6b�$��!�g��M]�dT���*>��������/�Tʪ&	��ZH;��{HX|����of��֠�LE��q��H���(���3���=>��'6LLm�Ԟ����ƪ觾��9�ꙥ��w9��=:��>��no��J�,�S|��(��9l��
���='�iR�ğ���^�I7Q�����N]�=U��}���>?�����}
�ګ����hfC=i��+E��U6��>i�+�/*�`�:}�4�Q7n*	��z�����^���#{b����)H�cx�F~�>�p&�!D��> �F%�ua 4��ma�ݽ�v��Y9�N:��D} `�s=%dI0h��ȧ�X���v���H�c�n�M.���r�A��$����խ̓�A��5S����������#0H�]�̮�)�*�cXI'���;�g�K�SZ�g/��E�N�t9�W��stY��R7�a��g�`�p��Lئ.
Zt�C��{יU�vǱ�-��IDb�O�(10>�� �}5n�D�+l�Zz�z��LrS�Eڙ��L��H|J�կ�B*��b����c�{�	EF)KMKM��kZ/��}Gm�,P��]T}g��U;��O�����L��k�n��1s%e�G�����;�o��&�r��י��'lH�������Zy��Ӽ*O[����է��3D-y 
�:Id\��,}&p�4�yoء?�nZ��3�a��b��ٷ�k��#�~�1e�A\9B+�o�,��:���i�27jQ�$�;��U�A��C���Zŝs��,@���)+h�O! ���G(��������
ea�:E<�1'!FG��������k������1B�>�{C�tQ����� k�$�b�u�BJ��+�L3o��>�=�Ql��3v\vi>���9��]i�v�П�l�D��(�ؔ���mb������$1&j.��ے4� ���dl��ު%/1�$F��o
�_��0J��֖հQS���<��b`_F��"	�q�L��@#yZ�� {���{��JɊ��#�͸:��2��ퟣ~UU���J$����}�����o�˩U���<��D{���So-�uDp�~k,J�]�!�u�Tg��Iin��Ï��A��kk'׉�~�\�͂|@F��M�NJ}y*8M z���r���W��>[Ҫ��WJ��-<�<,`�T�k<ފ����&je�j`Z�_��O��'�T��Iˊ��Fԍ�QNM��|�J������~���4����+�x9��S���&�=��3��y�N�q"���$���������4IP����&�x�	q�BO��:�[>B(��h���g	`}OW ��F	D�5zPBt�$�O߰��'V	d��eIu��F��B����8N�Q�0+P�Uݞ��o�,0��ſ��9A������ϕV��y�k�H^ 5ƸgC��(�\�$�����H�	�2��>� b8FR��¶�CϽΌ�Y�v�� �*��Ipy�H��\ǯ�M�1��<[�mg�%��*_�/L��UTk\ev��q�HKjd�ut��3�.�5�M��䲳������O��p��u���(4�U48{���U�D�=ǩ�4,u�ԎM��L#�oʉTj�q~��LG������v����u�T��ߋ��� xB[��r�[�~����� �\��u^7�94��x�Ӄ�׃.�^�Lhac���v���)ֆϝ�xV'h�&)�P����<P�C�
h�w�����r%�-��*�`i#^����7U���e.�:�Y�h����������yYz�l�ٽw���0<R]�iۓ�+�=����h�VJ��[I����P�j��)���v���ˑ�:��cm.<n��ة% ͵:0�pu�+�0��(`6%nTruq�XEu0�1`[?�o��K����_�����t��ùA�ɽI�q�里zM&m���0S���E7�ƃ����e$#��G�N�} :2������A���}^ܣ)��:	{;���Y�{�7W\u*K�U)��C	������
�����y��`�	s#t�I|�P,y}Q=�Aph+v�o��0D��6�Tgo�>��.)���Eq�u.L�	�9��&����k+0^6�¶�	k����Q쟛#U���g(锖9Bد� �)#�ў[�=|�AC-A��~�(=����r�%ߔ���-,.��a�Ԙ9���4�xB�<{��&r|��z?�}�	�2��r-�|�>Zv���%_E�� -�7��[�I��f�XS�d$H�{�47Tv�����H솦e�{S�QAD��?V9���>��}`�������])?��&e�]�Yd�QH�
�W���%|  ֨i�*�%���?WKvX�&�O�
��?7̂#>�H��zKj�d���%ڗ?����H�Nh������X�sDd�@)�vc`B`ܔT���c��5�2��fR�yO%�6��_��M2����|g%��)��5+}9>�]ޝ~�>�s~K�`�5��ϕ� &#�|].����A��Co��
�W�^U���r8�}ԸRK�}��v4����:1Q��8�O��`��l�;4B�,��o]A�ܺI�rXҼ�zX�Y�ٿ��M>me!��Ĩ�����H��0C���V[��8��j��I���ڝ=�^�����
�. �O~�Օ(���8Ժb�%�T��8�:>���H)�T�=�)-d{SGa�F�b�sH1�����aڀA{�D~�;���y]�Lw��#vi>�9\��EV����،�������|';\J	c�����]D/U
��`���6����!�@�

������mq�����L���N ���
@�j����-�����6U���;<��Xl��s�g`�����(j%��Q�	��ލ��(�L����m�z�i|$��d;/M�W�b�\�g�:�r�<O��Gw�,rV%���2B��~��<Q>��N��-@�%��Ț�i��0��(�xCn��r*�t+C��q�w��6ϑz���w/�����`�/�&Lڥ��Gh�F�'	�e٪M�O}]<��'ڸ2����Ө��k�R������|'�I����ymSkB�(�[wn���H�)�0�գ�w�<ω����>ٺ���c�uj�-q�	|�V�� 2y��l ̌����P��2��\���$�uO�!L�Npa4�~�gd!�)�����`�����V�6�	?��
��ɽu��}o�9E:�9Ͻ����yi4�l��n`?�V1�[�����B�t�;="��*��EV�F�w4���df,�ĚCe����i�A���hJ�r��솥��x��>ΐ��=�Wa�chx�x�/�@	-
j&��V�Ph�YdH\�}>=����:�6��O0��Dh�u��=�k��5.1s7��U���?�#��E����	l�G[|lSqe8���Ȁ��%e�W���TfKqd�
���-��/�g� F3��H|<���[E߂\kw�X�6R<��)J<�{Ę= ��
į�δ�Sg0 ��?��L������yȇnB��V
er���}�fQ ���Ay� ��w���Ϳ�Q�-}�d���]��l�{r`ޚ�1Y�IҤ���31��S���·ȳ�J�����Tqc�#��9�F��B{_AIS�
�O���Q��c�[-

�&�4�˩���,���^�nQS�8h�5�����nF��
�3CA���f��_-�H6�R�zjQ2�#���y)�C��9�3�B�D���jśT����a�����c���]�	}�w�Q_&�=:��}�z=ri�b�]H%H߆���׊��Ū^_ <10ݔU�+�Ð��<�O�P��_T���S���9�� Pb��nt��ׂ�&� V�{1�.��nR9�wy�"=C2c�(�&�@�\�%��ߢ
�v��ܢ8���j0�f^�S�L�4<�O�b����r�S�<�f�Q��w���3�ovj�?����\xv�;g	r$-�y�\���-�MM�ŝ)idp����Q��az����t��)w]�Lt��l"�a>��='K��@�K}��	J�9���FN��߬��L�)�eܒcS�q�� P�Q.!x**5����:H;��7&#e9�',w�(�ٸSj��;2v�edW����|�&\SXl=-\���.J����o��_�����E}=�x���l����I�L�~@o�e$1���/6�D��}3�b�8���wM��f�_uqp�r/5$���'�W�l�0�{?�,�8��X�؋�R��A�xl�ݱ��(��:(,��(��~Q�c���֜�ɍݏ='���,	7m���=�SĘ�|2�l�"M�F4Y���,OpHxGA4�/���z'�f�vN�9�;�6��iG�U�0�AFޖ8�
�g� ���!�nekt�~m@�p�h5(���IiA��«4���aO3+���7)�r�G�"���Z6?������6� V�M&s.�f�_j�p��X����uSHO�����l~�-��[i�q3Fi���*�W�@�_3\�n��!��Υ0=9[w�����f�������}�����xs�-TQ��w]����W:I�F&]sn�8qgp��Ǉ@q`�q[uOx�d��P�	��117R�9�7׌����њ�3
@t�C����X⊴c�f��Ts����<�o��pw�?? ��l-3�23X��a�f��N�C>��U��"l�߯�k���+@����s����Aup�>ҫ�҉�B������1\�eZ1�u'm��9X�s ��ObO2L�����������8���t��`
ʤՙi&b^��YO�����^?ƅ�tD�tU���6�5�^�ؓ	p�|f$xotU�dހ�����n�n��%ps��N��G((�\��Y��,�t���\&�e����6|�=�̬y������!}���X��Y!�qQ����`�Ku��@F�RU@΅��iP���r��Y�vy�9a���pmX�nOb��D�����`ʕ������f��B>h0�vC�LX�����3�X�k%]/����������M#��D��p�09��"��K������;����W?R�� �8�ř;���cn�r��)ӛ�����R���:C&:3>�|W��!�J���5u��ɂ_��:iģ"|n�%���Ȍ-���T�_jg��i��[���*�T�-eAB�@X$$�۞� �������^��:r�Ʒ��mƗI�չ7�!"����&�dm���_l���'�J;��7��)2��]w��*��^q�&_�m�!��?�f�|0��E~�׉����	��4@���>����xxeh/"kΥ��ĒP��c�ܟ�f7&�����W%���ćc���npD�����Q�ա��G����Ş�Z7B��m����䃲aÉƸ7�!5<%Q��K�Q;�����		����3�@х����I���R5��N�u�]%:#)�a}�i������ �'�`1ҍ4tʲz#�� %��;��-����,�

��jS=�\f���)9q���<�e_r���҇`��ǎ�_��HX&�b��:���S����`���@�r��J�[2_tO���j��I�p�`�@��+D�ZzB4�B��T@�yփ�� hY���1e4�j��@�hр��S��d#��J��U���t�J3��)��l�kш�e{�yѓo=�J�ǝ~��OAqGAN��<GR�W^�H��@�FE����(L����3�-�����Τ����b�2f��p���RafK- Y-8ј�����Ӹ�إ�u������õH�E�!y���ycWO�F^��1��!����m"=^B�j-�� ("\���ɣ�� :����x?oT�#��#���L:&�����*9�m�Ԟ-�!��o��ѤbDf�H����;45�[F�������>Ш�0l���ٖ�TC��-��-͉�?�JX0�X�6�{��w�\��p{��M�f�8��Xf��>x�z �+]����Ykݾ�9Z3����׉�xu�@�B�zZ.]�H��ú�á�[�u {d�]�baW��C梠ѩ � .a�)`g֛��ٳ&a�s���I�GPv5C��yO�'�juG�t_���B.z�G�7z���o�3_oYi�#beEt*U����P��2��)�$�#$�͗Tx8��4�aV�D�di�{�k���m��f���#7Az1P����v�q14�I�Ʈĵm��.z�={&��F �C��	�nS��Ek��
Mi& �,�� N֤�����+�%�5���쟾�f�D��]�<���\wS&�w�K^w˂9<�RQ�p�y7��:W��k�r�����v��t5j_��(���*����� ��[�dE�+`�4>v?̂9I$],���x����M���|a��3\%H5̫5���t] ���7��aK�pF���Pu��<1��Q�֩��i�5K�dD/�(��D,-i?�HH�wS�T�w����o���1\�.�`b��I6~s"NS��<�
:B�(1;�3�'I��pY?��;�~����(2�>�N�K�����K�y�B3O �^;�]�}����I4�|��N5�BAx��������|��2�� �1�����Vk���ݑ�+P����$��!��/��xI�֘�t<�]n/�GM�%'��9�>���y�VZ�!�y�I�U��NC�do`�b��P���)� (�^���Dϐz�j#\���
��vJ����u�%�O�ڝ������Q�wy潵5\6u5Y�����{�t<h,�oaE{����>�҈C�w{}��_�k*h���9�r��kDw��#Ά�5{{{���k��3��'�3��Ue"CD��(p�V	�Xwz�GزX�|"�A�| ���3���tw�)��x����,&tA+�V+n��ye|BT�:�aBp��G�"��iB-y��6�u����H�뉟}�-�8L�d��#GX��ƿdpzN��?�G���'��׷�k����e�q�K���P�X���ibt���RD�f�������K��+`���nتp���[6��0���U�i�J��/�0�lq�?�X�$����0������.�3�@X�LY��́�����䘽�5i2i�z�B�c�9c��5������,����>'p.ٺ���<P��}z;�/�n��	��an�o�A Ө~���BD�@N�Cm	~�L��+T,�9�#�ɛ��X��W�o�q�=�ڼ�����������}��*䯛�o��pi��q��S)�Z����j<h���\�����+ʤǨ�8?�Qؐ����=�:z<v��
��i3X O���w:���@��K}J�a�C���] �bFK/��G�%݀����\�q��ܨ'� q�c �X��pl9gOE|���� e�(�p�h�\���2߾۟F���v�E�\�Ir�E."I��I;&�齉��0Xԛ�7��Fr�|��)b�`0�^8�P�<?B���LD�U`�8�����rä��+���l3��1(���.wj�H 	�ǻ"T]�u����6n�`L�iÅ3��������{R=Qu�8?t��[���Y�$.>���n���k�~l_�8�7�
�,Qm���]ҵ�R(�lskGB�ڳ���6	;�^d�b�/)��r�n��@���������%0���6`I� �yp��x�S��+R�H�θG��,�SM�SaP��(��%�J ��$���^�c�f-GC�c};�1Q)ڗPd�i�Ht�.B�8-�aF�0}�q�ݿ��`�;��[�A��*�@����2�]9��J׮�!�<�����2n�� �8�����K���I�inb�L�yu������	T&�b��������YgH:S	��ޅ�:P3b =������:{t�n<��Bd�25z�A�m�F9�(�`��������q�U�*����%�3��i ��$����;��@��иr\���Ö.��EN�T_�ĳ��7�ݪ�� ��Z��"ZQT����}��%�( ��W߀^^�f.��?\5���8�er����YOT�@.l�E,��c� 2ɕ$V7^�J���
��k���t���#�&����g���jJܘ�)̑��J� ~.��������I�a_Œ'��
�|"|u�(�MdڬZ~�'����[W�˿Ǒ��Ъ^ؼ���!�?�R�_ݲe�~�ES?������\��Pb�%���~�\�͛T1���_z��#t�v�M�nR���qF�ϵ����Z��F�\�yC�m����-��T`\�����}��3;�}��"�Ћr�u���+�]�]� �Κ�2A=$QM`si���Ao�i�4���>Z��*%�ٴ�Ʋ�i�B��#l%5�+�z�ǔ��a߽�@>iw=C�M-�鹁Q5&����۠7Ȏ�Ժ\S ��+h�Τ�گ��|=��t>TJ����~3Q黙;%��'
l�Ө��5��1�f�<z�(rֲ�;3,��`���'N�S���Wn6ﮭ������Pc�B�=��w��s-:90�Ľ�]@|θ6.��T�DE�_���'��� ��q�4PWf���c�@,��y�.�@���ۚ3Xf̅��OeL)GS���z07�%L�S��H�}�������~���p>�\���f�+���}���,w��L]^)2��[y
�Gy�@#���K�������rE$��>ŀԠ)�(�㒈��e�8�~�p>s��<!Z�r��YtCd��_(����ܰ4%j�7�?�>\�ms�vz%Y10�{�4zl�#���%%���,{��h:w7���*l��x��'$�.�a������rq�"v̥墷1�3���1P%�F��2����E�@�F�����Y4�l}�U2$�/5[I\e������-$7E9�ɝtx��q�rU�+��֔GM!���n\���s��CwD��DJ�+����0��*�H��������1،p�V���'(�O�1��Dfi<�=�XF�9��a,j�8jp��tٔ�+��)RTv�t�*�tM��C?��v���d~�C	oپ�q�ُ�]a(;�4S��~����6T�p�/�S���Z�1(�_C/���S��7�m�J�BJ0߲�9 9.�e_7��D�D;駓�{~�����Q�X�*���>������p;(Uy�k�����`����.�al������2XK:��l�i�>� �H%z����kG��=,l�����S�0�R\*��_�|�! x�L�:,�i�����g�d/�Q�s�p���#�Οrd��ЕAz�::�u1-'�v|x��/-@��[)���qc�f�)�0z�܀=O�� r�-�7�˪#�"^eex;,�ciЪ�`n$�K�l��'�i��6 �0���?DF�@��d+���o�L����;��Z26)V�%	�Z�X�'���8;�7�Y�_3�!`���H�����
�=����* �O�OR.�ȍa_n�m��