��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����z'H0-R��Ò\�A�֙'�����?��c��_�)��Ӌ��	��VN�>�ZOD�h��-@��y�e&v[Q%�,@hi�_�o���n���\�oտ�jX�Nw�<��0|�b�Bs��� ��d���~�-N�s��G�
\
��vR^UkA ��g��Ｙ�;!�P`�z+/Z(�������(o��&O8�R��(�DA
��8�ԕ� ?���Jv��Sψ({����a�1i�	�qF��U����7��� (�j�d��T�|K8RZ����M���Zl��E?<��X��@i�N�.���jƨ�[ ~l-Ƃ��`
�[�DEg�ɉ���O	[����ծs���<��ȰE��F�l�O�	�e��O� �c���V
7�@ux-@��HOV5i?�
@��w���Й�k����Q��f2oQ�b����V��jYIǶ��J]c$m�W�R}��_

,�I �Ʈ|,H�x�^�*�li���燏޴�[A��O��*�9�a���Hbm�K���|t�R�\�[M��$?=���|�R����G `����h���1K�|׹��7��V�B�9�����PX�^v�$�'�Oq蕥?��$�F�����Q3S���ȲFX�����~'�KT ew���R!�OK�ON��gM�����{2�����L	0+Z�#S��m�'�>�<1xGK��V_ ;+h�v��ޤ[�}����a�<��V�'��2c�A�n�P���mrW^kC}`8K�6����f@��O��'(hc���o�aij��H�rv�� ;�}V�D����h�YY�1k��� Hdd҇S�%�\Y/�Ay��n�h����T�3�H�j#U�H�'g�r'ZG�C\�gۭ.��廤��]z��c�Ҵ����hK^����V[]e.�}<+J�t������O�����)��sRk�A�
dy� �#�!f�G-��|@ji* ۙj7��t��h�)g��%�����2m�Y�s7�Lt"�E�������-�Gb�p���1�&R���2�.{f�:Ӎ�D���0r���lя�'G6~~��,^�>��O��� �??w����C�9��W�d_m��!�_I���֭�T�ڊ��Q�oK�f��*�����[,���̽=���b�P��t��#���Lr ���k��Q �c�Z�!ȓ+��|�V�ܮ=(^��pO��v��ˀfA�Q[�\tq���I���V"�LI�O����^ᪧ_f�d[7��y]��[��n_pC�@���*�6Ƙ�^��Ln��í�'�@����e��V��['��B��pzLcp�n���n�����x��٤�PY�c�j	��ma1t�6a k$�ܜ\�ؤ��E��z����D/������K����W��0�C�Pi�_�xlT(��������)�؎B��.��@��[Cn5`����ٶ�5��2ő�]�p� ��8��q@���/�H����5�YM_���ϮD�2�ޙ3���^����0�\D�yt6��"�B�9�dj�l!����A�b68���B��m�<�Gy�+u�,��P3w�U�����x�ej�-��JL8�Ĕ�-� �2�^��[���S0|h�˷�$���a|���!�α�t_��Tǃ>�%ŤVcJ~GV(u�����Q�h��6��#A4
sC� ۙ��D$��@ y��=?��7Wn��!5vA3�YD��yi�v���6�Ox�0T4�I�@y�9�-����Mo��PC�Tw�A�T��
)%�󱠊��Ώ� ,3=[� ���>�^m�Y����:1�n�k��-SS7w4naS�Q����Դ�T��Y��yi/d(K1�F������¹x�@�5n��!�Q�عFT�ݸ��#�0Z%7u����K�K*~�OԌ�P��ɏyU��7~���T��w�"O���?�tK���_|�EӒ�O�E'��ǎ��i$�V���%�p�dA�k+���:9ͅ�+;���o��JhHcޚ~���47b���I�V�H�S�zf�&�z�EÝ��'���T��y^a������:�H��Mrk:Q�L��g1�e��_��{:��c�G���	Wq�Z���ce��-�4bd8��+8�y�#&}h�������yS���!Ta�E�Յ+q�+ q��Q4�#n[Ў:5'��O�[}�V�~��y�nwp���X�1���%V���pq�h�����G����m��pl[��r/�ț-�� �=��-M;"���_t2oC�]���x܈��\����1Vd�R��{,(ʰ;�x�%��yS����a��t��{%�nL_+����A� ~������"���c�|͌��D�l�S:�y�Onn��
�a��z���<X4��
D���TL�"��E�e(F�kq��l�?�s�����v�ϬЕ�$�EEj4��S_��*��2��n����=��Q%��VLx5��o>�LR�N&��v�w�T�z`F��]mG��#wMB�I|�ܒ����F@��}E�̹h�%N���i�,I��R̀�X�^ɝ�h{�D�-ly85��_r�SA��aW]��S�L���^+�da;^[��$Y��/l�����	���^����\<f���_�����Q"�w}��"�d��qC��zqޟ�Sa�xۮ�v*8��lf�/ ��D<����Y��3Ho��BQ��CF�J��4���	�m0/����b���?�wo�;�p�މ@�!�l=��"`zV���Tmޏ�iH�)��A �j��UJ���v�%�R�"a�S=�c)t���Y��y��O@PjW�3�nӖx�l"�E��$)�#'��%�?+��&�����^+�tC����O���������~�p'M&W��-�<}�ל�¸D�fa0�Ժ�tŀ����A�d#%õJ�VQ�ؘ
i���M��:����	�"&Y�q�w�B���@�-��b�LT�-�R%%�%���"�&�(����W�ʈX<�����2�x'��8�C���c�^�2�f�h�Z���+���H
�����E�{U�g-V�_�\��ԭ������~��{��������}z5�w�����2�OM[�z�1�:AO�sOǐ�O�#pXqI��xw��丼�a��w@u`�aí�.3�^Ը����}rl��9�:%����'����'��5��	d�oh $w�d���X�U�&�bۃWO�w���[(Fd�y�����,6x�!�n`{W�a�x�
���~|)h��a$��p׆�Ⱥ�%��JΞ ��Qc.�+R��
M�J$�gkO��
�=@+���_� �e���(�\���u�]��베:p
�U*g\������&�-E�L�'b�3���"�H���%̯ �UV�'� cr�6�u"�hW+��@� ����E>��ZV��`y�e(ӧue���Ad��j+�4 �و���E�fp{�	���c�Gi�z�X 8�R�<�+���<��X��W�h`��;2��i�b]���m���C��Cel���~\כJ��Ǽ������� �8�'9�[k�sW�g��������ۼ��H��m���!K��π���c���D�i=)�i7�HK���ŗ�����p��θ�^{�,�	� hUֹ���u���k##�<��q���'��q��5���ܼ��#���N'�~��͝D�'kY����I�,ܫ1I��fk�T�p������vG�L�t]��@w�cH�!s��a)� ����m��B44�Ap^�u�bE�E�Y��+s�ÿu�X�@�&B-�s��_:�ݶUW�פb����p�K��z�����9�}��8a��jV`]��5T��&����Д������<�G5�VI��J��� !N/���̦-E�K�RG[�=�J�%vD�zl��r��Yщ��_���	�AM'f���{�w"�~C~`����v��ָ���W!���|
v]d���)C�&���j7���0|.���m�)�,�Zo����+������)�	���GU��<l2��"S�.�,L�Y�Gy�����l�B@}�5�0Lͤw^e�	nү��b'���9�n����1p�-<�A~;
���?�D���6�#^�0�z?�NYbI�Q	G@��n����w� D���z�`��{���ؘ`7�<�0��[^qD5�����z� I��|�P_֭~�Q�C>/�BZU�X߱�7���Be�AD$Es���9���(�����%�=�b�Gi���$@J�k��t����(�_��ȃ����� �T-�7���"��Pd7�vX��Þ�L��L�Z���;�u�}L�F��M��{H�g��N �d�rנ!X7j耆L���������_E7E��QQ�>���Y.����Y��D$�L�(�o����Q(�93��X�9���X��k3�7�V�΋�;�`�2Y�P�X8�Ccj����x�ɨ�p�8����[�f1���r�K��3I�QP� ��x:RO�V�U��C�\xUV��m�)�U���~�SR/:�_ ��&��9��8�C�� u��
De�§�x�T��4)����G�BʘWt�
J%Y@�"|�B�[���V����H�G��>
1P�i�hjD����*�Hڧ� I��-��Zi�(#Ò�6�J��������� ����2��!��Z��`L�|��'�)T��AMڜu�� J0�ckhdr(IJ�
T?ߢ�P���'#������G�<
�L*�MBV-�O˟��\���>���g��p~�c�츴�߅��#�Mb��u����Il�8�-�۰�s�S�tU�Y�e��w���c�3���ϞZ�^��w��m)�	��7/��T��/
�J*�+h�ebpY#p:���51ó��b{���)ü,*�����bj�q���,�e��no�M��L�^J7�'yUT}��~��x�S�����`���%.�>�E�c�N�B������=B�. ܰ���?��dDp+3[P�)���m"�|�QX^� c�������Oa{��V1W�&�O�F�iQk��o��)�'���T|�ԓ��P��P�������(��\���42Km�I`��]L,�������'P[ �KT7�9V(��d�^��w�a��Ot(Oe�Y�B@%q�pTZj�&'�c8���̐�IӬt����cLO5�?�Ə76~�Z�FA�/Ѣ|d��
�L����pg6��㱈����7B�Iެ?�O��QU>���krO9f����C<�k
%�w-�Z#^���L�A&�o�z��>^�ah�+�O����K����a��җn�z�nr���x���s���&���F1��󋀕�kE���a����BQRܱd��B)n9e
$s`���Ԝ��N+�3�(�|�8oU��J�ɕ;:]�m+HI
�U��{<�ǲ��}
��~��D�'�m�DPO���z.��ke	��($
lp[4�dbl2J�r����M�ۭ+�ę����X�O0cma?g�J���:û�煣���~Ǖ�ڹ���kPD}!Y���RRQLx���M�h��;���_6^�,�x�ѿ�S���ߴ"�֤xU��/��������v��Ǻ�&����U~P�N�8��xy���i]Gu�4u�_ۣ����MG��(��a�I7�Hkj&�n4����j����� 4q��"o4�.]���ݡ�xlUPD�'�1s�s_�7�]���Ծa��T�
y�]���K'������
w��D	O�^a��w�W�*,���^���!N�UZ(�Gf3'�S�Y�����@p@6+���������J��-�u���vx��y�_�e�Pr�QB
��cR�ّ�	�~
���_<�!+~�������:�a�y�8����w���