��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:��������uA��@��y���<����xDET>��W�����C%�=U����3v���hj��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��pSv@1�{=�\��c!?Ƨ�'�G��q�2�4s�_�B��W[��Iz�ߩ�_\���`G���}���}�7ү��-��T�'�kf B=ٰ��R���l�ta�x�RC!�*aq�޻+�z�)ƪ�!}P ��w�p�9u 굳����w3@�j������ʢ�u�"c�=Ǯ�1W�xCM��Cz~���/�W��(X-x��3��rW��|�BYiC����O�NZ��Q�����2�*����Q^�&�O+ �/�Gb����@}�;g���O8�������U߅r}�Ǎ���˪Xt ˈR��H����<s�-�$�]5%�iS-��~tO��V�=��k�uZ^]�R|d�k^w{���܈�kR�����C�r�v�ja�M�C���uE\��w��9I�D0~u[NHC�3����֦�cm{��x���8'�d�ج�̷��B��4i��-4���tSl�i�U
"g7��^��5�G�g�?��4�ר������a1�Z�<�5T�Z�F	�/Kѹ����U�A��IyNR[�8�p��%��|y����>�3��J�����:��Ӝ� "c�G4������0 �+h��/^��LED�x?\L5�j����~XGǹ�&*�ݯv�p�-W��RLFp��(<-�k6��^\o�Pz`+��m�V��������]��͠f�Ͱ�r�!�A�zPNb�ߺp/j
�,Ɗ�W��Dj���Ş���Y�r�*!h*�\�X�L�dU1ejy΀Oگ���R9���(:�zu^���ޖv�#��] ��U��+���0������������P�C"��Hc���u��jO� �B	ACo�a6����x����,�Q	f'Q�����4�Kv�2������x�w��+�t�8�"�m�A4Q:uW�%4ռ'��f_ 9�:����I��=�V�����������v��h�?�O�/�u���9�Mq�&�mS.����#N	����++�j�+�/E��n@�hw��x�.�v-t/��1QfM:���ϑI`�6�O�pV����p���5���|/�׈4-�f���~�i	�CY��Vu�������W4�*m��B��3zQ�/ Q��,r���!�fo�׻n��e'й��~R⨜_�� �:�$�Jf���F�jO,㸩�e��-0�߰��^�Ρ�T۳�B��o��6���h�����9)D9��E~�}��PJ<� -z_�?_�Mw��ӈ��ikѴ������7�\���o���U���D���h�x��ه(�b�Ի�w��Ǭ����tX�Jo��F�y�e�p�!�%*��l�6�͋$V��ӿ�m���Q�P/^h�O����6\�2,}��5�o��$��s0�r��F����m+~:��wQ��4��0���fp��A�hrʝ�![�����~� ����.�=Zn/��+�R�UPl]�����ߠ'����>�∖��ΜYu-�����-|�-n��B̐!�%�M�R(����B;�i�tn�*����#�BJ�T���F	|�0�Y�Gb�&�gv�A������A�	qH�U�xE��?ja��0����[]���ub��mk�P�JH��H�=i]dw/���հ(�F�+~�g����cme�t�x��mos�
���^$0أ�f��2�P,>�{!r�y����K�t_������,���Zy�\[$8�E!����F�E
���u7�Zx�-�ܸ��n�)�	ޟ>M�t.��4:�3-��\���-x�1*E��Q�9O����e�p`"���|P�f��� IT \���7�x��J1ZNQf��Onڼ�P����Q)�1��ȳu�
��ux���9�~�D
IEʣ9����*F�v�P�Ԃ]��z�l����@�b90�>oςM� )���7}y[��S?���aQt&�,�Sݛ�t�i^��{��΄o7%���Ǡ����W���Q>�����v��2�Q�y,wᢎ��\������	z���M�)����e*V'`|�[��u�z�U!��
�O�-���0��,bm;
M������C����Rp��c�و���"�����A�qPʝ�Rqw��[���THꈉ:2d���ŶSu]Ή�/PiߒS#��(�>��k�.�f�zmE��7�"��b�=��$�m�=}�a�$Z���Mڶ�'�)���.��#�%HԐ�s��NYOLpCϘn�����0��h��iL�����|��a�$�A��ZP	2UAABC����ヺ�ǋ�:����ۈ�:҃�e���N�d�m�TGd�X$Eخ�<�D��'5�/X��m=�Æd�����.����;e��U ?�͔��(���4+?Dh=�Xy�]��5���6ޖ��t,�!n�7�q�kB�3NBm�k䬚�T�������m��xw��g�K>*���?9��:��s�����.X����Ux���	�w!�S�X�@ʲ��䅏.���+�+/H/�mQ�/�|ɉ}�x�X�(�L�� #�,����#���������5s7ֵ\����!�e ד�H��t�ס�aJ܆+�ڀ�\z��}����׏#R,ݜP]8I��]o�
�㊜�XS4��S��Ⓨvb��*.]���� �������mj��f6N◨%�w=�:hV=k�#�O�f����o`v�<�S���$��m���q�zu�˙���!�N��u��S�ā�r��w��쭴��#fQ�AA�	�렁��t3�����UA�Kk�T�H���tF��.( axO)��v�⫚s�i�G���
-e"� x��a�L��I	rA���n0�_�I�m.	����Y#��XD�Ԁ1ϡ�q` �IEN��4��,�/M�����gkP�:{ň5���|H�F9��F�L4覵�)��}Ċ�E3������t(g�'���]d[q,#a����)"{�[������Tm�Ə�R�M#����qwhJ��t�ūx©
(+-����B��A�HƲR��A��-�<�<�Xʡ�A���Y��1D�~y��-�����f�{�*�A4#U��YA���,@����\���ԫZ*Q�	ف�;�����5 ���s�lH�	x�/��z4;m�Xvσg�p}+��
1�5��0�i�OW���ިok�7Nc�-d