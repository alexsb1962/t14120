��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~}:��<#����OY��ru.�!Cn���������]h��j�8|M�)��W�V4Ek�
}�SA,�ȱ�o_�w����p�~����`����ܷ�;�<� �����Z���òf��ۓ��)�O�Z�{F�3���_���M���s+�+{@�>"l>JK�(�r�u�����<JT�]���0�M��0�T�iu���ˮ�_�*T��h�)�%��g^�f��N��DQ\��j	��8�m�x=¾���Buee�?��E�c�lO�B(�<�2f�/���E���+jr1�Cq�#<܍����J��Ou�\��GPk.rD�UK�ش��Z��O
��r��3�Ҽ�W�ڎ�t���&�̣�vɌ[���+eT@@"�<�Q|ƈ1���Ip��1�<��fQ�l����E����l�	�Dz�L���.�~�^�)S�'Y�%JG�E����<�m�5�s�f#��s�����z�'�
�3هݽ�/�����9�P��]�[����\��5W��d{ԩQ+�,��v��4�r�ׅ���V/<�'�$V�_����u�m��K05?ޙ�zh�:��Xc�.�����b`��)��ة���	l���� ���EZ��`c��}���a�l�p�adcLWN�U�ZxQ
`���e�~��<N 5��ZT�z\���M�Y��\�������H�s�>�Ny[9�xd$x�sݮ!Y=�r�GF���P�B0����4�h�t�J�Q��<Z��벘;�o���e$�ua���KXAe��0�Z0-GAo<�A<��X��d�2�d;�%]a�l���1p���hɐ��t��	6�j�(�S�`�/��4���WZ�+��׈�~y��~��: �S厏�nE��>v�d>mrb>���G�$g��^��j�}ꁸ8��\o���ZLmM+���Zڑ�un��3�?��Z���]2�����8I���&�~u���=�b);9���Gn����wGm�p�T�(�͞���+#cSd��B�/���'��e�E�yl�>��F�H� ����hTDY7T�nS�kK�� �jCVA���[�IW,������^ e١��F��{�D)=/���Y`�d�R+,��L,��@���>�T}�P�����s{�&������H��V+|<��Waxu^�f�d��g�FQ���s4�39����%CS)�Yy%[\�����77VI*�1���:�D���E*�_^]7��hf@���[UZ�o��dGRv؍�b�pp)X�5'��#"��2R��?BO@�Dkٛ����p32Z�0l�����+�A;��3�#���ͬf4ӧ�աo��/A��ٯZ��-���҃i����;$��SZt�e$r>.��᰼����/�J�+p{����-�-U 83�Y������k�F���B������y���F�]�]��	��+�LT{,N�P��07���>��������zՙ�s!�׿���@�����P%TiBm�T��lu}h
�Ƨ�XB1L�]3�2���t؄ң�<9]g��J��y&*�5{U���P���
��-º�ҍ�lUȈ3�! G[�����������8>�$z�
hx�38Oٌ�����8�	p�պ�l���&�Ƈ���C�F�����f�ź��	����6���n@��8�/���s���5�V��r+�UA��� ���/M�vZG�B�;$h�^@
�#��b{<��rkwE�_�]�8�1��&��a�/���F��� jI��2��j�`����V	<��t��@&�y��Ǝ29GTtW�=�v�f�H0�)ݗ�W�|Y�.�-FLL���՟6}>�i�Zދ�5|\X���<44d�$P��g��P2��`^�W|�;�M������Da���t���"��b H���7��"6���6
���py��׀��6�OF�O�T�g
�����q����<�P,E-�_�Ʊ(f�-��l��O�M�,�|Ƃ{	<��d"Ud3�\�ƙ�ۈ�Qc��Չ�a��A�/�g��Ҙv�F6NX��C~/���9�m�I���v���b��Y��6���9I	�5�A#�<�oA�D��B;����L�R@ڳ�f�fW�.���J�M�����W����`�M�X1��+���K;��W[�4��0�@G���?Y�!oP�)��ӟ�W�ؙ�S	)C_d���xt�dp��%�N]���9@
����m���B&����qٸ���n���IJp�f>�(�c������?F�<B��A|߹�����>;	�IH���-!{�f<Hh 1aH�wO23�����>H훋}.N8��Q��0��	]�}�����f��	�^NX����o�ySQǏx�^5`r��e�������].z<t}5�Qd���a ��z!Nj�"'֘)�������ǧ'��gR���P���Ή+�I��f��!?�������9?T�,���zw�&�6p:����Z�5��D)50���][2���{�Z{�����^� ����U�ah�B���y{�'����|dky�Yi'�ő�AI��o��82���fꃭ��==��V�,8G�Ba�(�O�ː(z��a�z��i���p�J��������Z	�H�8��j�	��9�&:̛z!�gW��E�X��t:S4��!<!���SE2a�x�?���7�� ���La�>�ZS�EّC7_
� �a��JH��Rã��s$��%�=�(�����4I��԰�^��N�ܯƎn81U)%�{�v}a}�v�<�L��ᡣ$� �p�� Ԯ�}�<K���SE�B3��_�|m
���S��baQ�*���������dO[y�=+)�-SbZ(�~�a�%�d� ��xS�<��m�__���2HaW�m���I�,{8�,��Lh���G���)��a�ۮ�=������/mhk'��*��/�S��DeH:�AY�;��Hc0g��+��\��8J�l��[��G��a�X�_f[onG���
/�y�s�ь��K�!\�� �i(�<�a���\�n�s���FԢ�LJ6��5z�V���Ƅ�߇K�3G?7�俚[�v�x��!8X�؛:Vm�Ǭ�{��l�����ܰ�؍�L �y�fnb�jй��_��h]���R�ό��Xa�-����qx��I[��:/��1�����{b�GJ^�}��W���vR��^7��w��]����͊�|F��|��z7fi���O�d�d��?2F���&ߠ�e��3�5����[��3����$�`��L�X����Փkm`����n�����[0�E���)�����q`�	��&3�Ț�L�LA��u��!]iz���=�#���A�]�[E�v=��3���Ɩ΀�9������H]�r�[�00<�����,)���M0�����H��r�BVL ��!�'��,r�{F�
 ��ep����/>_uE9ُ�At����s��P���O�s 8��)�p��u[�H�p2p�ۯ1��0���'�C����`�&^��B��\�yi���)����ʹ����y�@)u�Ȧ��3�9�,�ZU1zI�5�P:��KMp����@��y\���a�iFg�z�7�8U���e��}�)�"���|2�s���a�>8u*��&D�K����"��
�(R��֟	��T�cT�}jO �1�{�7�)ci��%It���Q�yҞEA��^Mffo%)x�ыQQ�5m��k/�Sbj�������f3!��Te��=k�	1H��~ƃm�^~I�L����Ĥ�b2���U�E������}�w���!���շ�2Wn���>�7K0�t
�=�v��{�K!�b^�0X@�<QéSsr���%�W�iM�<��^�������M��&��n���hpt�����ތ������(=�h�[M��}{�q䃷�Z����Zw��l={��vUj?Nn�)G�� ٿ��D�}֌O�����w����{Ĳ��AD$��z��%%�2K;x��?:�]�F��_�}
���,a�ULk7��w�n�� �y=��r{��c*+���e�!�;eH3��2o�1W��m�R\����/���I����A�m靫8۞"�W��/(l���.�����i���Fu�v+��Q��,ǔ�)�3AI���$�M�u�tyŅ���V	�vU���/�r2�Q#��i"D�0R=zƾ5����^T;-&G!�@���a���E!��R� ��؇�>�� t�Z!���w�\�sS�C��(O�'Xs<"A�k*4w�Tu4{KD�ww6�򟕾63Wi��&B��i?�_�
���Ƅ�cW�"��캟�U�a]R)�o�����t�~L>���������Ꜫ�$˲�]��3Mk�m��'-3���M2V-[���~�.0�dG��1\����0�n�.mc�H��IJ6'��a�F�(�鑷�` ��B7���9d�[�o�W���]!en@Uw��?h-ϑ~���������8/��>�����.�`^SX|���hl�j�f!F���[HX���23ף�]�M�5lh�,l
V�6���ir��\X��{>�S]>RՕ#��s�=WF&jEӱ{���l���P��h��h�z�T��K]���I��� Wq�,G:>�n�+2[-1�zTc��{��	a��'��c�a��I>���X_3v/Y}��@mxN�q�(�n�<�)�L�z�f��4���v���2��v/J�� ��w�)�iB��̱��_�F��0_�2���s>')�AbO�L�����If�yS����0ڞ�݅��c��������_wu��*?f��4��m��1J��A/�C�r���f�7m<X�P�b??$������s�QLFӢcel�u>��P.ڋ���;I��~�0澴�0�_�fN7xW���IH��n`�6�����6�q����c�����f�Ӭ���U�A�|��*���K��bjbk*����HQd�u�7/�Y�uqg��%���W|��V� ��jϿ��ҽ
�Z�8iAZOmdٕ��"���d��X/����H�0?ވ-���v�~ N��R���������v�$O3Rڷlؠ(�#hbL[o�W��'yiX}fG޻��XPZU��ߦ
3�o&Yi§S^��1�6���x�I�;��_`ܽj��ц5�0+��z�hpj��j�<�.L�����s����=hCJ+h�x��l"E�{�1Bw�9"��Fգ<�*��f���>��l��fu0��e���_���f1��!����B�����52�a�^�.�,�v5���d�3'��f��şWε6������R�>}��?A Z~�S�f�O���
��&�KWǎ�+>����3řon' w�{��s�*�ġs ��� V�����Yx�-<�u�!(��^ۦ��M��N-�x*Q�^�����F�ŜI@Po2���mfwՇ#��Y[�D��8Ƃ�(�y�c�=�{�

�ӡD�vSa�D�[��i��F�<���u�4~���4F4#m�6�LܺHd!=Z��l*��[���bO�M!�}��n2���FO~�֌�����DBł���WG=��;	HsS�A�}t��"U�'�Q�"T�f� �U���Z�N�x;�Ft:_c�ɤ�:�r�g��Z��V��N!��ٷ>�[lEX��i���nآ�4����Rǜ>4w�x�h�@��AM�yR�P[��~�4�Q����Ӱ���u0���>U~�����u���Ro_Db�:u��חK����u;:Γ)�6L�m�Tx��vp�oq8\���Ճ&S4��I���8�u��p�_b��h�u��Jdל�v��A唭������Θ�F$���A�\�7:��X8�o,,�r�:m:mJH�e�o�[�L�O�d����h�N��jbzǋvYM����	�WX�q>ŶS��-�����l��$���z6G�5q��������zv���	u�^Bّ�Au1`�kㄌm3+E{
I�~{a��*
n6�B��Z������ ���7�A86�S#���/o�u~Z��y��qŻ��3���K}�{�m� C��RI}@��a��}E�@K0��Ŏ�_&�T�5�X��jk'��[{5�1ͼ���� �S��Ć]��s�گj[��+ÍRƘ-�H0��j��i^��ƞ��҆�?�I(��z��B|��)�������~N|z*�$j����cN��('��P��B /��6�?.�a���8���4 bPh4��m�E�^���>���.�;�%�)Z����nB��)8ޓP��o5ʫ�3}�0(.��T�C���'k9M^.��:�)/�!�SXj�݄�?'��D�t���ST��'�����ɳ�<m-@�\�{.�u�{���������<��_��b3̪x�h���=:G[��$���Uv�q�{�m�G��@hs3d���h7@�*���wݖ�t6����t�p��U;��s��K�,.�>��fw��x+����}�zh���5�f��ٸ�vx���U_�$w��h����ώ�S��4˷����w�#�e���
�` �M����������\P�Mmq84�)�k g���`X�i��E� �[c���dt"�F���B�T��t+����t�&#�*���c�%�	s�?��Za.�Q�2�6��xo#���2|`��Ļ2��s�S�Q������1**�:0_�
`
���PV���E�7b�*���%���P�����!��w�a��Z%
��#
��6a׆��0�Q�A
g�y�Q�2�:�g�um�w��(qF�@7�kH8s��:b�V�:!P�;f��+�28wVM�V�ߜ���Ag�i����wu0�J�H�,��¯d7�`:�����^6�'d8[ω��E�P�)�����l�N;�v�쒽�<#���`W�+(}&\���2�������#g����6�8D��"��������H�P��QLU�W�`5&Ӻ�+ǣ����5�	��ij�v*d�G�V][�:�pς�Y5��޿&��GH}�c�>��=��$of���ލ ��M�zZ`�k��T�:�!jp*~�����[*�X �%JRQ�Y���N+.�eWJm�8C���	��ؖ���������e��6�GwN28J��&e�� ��RD
�\��e�2^�a�tl6�b�$m��	���a�0:X�[N[##Rao'�z�U�R�xo��i���#I!f���c8�f�\׏����?X$�>\�^x���	M��叉x�{h,!��=�ͅw�"�Ā� ���}���W��zˌJͽi�x(�/x��l�P�ԝ�뫙��{���?!��́�h�����!�UQ܇5��7�Vf��hT�T/>k�NAU���[�"�P2`_/t����e��⻡�+�$�����$]�fS)����?L(i�n�Q�I���Z�-T��8wwd�����)X��vc e�����.�Z2F�<,�7a`�6��5��%6j��Lj�.�.Y�e�sߔ�ϑj�5θ�)ox|;����z���#��w)A�l��B_�H���S��L�0Q���P_Ij����j�{�Ǩ�Y�*����/���[�i|��0��5Uيy�r'm��{���`-'tw��	��:u����zۈ"�
���H�+r$�S"��犪{*�75�.f[o����+H�6l������*d�Z��u�M|�ᪧ�� �0�����߻D�BJ���ؖ�@'c�GTCr�@����oQ���C�=gH@��`��VPP�Y5�Xn��楿
���W���������j�w3ӛp�Byu`�j�WZ�qS^e��e�1����hXcjގ����:m���r��Kӗ��W�nS�!�8E��ѳ��ݸ���H���nB�YO�/���p+�?�����iI���M�z�m�(dM�YY��'���@S�L��o36}�c�_F�T�H�`#����{�R���|=N�P�C;q+��c&�±3�1�fe~�
['*4I�<��c9���(�_�G�LC	�5N�A.	;�,��G�&
�J�^wx`�l:KJ2��nn�w������cጐ���tJ�����Fy�aи�.��E�3�k������6�.HO�,z([��9uu���o�$�v)�ґ��n�*鮳�Vm�v��j�0(��
.��!7�z�U��9���1��<\4�����(d��C����c�Ç������ae ���X�7�ԝx���0�{�0�</4}��;�/�W��Au�s�˖i�fd6�����9��R$����C�h�9F�������,��Nj�0	��YD���B[O�Դ�[�V����U�C����v,����컇��LR:l�HJׂ�D \y�xG���}o� s>��ۄ��<�����-D���^�g>�dд  �������cFC=�&���l#���?� �'�@��3]Xb�����zυ����h�uxG��BF.\ P�J�?��� �v�ݑ���=�M�	�O��R�2���!�m�u�5̱���yu�+��*66V��j?�ȣ_-W��S�Y�*��Bҭ��cA���W���@��6{p֏A2ur�۸��Y�-�֓ԾK�1	� ��N]3d��~(0�ώ��o�H�=`/FG�ˆ*R`�Y�	<�3��� q{1�F������~HX]�*f����H� �f����u9�4�ɐ/+^�|dئ��3�(nЋ��pk:�?hL(̦L4x� "(��i�=��G����A=[+&�mv,�񩝮e���?���rb.��C��="�X�
��pp׾�G��gY�)��K��y��䫄a��l�G����C���2{��,9Q�Ƴ���0�7����O0h�d���
�����ŠV���
��$ڃ:�@�[�]M�j���Qi�!���q��������;§���Wq��D-���u�����ᾔ�>�ןQ~��&������[Z�P<�PO��c��Z���P�aT���Crf1*��V��L��甯�nJ���X�E�6�����߱�|%Mr�<~�Y�"��x�n�2��|�7�F�ͦb$a"�0�9w�u��e��f��uܩ|ۍ����+���� �M��\x~܎����ѨFj{�f�x��ა`+��b ~2��Tz����R��rW�G~����GQI׎����ᜁ�y��$h��V��r��,8
$����^�}�t?��"w#��-U��_\ �ٞ���-8^�"mh�����p�7-�_)��+n��Z���+���)t@��U[x���qtj�63��&H�K�@�؛�w���99��ۓ������}����`�pi�WG�=ʡj�85���$��v�����p��n�o�۽A�&(k���Oj�دt�9��NY6��=�&p����>���4r'�g7��n�Y����׳e��)B(��P<<�1�&�	г��=�puf���ς9���r��;<�a��I�Ro*A��bBi����P{;ó+���ST|J}��Q{�{�쪴��,	�
���L0"$�!
i�˹�f��?b�'�5���#q-�[^��������������xZ�,igÑA�'H{�_E���Q�1+RP��K�����G��%rHV���%�O>�Co1��h2�j^�W�;��}GF�V�Q���;8O�2;����Du|�'�L���XVO�b?�8��G����}H��B�s�p
HuEJ�º��������7W��+�O?ZM�����V��"=��:uK�H'����%M��L�(4� U	pO�"L�P?�T�����V*xr���o��Q۩Zw���/�?����	���yE�-�E��~�n�U�@ K��1��^��0=���,�ښ�1��s��B�3`�S@���1��=[�˃ܬ~�qȱ�r���V��6FA�� (�I��f'J���ؽ .��9��J���ٔ��3�a�5��8Ȳ��!"���})U�����Ģ��C<��ǖԄ� ��<˃�.�����>�ifTC׻hXD���˯2%��j�#���:�337���ꅄ'O���bI��g�����
�]黊�cqyoӄ{B���:'ځ�8s���)��)[��a�,.�j ��v�a�7���T�
 ���,\���,��dOZg) u[�N�y�hŢic"Z��e���!l�=k�&tW���SZ��:쩅��d�K}g�ZZ@��F�k��
�R�֗�����q�Z��ɽ-=�!>���v�x5�X[^�_O��S_�g�X�_��b��zƦ��p*w(�7��	4�S��rd$	����t�}JQ�����r��!�	y���J�o�mHT�3ZFd�E$j���5D���b:�:[a��',M��� ��}����������p��
����� V��A�~V���7��Bp�S�ԇ�B.8��Ҵ���ҋ�,s_���ƀ
��F���M���������1~-�`�S�������D����3�
����zM�;�(��N���U�$u��L�)w��d�g6���Fd�γO��� �$E�Q|LPAO2O�|��j隌W\{q:(f�Y)"�]�&;=����vL��������)A�vo�{��(�|��q���F@��Ȕ�)>B�fY�1e>9��>����SH�gT�����Z]��th����2��{�Au��r�^��A��}�)T���_ohֈ`����/�Z,�+j})��E�����hB������LD��n�_����W��5N��{��;���C�D?=�:q(��
D|�ϐ���Z�]�n3�&lbL�o��J���ΛJ������S)<��ӅҮl�w��x�й;�	"��`�Ж�tۖ���7�$�%��8S�����*�`�`���]��=_��hF�!58����f����	s�&����9�Al���r�C��:Ƹ��tD��	(ZAUn�A��w{��� 5���W;(�*��	`�T,��]�'��/xxB9����>�~|_P���6>k��[:�b��6�\ԟ\-ܰ�k|;���eY�
W��m�U�!Z�s������y�"�DQ	'6��qC�L�r�~^DkI`s̳|��{���߉>/넹�w���v�-(�7靉��H_���7?�ە�1����Դ�DԆe����5�
�O�.ѩEY��J4��I�Q�W� ��HE��s�<�u���$s`A1�OEb><���zY�G}�����E��$m����[���S����V��S�f6�m�O��0�G�s�M[�iŪ��j�ք�w���pM	i�5N �`�5O�j-{�C�� ������������"��@�� ��2)$)8�e�@�+R��kM�6&�̬@���j��~��Ӫ=����(V D��v��� �+B1�j��o��BC��J�(�΄���{�� �SL�Ɉ�8(mZ��P8{���C�N�n{�����s�^��K$	u�ç�,��3��;C�a�C�p֡Q6��r�����+7��|�V�m.9�3��{��Tܸ�$r�)_O{� �S��|*��ɕq�<{C�H�%:B�aї�~ɲ��_2]?H+�f�I��J�r1%�A/Vӯ_��R�=&x�2~�t"�( )���|^��<�חK̇�.T0qy���\��kr�OI����"�b0�g��W�fq�?ҌPKr�@�b17,��(t�z��: NGQ�O�N��������b�laS��PH�31G�jy;:�[��#�#`����oՏc��Y�����)����A,ĩ�I!>�Ѫ�W��R���I�/���Ð�:6" %:;"�ap������w�}��"*��@DnR��_o�rqVQ�_�����W��P\���$@I~�N��϶�R��$���"	��J#�!O�!7.|�̩�Mb,Z��$������1EˤK:w��cVҊ�16�zt����k��x���]���7#�	�L)�i�_�oh���,�	��e�9����<��A��V #��7��e�P��ۻh`��[�����3^^�����\���'oz�j��A��%T�`��KIRVIM�ɒx~�ծ�����+�8z��qr��8-5�m��P���lY��O���w^���,����:��;���ʀ;u%Ʊ�"Tr���@�[�!�Aɐ���7t�M���;s/]���u��;��F�	m��}$B��  ����"'�n`��Zy���3��9�"���+)�zO��<?z+&�@��{d��n�ԩ�0(wb���Ν1�oGA��\���d|�B�n�BG���D���c��C'��l.��h&��^��N�oR7~�d��#{	>���{n(�;M�x�q:���J<�l4%1턕[)��vʫ�Gf[�=��;�H�K�O�G��1}�D)�ɴ5��5U/:�G>�I�)�`�BF��Ƞ���K��{,���yt,�	V1�+��qK�
d���i`^�v�;?��W6�Z)���9�.<�tЙ`����Z�r�!�l�\a��^k��Jk���r�Ί�T�� }��T�2p�cs�s�>���qY�cj��%�����z�}� �i1�����c����k%��-2 ll{�"�ŕ6�����^|[��0���{B]�Q+�w_T`�|�V�Bpm�n87�4<��jkP#�3�=�z(�H��s�AWbr1?��G�=��HC����=��>�1��$l�}���B�N��B�h�;�(�<��3t�� ���E<�I�Q����Ųl/�]�F�5�+��U7��Ȑ�5�&Ġ-�w�aK|_�)vp���9O*"&��p� O��n�7�}�(�!eY���JCjE;
��R���k�͑��;�"�d(d��L��`(Oj�(��C�h������n�h4��n��~�u~�DL6�n���1(r�٧�߂+`l����RJ�y�e�zx�J}�;0�w>7�%M:��L0a�l=F!3C�LѰGz��~
�+%�gH��.2�������*Ҹ���Jh�����Q��eI9?n��gbQ�m�Ww3�K2j�8�����Ć�S#��?���CB���
mX��$t�/�+�?KX��j�t���Z����h>��ܪ��BN���}B�r��W�[^ �u+�e�Q�A�mg:a���R3s���$���k��ٿ���;�զ��a��1W��-�9�J�S}�V�Jz[g:���pe.����}���M˳R��������s�+ҠБx��1]m�q+�'1茶̊'�9�.�8g��iW;%1�jD�،}�����.چ\K]�>���@*���K��J�a�`���P&e�B��"�T�6|�k+��,��)�����u���s���p�y+6})���@0"�����8�h�5W� x�>�q����,�*J%�H��<�xQi~
`�ܲ�+��`�O�����V	�0[�Lmg����h&cB`h]��!�ѯʆu��X��^}o�o�$rq���lWT�G�#��%��`�/G(e��S1s�/#K�?t�贁ݶ����~6�&���l*���E�553�V>з��qy(��O�C�b���fł��]��zX(h�nJ��	��Z�����0a8g����[�m�zΐ�Z�A�`���4�&��v�Y�E��Y����e����x�G�����wLM�n/��hd�w�j��ʴ�Ǝf�RG�(2�����b{�0w��.��*�4�YW]9�^�ͤ.��5�-��jfN"��OZO�	����[����j���H&o��d+�ܑ�W0��h8h6��N{�S�=�Y��ra5KC�z?d{�'���
,�-��^�����<#�~W�P���B��{Hh@w����N���
!�/cA��<�􋭺b�̫���@N�������Q�UV�_U���#l���h�4rNaO�v��x���v�ԏ�g�&��e9�w=$l_���1�H�3�����B^�l�ރ��5N��F�a�*$D�y �.�cd/��ߊj�q���� v�xJl^���v��`m�>)�ЮZA����Ց$�+�T�#�S
%�J
�!_d!�(	b���=P��>,���֞���Q>p"�-?�,x�t8�%7{9���QZ�W��{�)�L�E������A�D�<���7��m�(�'�
�s� ��ʹ&�@���jy[����"�R�_�/]�(4���n���r�@�'�mB������ki�C�:��_���e����ȓ�OĢJг�$z1$�'���|�@O�'2����+jR����*�� ���f��zO4�_#�M�a�SQ�0L�����?f1�=�J��A�0i$-��p����Ty�|�d�y�ޚ�;f��rl)�?��	g�H��u�y��d�
g�� mpn�Pgf
�[��T�7�
^W��E�jʽ_�&���V��UG
C����1UUB\��3G]��<\ѹ���Mg	p כ�V�W@�b�>���5-]=U�*q�ԥ1ߵ6'q���Ptj�׌��EԲҦZ�E�WT�n�잁��� 2�@;������u��v����?�~��6�G�Kb��|R���AՋ��v��y�ES�D��Iz2�k]�I�tBL�!f�i��g��QHs��: ��fV&M�Y�h%�z?�mѨ����E�	��A�	i�=.�-L��>����,忺0�pQΥ��<�ֽ�T4�:�����p�$�ʮs�g��ã���d�y�n����i����r	<�f8+U~�R��t���F��ː������A�'��@RRg�D��!	�dP�y7���(윆���=���"���U\���ws�j]6}��ᩊ�?� �����Z7$-�'`?n\��*Q�C� ��[446�s�>y&�c��m������C�u!��*���2���0@�W1y��+�7p0��Fy��o�R���	b�%aψ*��O�F�K�� ��6�s�<ja2ψ@��ۯ�j�S�&ҿʴ,b�>(��Z�)�\��e)��Ez�ʅ+۔���ȥ��~�g����U L�k��
�	iG�w���>�ڣ�A(d�>Շ�
r��u��(��J����+���ڔ0����4ܣj7�PpK�X�����,�����(kr�C[p.�lJ�A������YC	�J�Gᕰ��Rz��]B��4�pÁ�V#f����x42�Դp��"��a��;�x�Fcz���0|��w=��y_���Z��1�L��ad��i��O-t�� �ů��Es9)z�o�/i��*�5t2�^�|��|�*�W� �g԰R���Ҿ�q���Ú�C���e]��}֥q��8L;E����ьۡ0_��0�x�m5P��+�����s�)�J#
=Qm/U#�k6�Z�~<��q�Cί��5�b��\a�����ʬ��5��ժ����Ȃ��Y�ǵ��E)t^�٠4�S%c6q�6NA�vn �µ�V����R�Z���AH���A�+���tto̩��IރsM9�b�ov�~�q����Rk�s��Oz�c-�+�@�R��=��0�)�bN)q�J
���t.5B�X����D�L���V��m����:���|�?t�?7���AÏ��a�U��
�����X_Qj������d;p���<#����Y@�^��qZ�S�LSC��16�t��{hh�#M����s�!��˖�,^����}c�BdY�o3�t��.�5�+Hy����-���p^4$�FO�&=�G��H��֒Fc�q:���:H�w�]�w9�-+�2�^G18IV�?�����u����jYw?����l��0p���EK��R@k�*�X�]`~<zː�َ<w�.�������G&} ��dN��VY��x: ����B��������b���g�����Y"AA�ɬh�G��c+��0��+ˊ��>�2v�>����B�m������;{�O� �M�y��\�۾+�҇'�lȺ ��ƨ���BD&�(<31�?����ݳ,��\,
�܁��E���qu����[r�2��O�X���n��2�x_'azj�ƿQI��tH��� �H&a���(��?t���8\�<�/fաێ^���`)��;�J��P7��u<��耰���K�

�!t\3o2wMȻ�l{]���i
����.��Z$�e�$�v�i���7vm�m��)��X���%�F��J]Edd�p�:s 	&�T��Q*��U�� �K�I��G'#�
�A3��b����&���zO9|�Ht�B�,_�n��F��Z:\�r���F��T������*Ԓ�m}ʘ��F�O��.%)�/q͵͊��xoA��H�A���(���3�ȁ�«�FS9�N��!�̬ܪ<":D]f�n�M�U��6N��8�r�Ƈ��R�19�V�����!f�Í���₩+��&e�6�AD�Sl�
:n����6��q���[��3��դ��@Z����S�7J������@�c��[�[/|X���ͮ�5tٰL�8��A *'	
�=m`��W�W�,V3=�+4��j\*<k	����O52�1�"H��G@�~�i�|(���JA3��>@U�2'J0�!��N�}Iq˳�?D�?2���|���Oi�ƚ����3\J;bӎ�{߉<� ��Ja�#�`�{ 2]Q&	��r��-h�+���{te��'@��+(�H��T��y����7�&M��~׎�I5o�f��_�G�PI�O�#�o� A[5Uh����X
4o�#�����NRE�A@eTV+؊{󟱋�Q�����:����Z���ʶ�Z�ן
�|ۍFG�C��aé��j�T�q�Y��� !���qSUn���A�E��cwt�G��M�QE�%�ƧW�|��&���^5O����r"���Ju�cw}�۽���s�q�����{���D�ՄC�-�]���m��j"�&d��^�q{d�<Z�"ͣ9Bб�M��|�3�G(�W��P�"�Rm
��9	l��oYP2�F3�饯���Z[��S�6�A:���]�c�X& �)�e
����s���\�=��	�K��z.�,�O�{P�(��38n�b~�Q��֝0�r<�.-��Լ��
�:�T)n;�$p��x�]�XAtW��{�M$J�2t�/�Zj�q��l�Y�Ʃ�ɠ����U��W��S�q�#C�dfgCz�;/��y@$�z�d�Q�w�'p}D�X�XR�\J�Ԯ*,콳C�M��D	dGp��E#�
ݶ��&#��^)ȡ����@q&b-�!���j��G�re/CI,o�������D_P���]�G���W;?6����S���Sag���
X�sZ<|R�ኚ�b���}�^�U� e�l��f��+B�r�jY�8�Ǌ���E�~��_�NϿnr�}g>�������U�ۍ�
�R��S�CF��ST7��z( ��y~�4�b��K�U�'p��]�9�'D	��;	i�r��"�\�~�y�M��v�Bn����������_ �����:0�)]/R"�AODܳ@��z�hH�I�EL�4�w]ۮ�g��|�rQ׌�͙:�K�n0<6���XvLLAJ aXNI��=TG��I���@īV`Ja���}�_��m�<�R\�q;xLoR8����2_�||��ܤ��D*R�a���������G*:�� Ö;��7�:��� Ġ-F�ӹ�z&Ţ�p��=�h����G���̢[��i\<�Y�t{��Y �"���w��05�0&/���@��laJ��x̍�l�s9?�����W8K�eI ~0f4f /tL:�L�Kun�D�ib��MVOc>@��r��;��d��9=�x��\��MQ��{unS���l�c<��^�=� N��v�
548꛳K�ɨ��_{����$��|a�7WB����"�0�4!���	;j[:w�H-G(-�z��J�:'D=.$.H܄f+Q414�g�)�
������ލ�cq`z@P�mM�
�`�L����)�\���$�;�2�U|"�Ў�uH�;���`��Վ�Oٰ_m��_ۙD<�
e�a��8f8o��U<��TC�q:�"��^v�"�q�0���Rxkԛ8��pwYN����O�i,��}̯�(�\�ai���r����#d� ?νH�*,O#�Vȱ�8�3�O#��.A^���L�!��p5Ňנ���̭��M[�~�gև�i��|4ZX��.SJfU�gT�U@�)�%Ro�9�$��R�.�>��V����rP��}�V���ҁ�Z��>އ5�Y�Oi�E�;E�"�b^[�7��N9���P袇��(�#�r��;�~��1��o���l8%����U�/acJs��Pd���6L�2�Ғ�)kH�`�Gĺ�A���tB<�7��߲M�Θ[�HU��4Y+XE������ ��S�� ��X��yHZQ�rߕn��]Oj��Ǘ�w��2�<,W�I�K�ۄuC�9@��}&�o~sHL=�2�BE�H'c���=;1�x�.�I�`o4���p�R�ܰ�����v7�yr����%�.�B��R�) 9�����3��U��ݽ��6osGt�l���)�QJ�T(���=쥵C� �̄�\ҹF,;�w�6k�?�G\�7<�~��1F2F�&;W��z�k(�Rߟ�c=��[��į��Ɠq��ݠ��W1�9�׈��*\������6xE&f�|���<�x��>Y,qu�y��=�[Y:�x�ھ�Kޅ�h�[��p��V���{�<��,��̺!�y//穁w�_����wM�-�ޑ��8Px�#C��$u��}��%�@Bũa���)9���=W0V��O}��`߾Xh4��9|l8{E|L��*��۰�3A����=N�&%<�=���u���E���e�(%��?�=��15�j+ �l3rT�v�*�-b{���`/�w�e����I�x2I�A�b���}� z8��� ���b�Se򫄷琖U�'��O��q�խ�]Z����8�a{c�Iפߨ-->�X�5��2S���)H%��&�>�L�K���Az� g���!�dŔ��m�k�_��)nb;}�� ���]B�;d������Q=!��)�$<�/N��)�7���j���	 ���/�Y�#��o3,��;�NN�i�
o�u��	�����D3  Am� ��m�z�O֡�"�����h-�F��i�o��(	�_�EM���(�J�V苼#צ����޿:��UZP���1@��%kN!�g�r��a�ղ=��~���w@(��7=���R�Ƿ-H��x3�%�y(�L�r�.~���,��g��0�5s�&2�՛��|s5���ՏU�qE���\/�`c����<���]��&�(�a�iw/�w]+�Ș��9[{4C�ؖ�!k�����my\h4�w��vv��rDlw��na�����9c���ݥ&y�#���|��R��a_ �
9�ޒ�\��_� 2t63��Q����PPF�i&��مv	\_�f���#�����av��$�����m��1z��
9�{L@}�kN,�X�1H����R^��9l�_ .�N���� �|�Q�As�	�Q����߷� q(N$΋\�'y����ݬ!�b�=9��ۨ�k�A��'�L�XYoF򛩾�c�o9���y�7C�W��e@�w�M�{��5\�&BdRf�:��⃕#�i۷��Y�*=�k�1[��A�|]���\rkux�����H&��z=��'� ��.�G}j̗�&~�oo�E�M��\�� �����l�����.�^��{I!x��,B�N�:0�쫡��R�Տ&���i��~�\])��k_�Ɔ ��&�.�ߓB��K�6F�}���
�t>����5�Bv��6z���m`a3��\+�O�U1�M�����8N�e�?�HW�т��� ��m-H�*R~��C��u�y*�}��猈2�7�)�ZQl�Lʗn��M�'�x�3�I����|�}�	_�l�A�h��є�2lJ���B�E��+d��I�[�k��H�SJP:�H��e�>��y*D�%�I�`��6X bn����,�����E����M�� d��%���h�I>j���}β��i1;
���<&j��?,)��LM�$`t���ޠ^[p���nlx�}�#꒴{&��pݎȣfyd�s:� �m�,�0!��aH{�d����_�VQkK~�ʍ*
��Rr�[H�X�d�	�F�ta����#�1��!���W�w^C�*A%@%��S.Ō�5˳:P�����3V���=р���Σ�Ȱ%�C���#�J�([�X>�{����=�K�0C]��	�KW�~��[��X�_��$�m�X�y"�p��i\��k����{nS�8)� O΀k�C��i�o��[(Υ�-�D�rk[����5r�Y���!�Z�O��l���kJ9?q��lh�ŞmͰp���]g�]�)�pk�j�e��]�<�wt���g����3�C1�Z'2a�2�-^�E/�Ӳ>5����҈�f��Xs��e��n���K[�yv=�HS6 �d�]%*�{�,O�C��)���P劖�J��@|aj�7G���!xF�~Sx���9D�k�!�o~�I�*��A/�-�]0���[%�8@������ߑyǓ�`\	-N��@���:x\��(�ܻuce���H褖�2�[g�z�{n�SZ��+���k�NV��D��i��:J�f3���"���w��)p�
��?}��N��v�<w>���T���/��V�ک䠿+��s��*��ϲ�kI�6���S�H��
S����S~u"o�:og�%#��Z�1�]r�WZ��_R,�h�ɤ���o$2�K/켰�4��w�գ�ؒ%��з�����I���k)��j�@��_v�gD��~�D�� 
,���J�x�jp����������d$��B>(�^fiW�;*Tn�b!�Y�|� ��m; �E4��5�l��%��R���8f�JM����'Å����ʰ����T3�Mʹs�*���]+Q�U%̘zp0��j�4�/ݸ��p��r�v����t�:DW*20���1v�5V�$����G0���|���e-ݞt�h���DN=������'���	)Ր��tK�Y����qאr�6�,	+ M������3��*�4�ʹ����Ӄh`T\տ���K�[f��s�׏�ӔM �er�-�޾�;�/���)��.ӗ����t�L�ۤ�P���՘���Źv��H{6���Od�.X���gm!۲�h���Ю�_�*6N0o�֞�Q���Y��X#��̰�9��UP=����]X�0B�e� q!�|��)#go��Ѭ~�-G��ܩ�q���e���SjWr��M�dJ����N����N�����"������//r�t���KF��ݛo�8�Zg��$Mh�,��sn�pdz��j2{�Cl[��d#�Ŕ?'{Tp��`$���$</�`�)�y�2���;p���L:�hy1%�����E$�59j�̴��0�u�gsG �z�7�"��(��澀���b�u�@��n��.�`��gΪ�m>/_���¨�ݶ�* �D�����?��C��KG�G毝Ǟa/���Χ75Y\33�0�<t�ݰ�B�m�,��a<e�ɮ;����p����L�B?C8��?���BJ��HUx�SG	j��ZJ�6�ʊY�װ@�G�M4�Td�y�E�L�S��I���\u`h�������J��.��=��0�! �t��f_PSv��0�՞�24��Y�� ��P�Y-]H�=iX��._���6r�8N�m�\l���'�50�[PY��ѡw�w|���oR�n�6�n�2��O8���.��!>��:�����؍L�Jl�W��S�.��Z���쵼�[�פ���I"X<�����i����`�<9%���ɮ+ϫ�]�.�{�u{�Y��t.Q�s�>��j����"6�Jʐ =)c	Yd�S<���1�R����*��X3q�*f���+�n�Պ�Sy���L�Ǻ2ʫ�ws�5�H������[s1Q���>\� ]Q	���&���Z�gb=󺭡/6������E�o&`�Y�]3c�2�5^@T�V+*~+H��MV���o2��/j��o�i^F�Y=V$	���p�.<e�=n3)� �ħc��}��N%����?#�F�R���|n���w���5,��-3�!�q�Z�=pg��i�����Z|]c�n�Z&�"q�8��ݑq��]g�ڪ�ſRkĆ�R��yU�z�s��������_������e>���H�6��]~��{���:����'�B������ո��ܙ���F8'Y#�� �PJj����ק�Z_��S\kc.Y��k��F��rƞ��h+шH��`k�������TU}��iY�	'�����A:�uە��.�V�rJLhpB�eo/�CMY+���$I78J�I����~Ps�R��F�f��S��o� �(�2<.'QC
��I3@�����uv[��j�;��R`���$r_�R�3*_y��;��g�~"A}�_��/�1�	�SB�"�V�0(�\�p"����V'�����Ey'm��"{��������.�[N>�u7��C�}"��˞�Nn��h3�Gu��z)鉯;G��d�x
�֝�eإ�F��:@M���8�$��谡���K���g�|"b�d�����
�tؗ�����#���)�^�3�-TM=�瀞NCx����C�=�CE��ӱkZM�E���:\��.˝�����#�]|�>�6u��7��9������ֳ0�,�^*R���Қ�M�ʿA�/^n��u��0(P-=8� ���Xp�z2d�*ީ�oS��/��F�7E<9Б
Sܰ��A��������m<�Q��֓H�W��}a��9�3+���~I�0�5Wp(9�K��"���Z���{r��l:S�^��*���>;��T��c�� �e)<�᜕�k8���C�Cq;!��uk�k˺���&~�\�'ԈÔ~o��%���2�*K2E��G&P
@�`EQF�����402��i�����ݧ�뺡��l�t=I�@y���qj[��-��CU,�R��L#(8��G]��k�0Pa��#��\*m[����{�!��j_�3��Q����h=}(�an�����4h�����(����^C����f�x�R)cXፅ��z4�o��{h� ���&L8:weM�s�C9ª��	����5���itگX�1�A�x7�׵+��M`'bR�	W��n`rD�6�Wړ.���s�Bd�U7zƭ8n+㎖A{�Hhܑ?�==�"�:en[�~)��d����#5�j�$vݥџ>J �K\��#�g�����p>�J����p����c늹Q)�j�ErO����ְ쳯�IB�\)FL���p�% xp�8�zc86�w���Q�0ږ`SV[�3�olR��9P��x�A�,�̧�P�U��f�lz:���I���T��پ���\mMz�Au)��6Y���OQo$�vW���'jQ�+�p�I�1W�G���W���Vi��(��ӭ�Y��'r���2&���Ac�����Ϯ��P^��h��U\��iE$��_@����.���DH�mK���N�T�n޾�5��^"���d�x���ǣ�b #�1�+t����Y��C�T��r#��w�B0�zC+�g*ք�m��X�����X*���mU'����H$׎H���xc���:���4y��z���x��F����;ĚHPx��}k�[�����@[f�}�a[Z<�s��agհ`%�O
���}(� m.I�n.ToI�׶.)�R���?;��X0j�B��H�O���iB��ă�hn�<�?�r���Q ���Sd�t1*W�9)���&��b�t3%2�t���a%�ð�I�O+���	i�Tp��3?V�Xѽ�^� E�Z��(�T��9�S�-�0�_p4�%�@����-�,.Q��yz������d�R��5�vRW�*g`r>���E��Kh��*� `�)d�_sW9�Ũ��?(�Hg��3Ln�D�b)7(4x�h��/م�M��*����q���(�>W�^c�%����G�%K���`�9�i�@�wX[�c��d�X~b�ğd@��6ef���� �2�L�"�������7���>�.�w��]M�b��@��[g��~=MC�*3?'h?aQ�].��0���;
�ׄ-./½{�D�n����p+�����J�jn�]��n܀��.��0�w��2�lxX�΃�~�M`]��1�����ݡ4|t͘�F\����7�Zù�< ���P/@�(��O#�ܚ���?HGk*�%%E���wHZ��(�΄��M��4���Tp��(������D�w�J8_��B�n8z*�N���ϼ �F'
���Xw�h���	ed ���2BD�>,EB>$Rt窋q��X�,�݃q��>�\�)��pU���­������ܝ̓�e]�k�L��&�����b�2:VC�A�E9�ڻ\�Q�r!��8I��:	�'PH�a�֐����u��=W�5�t�_D���F�i$�P<:�������?��-@(�)*�oM)ICM���e=��oO�"�q@�qo�;�f��h���6�%��h8)0�ȓ��0����O;Ez� ��^���^�����4M� �8�I(?�4 �,��s���:��Nf�m�_�7� ]��m��\�o�d��%��� *��N��������aI�����1�,U@�܅5M2�*O���1Wj����ceҜ[�v�g>8�n�[�n��ڹ7Y>sBm'��0�R.�:`�b4��ȕ� 7_C�V��y4���G	�#��J�ƞ�}��:����=.�?fS���&&�[�	E5����������~��fӶ�j���
T��ՎB���ze�=��3�aዧ�a��"]�4��.̩���&??X}��8TA�>g�_K�Dj٘G��5X�6b����ňLL~�P��o���D
�0�Z=��E�ԙ8�T�p��mɸyQN�^��aV�\e�}P�cK�V�}�x�U�(zzӫ.l�\����P�����"x���'�/�C4񒘆�z��/�(�}�$��vn��u�G*�!��4Y]��)\
��&d��$��s8�1���S�+<��X��|7��Q���Aʗ��=�D"��{�����L h߻��p|ܦ�^lKx�_����������aF��@R�d{w��	&��#	8��O�J��=0��Q�*E#��jB��+���n��$�N����Iߺ��B�l��U�G,�k�4i��f5����rT�}:0�q
tU�����M��Y�98My���y �ȍ���E#ty�zd:D��_-;E?>��l�i�Hb"�_ ���_��*�?�<y�{�U]�չ��L�~~=���������0���BF�E;�v[��84,6(�3^��d���?�W���0Te�U�ɏmnx�������%�Jdx�����>����-�|����:A����j���z՝?��M���U�.�Q@���^�C%���/�Vd�9. G�S���Q�!X���#�x6�#��h���J�AM�R������JPN�r�E;�P�>8�T�Q����j�����O���|�Ё]���f�ɫ���@A�;��ބ�wW3	,�(2�a�2�\���F?���H��w�>�s�M.�}��񰔹~��ʪs�v��{M�d�
j��{�(��1y�֟>r�#���;��6��^��!�@b���f���*R�F�,��B��.�Ii����"W�%�Nuû��(ikt{��.���M׆f�u1��L=C�2;���Yo7÷6Ɍf�9(�Х{� M)1h��J��2�#<�9���T��֞����kdl�D�n�ǃU����V�Sp�9j��
�E%�����֥�~�Ci���-����oP{�T���Ɨ.�j��Q>R��!��eͬ%IPX�����j�{4O�sG�_��%���9M�����%�?�[�
���� ��p��������C�\��M_#���;� �n�u��X:x,�Z�f�k�{�Of
 ��X�*����)y`�5(����Ub���V�80�FB}�:��<5�#`��a� P[��_��Eb������W�����N#yr�Ru=���q�DxEۈ��B�!W��
���AS^A�A��F7i�N9n	��Y� V��
M�}��mI��P���v�����z ���I�|�)ꏢ�����2(��J5���H���v������0v!�A6��#�3r��K����;"1sF/����`K|sh��afܱ�&��8��c��"��H�]8R˔s���� �l@*���7,��� �XKja�6��k���YN"�	��u��.]��,���m�v����}݈rbL��>�FNz��w&�hI�Ϣ�$���s�#Yή)����^^��t���w��k�V����n�L}>d�0ⰴ�����خ r6|����I�F��U	�Il~Ʒ�g��ն�����
:\uNF0�c�k����g.R��
5�1<�E�޼��wcQJA��r�ӪE�٣i�*���
l�4���K���=;��#��L?*G��=?��V{�Ab�����J�	?ጁ݌��o��V^/�.�B.a�ݻT|���4����c��n�������ȅ1�͸�(��6N-n����<���/D��;�;I����۴���W�e:�,���B&$5�K̰�{o%�ZB%��V%-�Md4�)$��kj�,X�Jtd�M���ْ=uň>������&`�<v��1��kw��L���U��W�i矸�GO�1|�-���D���]b/�[������V�P�m�O�94{t��W��2�d��,ڈ���"���B�]���r�Lӌf�a��O�*="��X5�\����︴͹������AM�9�#�(� 'S��U	��<v˂7��r{u�����ER|�u���PU����{bl�TO�s�$���&�!鰎���M�,���(���8�v8鴠��b���A�+A*�����q>V�b������7�'Y��޸Y��[�9&��]�
��&¼��֞�f��a��g�i�y;4-��p0�1a؊o����lBߏ�R�����>N�b�N��u���K�c�,�ܲ�ӹ�7YT�y	��X�ÓLI�m��CTU�c�#h��e�5�S�&",][��7X�Qݖ�j�$#:z�$G�����z�qm�!0ZY���HO������P�u'�I��u��}�#�e�����}�I�2��W�fVz�![��8�Ʀ��B��)@��'����b�5}��ѕD�"��T#-�����x���=�̈́�59��#ӓ������R�udWzl5V=�3a�)3\���$}r�Y����+U�>YR��6�6��3���Q���4,���P�5���T����?�(�
�?���}��%����a�'vo���䭒ƀ�����d�)��l�ω׉KU�zc�[���=�x�_�ii8��"b���.Ʀ9��òq�� xK[Ŏe�5!�vz�U�b�vr	6�Z���i��3���^�7��V�jb	@����A��	�6 ]ԓ,���Dӥ�r#��su�l�D�� �.<_�\
k�\��1���"̕�&�$�Z��#�}�����cV��O�t���)!��-~���^7kG [V�~3��Ύ���k(Z�چ+�O�lvB�e QN�x4.���^��G���^
��^
9�`�(��
�C��}ߑ|i�p�5�˴�km˟Q�D����l̡G�Cb�ux�V�?)Nҍq�����&!���W:0#,�C�6���)��34�l�V5'Í3��'!@�~b�:.��WR8��������Jߤ.-(.���1�=�{��J�4(B­I��������!|�e��[3�e�֍n�	���9dW5j��L"3�
s2�U�J'8ᪿ
���Layߧ�N
����a��6S�ܜ��z�,�N��y�y���"XD P�b��S���0v�"5�>9p�i5U�8eL�[�`$DC`Ï">W�Jf���&
�cT��2_|�01�T�.��u�.eL����g�uI��p�T[�At�(?�P�N��wu
�꤉`�b|~�����Տ	{��\��R�g�X�Gn`ޏ�G���(���YG����V�Ju'�hH����[��)47Ǜ��z�1�x�c ��T'D=_�L Dn�������y��a��+s��e���Ph��[?7�K�-%h��[�,� %��{c�4�5>yƬ��<IyY*�/�'[}#��e�,P��JO���6DJ� �ݶ9����`/iCf&��J�-�ڽ   h6O2�|S�U���OpV�M��ǎ����N�� �Xˡ-j*��QK@���P�>���Q�(hw�׏��,� *�f��������;֯w%�A$�i���S�&�&�p����G��T�x���U<� hnר<��Ѿ���)�ƙ{`ۨZENeFY}Rpϝ`�N��ao�nDߌ���1y��	x��7;n,����k����v���Ea!,Y���n�CO5���G#!�*��JB|�Լ �Mh%]�C���~��ïo6��Co�����Ej6�=yK֖��rFa���{2���h�㵿@��_8n�گ�o�t�q�|�\�8�]	zdU�
h� 'a,t�:NL�"�U��^�h���Rx'��Oڭ��w
�B:ʍ��Q�Hߕ5�]t�IRc�w��6�. �3RD�5L������֑KA��8u��*}�NH�$����U�ɘ>��e�_��2�r1P9�86_GY��t�TT�!�ǁ�3��0��_�a�O~�8ة���{v�ʪ������FLv��^�?]�Z��2���O�pU���l���q��H�,&3�0��I��w$��
f���E���]��[��������Hr�F����)��%%�4���՛�Jfŧ_>��c��qR躷�D�ԯU�U�Wp��pC'��x����X�gQ�������'�9��8,���/�D��!�rk�!�+�7�c��J�~��""E��A�;5�)��u�X����xʖၣS/����B����� {���><@��b�Ũ^0�p[���S5PG���mE���������w�0R��xaM��2�nv��'��1���j��\�w߾$0�6�ֳ$l$t���E��3�bG�{z�g	��=�̥;�4�rv5Jb#1>}iVڒ��r�sM���o�������.�p��w�qR0�*�e,U��"t���#_�z�T�oG�	�m^@�J˰t��m<x{�����\���	z+��k��!��tQ �J�d[�1�f5%�<{!���~Y�ӣ�]1� ����֥S�e i��74d[R��~+��8z7/@86~�**��2y�s�da�x�EU��f
dl�B	c�L[�F�t�n�s������å��2Em�fj[�F#$�V��z^�a�ފ>b��#�@J_�:r�POb�����%G\��}	!9=�B����7��mv���;aIq��8��Y����	Q�Zi?�T8���p��Y�M��O�%��R�≜�ˬ��{I�İ)�B s��r�o >��y%-���zs��m%�p%n��ou%^lk�r�|9
o�4��Sk[�M�p�E@�DhIg������k��݆�^��Z���b���±�҄]׫�����f��=�O�r��ԬMz���"s��d2��W{6�g����5�GTd���T��:����|�z�˾^aڹ�=�%�C5�������'��n�x�~�g�X��2�8Q]�3�Y�3c����ݶ���&�x��ro����`_�q����0��/�ȧ ��8�_��w�%^](�~������1g��!��;��inߘ�ޱ����T�ǂ�c[B�A*dl�0`%Dg�k�$����?�S�ǃ��Y�����H!�D�w/OLz!$gv�����<3���'��گ5@�A�sn�s�Y��kͳ�e�j�-�e�j�ۗ�'^�M�m'�]�HUb��˧�pʕ��ONr}`�?�������q�����d�a�si�y��#������Ԟ$�&�,���� ��M���>>�wBc��N����D��b��x_�����>�jΎ��bz��O%\�靬�-X��b���tl��]�)GLZmN �Ԑ��㏝��E��"Z1���Q���
����X��2n(�g�Y��Y�_7[�u���wd�bW�@!��(�DفƄ�S��BU��H�%˸@�(�a�0��CP�9�i��������b٩�c��tv���n{Z`�q/B����'�IA�,X�&��qMz���ɜ�Á�vJ��<i��8��a[�Q���I����	g��쪩���{0ԇ��=�|��cB�lO�C����F�`��Uz��@x��/��|yLq�n�gb��� J!X�E�CE�`x�y
�Z�~¦��g�ߖ��f[�-Z�����`l̙��er-PSi=�h}Nf�J�����t�n�b
%Cߤ����E݅�MƷ�#����0�r����
�#��e�.���C[m(�7e��Sbm��l.����B�k5��q��߳�����,q��R�U�m]]<���V��4h�~���v�O���^�c9^A�S�����E��o�����3Ң��?��%W�z%�787C����@�T����R�vd�Җ%��r^�ۙ����D7���| u�-�ջ�J�Wg�{��0CG9�3H|b-��0��<��d9�`\5��Z�}Ӟ�\�"/��#*ZBp���{�V��{�Z��[`w���r?���'
L
��T�H�Va|�ri������%s��*5�������0ؠ���!q# ��$�i��$���� ��u���Y�����CC�'#�Sb�HFI�ک�5�>l0�a]I�hԕ�w��~5� (�2ܥgM��tG��\� ���E.W�-2��L�p<�'�i���*\�	�qcP�f1�O��A�D�,��	 t��Z�&?��&�7о~�9�lc�!���?Z���$��!ܭ6eq�k�O6&�h]����3 ʶo8T�҆���v��\Ź�B8�/� oо��O �N�V�[.�W�ϻ�~V�訨$���W�i=pe�_���ߵ m�}"�ja�u:�ٕ�H�$ n��~���%��J[�X�Ӛ_�Q�#wtPqT�@}��;��Y�\�Ý��.�� �XўY�҉�Fv�C���
o������ w���	��y:�&�w��h�]��
�����)�N, ɵ����++���B�W�Y��9��G�v�p�Kq�q�R�Z���ZC�ԉ�S���qYA�z��B�`s�h���u0�^z�$��&<T�\�{���z���^|�'��COmZ��ݏ�g��F����t<�Ēg$/�w\��ǃ_�j�Ln��׍�Q����:O�B+�]�?��	c�҅��ݜz�؞*��6�*rGQR�җ&����|_��ɛ-���N��=G(b>h��X�D��ۚ�@[�
�����?�vꒉ�� ��77�~��i*����9 3-ke�G�d�2��o��H����o �����j'��/�g�/�u_�%O3��/���ڀ��yS'�D�T����`��E�g����A����a4'�7_��V�������>1�����7��	Iw�)��_7��
��bnͲH�<k��f�cO�l�h���
�a.~Z��:I�pg���<�~.O���}7�1��F����X�����(of��Ms�¸�Ê9�N1����^��%��ɸ���(��("���j=��ξ"�UK؎�-g�c�eF�1ZsdaKe��|��5͵���i0k�l�N����"E)�#���ngc�9�6hD�R�6h��卂��+�*��q9�f����{��o�RS��^hY1Kj���e&!Ø���4,E��S��'������'䶱���d�J��\�ظ���C�-��|X�	Lϑ�k>c@4���r�ے#������7��ǚ�Y��ܲ�v�%�i^tЈ��VگG?��\�<�E����Ԃ� b}�0u�˙:
h��|TPц�2P�nI���ˉ'q<y�W���˦�Mw<ư��4���ji�:A�֟�2Z"����M�Ԅ�1�V�t�5j1�&W�M��U���'�vo��|������`�%*K[O\�35�x�qTb"�*�6�!���=�8��E�;�\ [AlnaC�,���2��!�,ZPC��`<|+I'�N�0���0T>��*dm�q��X�"䌾��h��߫��x/g����()����U�h˒����V��IYS�i�K.)��,4����R��`�Ub�[�s/���ɐF�1ˑ0���^�� R;�f�C>6H�ϱ����{ %�i��Y�����-�,9��4�!E�w����6h5+�
�����ޕ�D�xJ1�C�P�4��~N�7��#;�Q.��w6� !�cA4h���%�
�{�D)j����N#ی�C�>t�N#BL(*�,�We�&�(�c�p�@����x_�%���z�Z$��-O�z�&u����M�%졒>��S'�'=�jPx׷qt��G_��g$��D@�P�&8}�|�ȉo��(+JYy~_�����5�yO�����a��Y� ��3����ˁA=��]�i-��7�_����mA�v��Z^�a�)!��9�{*�	��ș-�~���i�*�ddj�U����@q\�5�u�1��D��`^>�1� �):��8Y�\�D��@��m�<�3�E_�Iv��YI"{d-�b��b��'����u	��1�1�%9�Kv�e�ki�;��W����@QQWI��^G]W|�٦ ��k	�ζ�Sg�T&Ƈ9�.rh���Z���G�)2�u�_x�?�d!���Z���-ȶ�^H�&\��Z��:�8o佖�]��\����x�]�8�"G/���/ݖ��59!P�mtT�XF�2�E�M���XMJS&�d�V�P0�BW<�wrs�]�)������XޔZ߳q�iظ *e�G�Y�p���D�ڃ��5�M7`�r�~�;v�X}����dv�P*��ʗc�%͕Z��D�;'
�!�±�o��6{F0aEy����3b�	k���g?�I�e�ߨ��h?�T��R;����~
���Ğ�B$n�
���UPu�$о���EͲ̾e&�_~'�(*g��u�v4)�$L�&B�_P��m�az�ϔ!ؤ>j�=�`=���J#�b���>a��p׈���m��i������$ ��ț3�/�OA�X�ǥ4����~l>��� ȣ�;i�Mm�(g�H�EÎ@_����R�PvY�GW���p<J�v"�2�7Z{�2빴;:n(��i���*�X���,A��;��/��������,"^��4)��Z�.۶�����=����?(?�L�5/����k2�b>��Vs�b=����%�E&t���}V[���_Š3��Vg�:��J>��D��nو���D��gH<����g <���,HR|���3h��	QV�0w_]kǻ� ���a�/E��v� ��;�+�I�h��`�0���ӌ��q�c8���<��{B�Nk�=�H�IuQ��/������}T�Ɖ��5��̾Ug, �n�W�����c���2����Tx����wj"��tKT`%��t	k�?��Ͱ��1��<�ʖ�&&�))��2*;��5�|<=D���0PZ"�e�w���4|����֎
^��������퓮<~��J�$8�~����_��a��)��by��o)/u͐�JZ"ǚW���L��0W��ۉ�$��K<���B@�0N�/������� s�t�����k�s�d~�oCM��RY�V!Z>���#R���-� �}��4��B[�Ao^�Ԏ����$��'��&�'IO0v-B�ua�)��d�ӏ��=�'�{���[s��e��/1�]ޯ��λ��;}ES9�Rt6�����DZ�$�zA�QjZ���>�t�n(1Q�'�QFW�<AQY��싃��/�A'\GI�E�	e�Nğ�hv�_qSAi�l�0�k���, ?<kҦ�E�����7�*/�4z6����8F�	�c"���"[�(������3�3 ,��?:v��+��d�v�ܠ�(��I\���b%�����:^�8Q�ق����O���\��.U�d}���S����ݑh?�fHԾO܉j����@jx������n�E��!�TW�S+B�γ̳jXKE�0�bړ���D��Ȳ:s��e��n���a|K�������o�*VH?�����:�3B��~|��ʷ����� $�rJz	����P-���S���o=�^��'h�� ���5c���jyG����m���
���|rNupJK��K�D/B�v��#*�22D�-���˼���ʑ�<^�%��q �����e
7�ʉ���W�)��w�7�|���&���'��m�Wa賯ꋘ��>$����X���K/�:ch놨�ĵ>��)�|��k9Î���j�z�4Q�ˋ����c=6��	�x�����ƹ4~������1�N) ����O����\�?~�d�G3_*���<�kmX��7Y�2���Fp��(:�RD0��F�٫�Pr~�"�qIvbN�us���#��t7oZىaEa��=[�jB�M�m#��c͌����B�(�?P,�k,S1ۨz0~;K]��K�lVo��B���X��?����$�q�ylx�2���
��hh��?q4j�Ұ�P��Ƹ;��E�����8�c^��o����K3 (�H6��ݢC�\zI��hQv�N����A$h�2�99 1����R�e���e9)C��,P>"�g��l0Q_�n,z��1�Vo�ɐ��!e^�>ӂ�;j���0�� ������i\C��P�=�����1�wЮ��.��f�}�@C̘����SuD��ݚ���ҁ��c�]�~�8r"�����ԛ��u9�v��N3����"�T��U�ZJ�"����ܢH_�!�z��w�Fm�+,��+��JK��U"z/aC���\��E+�TJ7�`�a�C)���dd��{9�P\�q0[�x}���L�j�Mr ���w�ak�#r���a(�](y��>*❍����=�������'�x� �Em�Ҽ��\�Y6�����$`fU7�q_��	mK,��FSO�B1�����5Q��6b8o�%}�����סǂ�7$��f��*P�1i�*;��ee0����&����Y�9/E����ln�dģ�&��#��߯ɧ|dr
YӰ.�����g	m��dM'!���.D�ᙎ���%_!�/��Ä�v��]�Շu��p���J��+�!'�@�$�_m,N����F�W4��5�.�jƐu�o�[J�&�S`7$�;E8�`�9Q?M�xi��DX�H�42o�&��i�*�̼���d^V�6����&h���T%OǓժ�����f��A���h��J��e�8�¡pB�3=���o���Gq͖ϲS�!��P�%�ǁl��'�s?�7�œ�tD�I\w�&N�^�������`~},�/IǊ�"=jk
ϕdx1/����4e��u]~BB��*�� \{E�Z��je�{�s98�3I��<zi�O�_}����*��� +���y���.�U~��h�aj�O �z�����|Ǘ�{Ҷ��V���$�{�ԛ�U'=nz�bMv�[hn1�`!����N��/?�O�r��V� V���6���0΁��PD��^lHJ��EM~GHo����U�E	?Q:en��ĽȌ�AW �n�?� ��2��E}��-	�?����.�6Z��A������tu��m�S�������97�z3�A�3�����e��Nk�o]���ض� %�������0�_B>x��}�>_�w�O��*ŗvOQ�R�(k휄�Y���WԌ��������r}i2�٠9	B�M4[���0k{ �h��t���G+��l,D�������u>z�w	�n5|G�f,��aZ�9K��r4����<�&��������r��j#����|�ʐ�� x�7������0M���]-M?�򂦋ToV�x���Æ��@�.��Š/=�H�/ ���^*�\_�^@�i�eҹj��b=��F��2��xC6.����tVfq�}+{�o��Na���2.ؑI?�ӣ�4�E�li 9�n���L� �_7�&��80S^#Q������6�%�)C�g{�1���꾃}��%�v$�W�>x�k�y��k��Ǹ2Jv#�j@	%M�lB���;���'��c�꣯*[A��i:m��9�pְ۟۸�w������$b��(��$�}$�3�G�Յw�Y�4]�7bD������y2><�{�ֈ<�hL��w`P�>t,Sw���k�:*P��.�v%4F��#��FΕf�F�B��o����E���������2�pFhjK1�/u�n��jw^�2T�K
S,0�!�1��1h�[O�My��p8C׏;����m��M����Ht��U۹�d}�;m�Ǝ�8������܇b��I>8ƈGW4/���/28���ɜ���@�7��Z��,x�Br�ox%�$T*UE������u-DD~��<����,�w�8�]Ǉ��h^�[��s��oy"�!ۘ������ �꫽�&"�l�T@��S��`�Q�B����<��d���Ledzv Ղj�8��wz��oH��E���0�!r&�<���������
�J0j1�buo�Q��<�<���~�M q�ܸ��b�t�A�����hm��Xrj����ū�NPl�^�H�����_�C	�M!e���wR�|����ް��-�Ƥ�����{�/�E�0����k%ω�� n��Mgn�a�ג���"���p�;/b:�I�b�OAu�ol��vj]��"%��R�`�1iQ���6��-���H콈!��NP���rO�=j5��0_��j�U-�ƈ�r(�%ߑ���W�6Z�w��c[�^"��2��u��DUI�~��~�f�&�����v u�;"�)��_�ɗem�$������޹/����5�zü����!�4]��=�i&�@���=���A B�=��4�-�A���M���Ϧ�ih�7�Y����C���+?l#�=�S��x�A.z�����lD>d	H�u\�.R�tH��X�GoL��|��T0mp���D����2�ˇz��� �i�N�Qx�#xG	;k>.�D�C��v��m����Xe��[��Lsa1��S�v��@�%�41jW]�O��ˇπ).83o%�KPX!Ν,ЕI(���ԢJ�28u�^��֘Ȓ�]/gO�<7Ց����vQ�*A���H�:ľ(�:��5�L��)���E������������J���V�%������C���쇫�qXk�D�%���f�>��=�PV���Jt�e�민y��]VѺ��,o|2��Y|$m;Hۗ�T�dCc����L�S8s�A,	$ݲ��"����O$|�~l^0��z�Tw\�B_`��Q���еQ�e��g�G��!x��tw�k���{[�� [h]�:Z��r�	W�2�˷���q%� mӕ����/�6#�d��&QO��@�K�%Ɇ����ÔIY���7�{�83��nrUe�5� '7�>p�ݙ�v��G�~��1��c�-�t�nMQr�&��'����&a�{�)�K@h-�,xʭ������e*��U�T�'.�^��;�t�Z�v��ge�c�)^��
}c��jzJ��򌼾N�xQ`i�jO����c[κ� ���D�1 �d_C�Nl���������'��瓺�Q�`���@/�[Wb}��wFE\ܵ�r�_jq7c��Es qfoiz��WpG��̏��b����1B�6`���E�����_A���MsvS`�k
�sujGv�tbl�I���W0̢�YA���u(a$��C�������ǆ�]%	_���Pb��	cȁ�5.�K87�5���f�ѿ�zU�W$��O�ԅj���o���|mƯ<��-�{.S�4��ۡ��خ�Ǳ}w�Ҏy}䅁-O�.k.�m�5�io�)��%"��u���F���WX�4�]o)�Gk�zV`7��DG"~��q����y�6�� �	��p��b��U���3�l��5�w��r���u?$k�	��]n΂ٲ�lH�:��v���{(8M��&���1/�g���L��#j�u�[��{��\ݣ~C�WE�8��̩ޓ۫_��Ef�� Ǉ�V���t��4���	�E�7�EY/i��T���:xʿ�}�jo�o��~E��hy��8�]��a��@zAbҔ=���L�"����e�}=��uw��x �o����K��S��/�x����"��	_b��̈.���	Uw�R��74a����n���qD��$���-�����ܽ��hh=���
���򞣸���ׅ4�$Z�� �N�&�?���x���]�P�	ǈK�q��O�m���L �;����x}~{&�61�hT�)�H��t��ϸ7�4�0�{M�W�54����}8d�6���Zo~��q�y���Ď����j��҈L���*�&��]�������繱r��Ѐp�C��� ���d���j	�"�n��H�j�qKh&������>�p��g��p�k�:�ȱ6��y��O;��]dZ�G�J_[�*�*������ ���2\��XZp&oM>�1s,n ~Ka(nD�º�����uxi��ĘQF��t�7�i���"6�H��0q2���[}x-/I�8��{�I���8��&��> �a��U::j������I�
)~�s�R߈Ǚ<4�H.y�;2V�k�=��|M�6��Db^�:��ۆx�Oa�+_��S]���T09�����(&&ҬS���.S�-#�,�ԥג�~T��	�����ol	�/w����a	5�x��AkN=��Z�;��r��5^��8����ɷ-���.���Gb��L۽wPD�fF�Q-U�X	���I)k�y}����!�1��ϧ|75PO��@P�E��b�IHI�OT�&��%ew*C-�{%�x���UM����Or3�n��G?��Cdq�S縠-D�K�/��3mA�Vҝ��%U�הz0XE|<���=�������ܥ)��)|���8���u�r��3Zn�U�<�G��]x�R��W_����2��\���mt�eG�������_��Hd��\o� �{7z��CY�Nc���_��c �Z�I�>"G{�A ׼��q�>;����z'!�	��nu�mW�k�X�z��,m� �^9 d{�"����1��o�tJшaMP�P{Â��uP�Zz�p���H��8����H���9�L�Wdp��m��{��<SCv�k��y7�4�oB��q��z��]g��8�~$8��;M!��aj�h]VҲmZ�:�bC*���.�0ͺ�cvl��4fL	\��g����|
0��Ja� �?�k��y�6�l�c"p�O���(�^|�6"U{ KD���8E���f7uE�U��~4�|iI��A�m�qί~������KRMs�@�]dbj?K�	���~�#f��iӣ������LԞ�^��3
�!�k�W(cv�Su�N�e�2�m��C6Eٯ�p	-���S����}ts���V�œ���nf`٧[Ɋ�����}pg|��O��ϯm��^�T���%"�_i�y֗�>�ϗ�:1�m2:�ZY�/��1�/�ɫFX��zFn�2�i���e�8�_�dǱ��__��ȨW�~`ߟZ�:Y< �*�� 7��
�bT�p�͉�rf�h�u+K�X3k-�I�\��#S6.�+���oq�)w���unf���~�e��E��Iw�X�%��s�٢*�ѵw���e��3���>�\"ĂtԘL{�%)^9���Bk��PR�h!����,��;�[<b˙�8\�������|J�[���Z���#��0wK�q��˪�8�w�H6j��.�k[����\�;��\ɢ�q�LtN�Yt���բ�GxP�9@�~�����D�N3������6;n M��V3sl���#@�E
�B'B/v`D�G�r�o�`u�	2���q�@ڶ�ɗ��܎(N����JzpõQ�|+w��v�o�_����_����%��vҕ4(�t$pZ�h:�>�9�"˰��9D/2�`��V���/�/�Vq�XF��'^�L�Bd�c5u����|�Ř����P��4�C���9���x!&ї�5�8{BH�p�RΈn';���%n" ���c$��=ɭ�g�`�-���XIö���ψu�"���"1i�c���U��1J2'�2�B��$�D4|?J=����B#^�Z�(�a17_ap�ɧ"r�U͵�){ݤ���jG�(;n�o+\`hI@�Ӯ�� ԟ�dZty�Ƌ�;Dܖ����u[bb�V���.��`�V���|8Z�� ,"�ݛ8��m��;�{QV�����_��0\�3��x�S<��.5�b���!P�#�7d��w�.k�M��
<�Bג����I��?�����~���� ���֐L ����J��Lys��yW��V5���>en����X�iw��	���'A&�<�.�]�V�"��m�N�u�2MX<�k�T��7���&�:0:z�M��,
��t����J�1����q�\�����K����B�L���_2��[}�Y�x ���	S��aI-�Tw�
c̀0��B�
�ĒFK��|��q�m�64��v���8���/���Y�ϻ��=��u�N.d�G鄽-*�ꡯsz]k�U�Ԭ���SgaA�^f��@�0@�X���ȫ:�n�?'TL���[ta�C�!���_�¨����D~�9P�{��	%Re�r�'�;I�.�-�A ۶�+���0˳]�{��
��6
��j�6l��4���L^��AKɑ����Ja>�W�^��*t����\��i�[L�ܨ�ɞB7���b�S���*<FMn���e�v�Zy��8�1�I����\tA�����Ƴ�L���7�Y���҉8�+�J��ˁLS|쐅����Q�4
��}?���d�%d�,�:`4�-{��Ե��6�,c���j8���w"@���ѮjI!���H~4_�6�b3o��F�^�����Սvc
E�M�s�bľ����4:�W�!�d���@�Y�|�1s�4�����d�2X��a���@��Ygy�M2|�JY�1���X�Z��H����;>���q8�r��D�E�2�7�[-���e����ڠδB��(^�+���'�xd�K|J���,6�s��pe�Kv�jB_��r:�ØNYL�� ���ڸ�س�%�B��9�Yl��Xu~���:D�PK�0�d��}ڻN�f�b}�qC�|�p"FMB��{����w���Ge�]�7ހ��[�,?��?>P�X]|$�����l(,�M�QcYR~`4t�!6ݮ`e{���k"�b��� �����I)e�hr�ey���	���m���&�*��|(�y�*q
�}{ Sv��残D�jɟ���v6d־�ȋ��F��z�v���hOͳ5�b~e#��+�^�ۊ%�)J�P���s+n8�JV��l���Ø��1��rNj|S'�M����m��%���X�hfUcc��J��ά�ᬦ���"��0_��i�U~�e,�ˉ@���lD�h��T��p������xS5m7��x�1�*�v�x�B�yn}+3�����S5s��� V#��xnt�c����4���T�Y���|Ӗs��%]�[�X.�7Uv�I��@�5,���7�)y�1���)��~@?Tw��%c5kب=���k�q�����>�v�ۑ�����Ӓ�TIwPKr�!�<NX\9��Yz��lE87m�Dap��ZQ�h8��Ly�jq)B�I���[� ̭�lտ#�� ��$���C�瘉�O]A��I]x��l�,��$` 0�!��)7N��	�g�7�#�k�g�3������lvz����I��C\x�\c�L���o�G%teμ� �S;ӈ�U�X?ȧV����}���v9�N�mK핕bw
��P<Բ2��CN�*g���`�
��������(x�}�ÅO�TLX��T-�CO�ْ��Q����?�Y]�r櫰����д࿑����P���X
�[����,�y�AN�+�����V!������K� }�[3�M���@��=�ȳ�O�Y]8p`rG�z�i���r��o\o�S�q�QP�c{����-f�LL�5)�8�ۦ�g�� ��RiU��e�&C֕n���:"�)�f@�[fz��6_�*Mh��ְ6D���g�R"	긚c�$&�ј�P��N�7��+G�τf,,
ŉ]�*2�(�=�]���w��N�����A�`�{�	�2��<��Xe�.`�]���&e��k�>�K5��"n�d�$̾9CG�$y]�o�V�p� ��|:�x���mV�`����H�ܓBqOj$��^5e��	:8���Ѣ9߻�G������ޢ�q^Pe��\���W�� 8jt��p�q-���F�\� �z���z�H,�g;��ST��o%�h
�����5+̪��c�ف�O����c��]��t������~%�2��y�&���q�oG_(����:�-�9X/
m2�����q�ج��mp�s��4���8������E��+�Y�W#�_g�I� ǫb+���&�{��m"8�c2Hv�C9��^�
I}l�Ph���p+�%+Y� ��:��	/��d9v����z ���@�^Yoyd���r��kϴov��3���j�0N�{)�T�~��g�H��4."jcO�˨�A7��S�a��á
���
\9%��݉:�����C!�(jߦ�&Yȗل �g�N` ����"+ѐC�.�cw9�4VI�B(��`��:H����Hm[ҭ�ǯ���fT�:ly�/_�d߱Y��v���nA9�_i~p;F�!1k_Ԕ���(5k�ݍW[3�u�����E�����(C(�s>�	�p8�Z�!�qv��GMZ�`NV 
�{�����3�ќ����#�;���u[�o�V�[��D���D��뚞1qS,T��u_���$+q8ɹ̷NΕ�N��Z�2�15���ש�Jp�� A�D�>%9�-fJ(N;��PYK����v�gT�Qԋc��]^���.��Mfރ|ʔ>*���}1�i^N���n6(4���@ӗ�{p�:����}]ƒ̭z#2*{�;�}|덤.*P��@�!P�A�(I�wn���}�R�t9Wѩ�};o��@hp1SC(�=���B���]���7}�?h%���Ӏb�Ft��O�=�	R}�k���%u��g�@5"�ښ O?_"�q�|6��W4<��f��p�h�m5��Wk��$�56��s�Nk�,��U`Ŝ�0�6�cE,��fk	o���T������#�w�:a\M<�ܝ�|��+�2��[��۰�F�%v�ٳ���3��/�D[D�Jf���$n�XF��B[�����8e7l�
AV{+��8f����!��9~m�G�Mh�f��o�r�ܪ3W[F�LA䔾��
��M��D*�kfB��\�	^t~X��!�9"U�Q��H��@D���5E1!c*3����SOw��>-�Of4��wW~f�G��ML������j���[��Sّ�t��<'P��24�E����P'�Ƶ<:=���蛸A����Aڇr!ܜc��"�ӅhO��`ѦZ�3�1]��Ͼދ�'��	�O �l��h�� �@��#�d���9qo�L��J�������?��M=�#��,�>KR[�e�갂�`r$�W��'Zئ2=d�Ұ"�Sz5!�#Ƕ�0F8�i��y���?n��2�8�]K�-5�*�����N�&��e����0�f��ެ��;A%�6�a�_��6�(Vw���s�`B�[N�Nm��,�6�?�w���2��B�J+��:?/X0`oaړ&��y:��:",��u� -+���ke{�1�dcC��فṝ��؞~_8s�-�58���x�S�ҝ6����������9�p����<Z2��u�_��ɬ��F���E�����:A�v,g��Q����s��c��w'b�����HK�@,$�#����YIz<�����"���8�u	<% }�N��]*��v�C�h�ʦ?�6(�'�����$��aPT'�(N�л�L�lu��<r�[ۜ9��]5^�V�(a�a#C@S�l3۪)d}�GZq��-Po����~X�I�:�ۑx�V��{�~��LT�T!����l3��N��\,?���2F�tCa�"k�נnDja�0�hE�U�{�?,<4�ۿ�W�9�İ�m8J���@+���b�Y/�����{3� �dGZ�cF��䬄f�s����譥?��Fҕ�R\��V�����{��ĉ ��O��T�U�'�D����p^2*Σ��Ut�������TduđLZsl�������>n�k7�
������؂-�6�B��4$*�"p�)U��^Q�A��P�x<��7����9�x�� �_�v�U��,?�X�.�d�1��ଠ��S�P�����zE��t"�O�Dsd��W�9��.8Z}O�X��[<�7l��!cpe�6��9��,����1�<Х/��`������cp5���"Qq����c����<�����z��.�<#�0�Q�� ��c_d�&1u(T�Y7^��X(Ŝx�w���4� L�A<�f�2���)�&#.+1��$Gz��P���8��w�)v* 1|
�j\��\�:xkT�a���L�Wє"�@�:6$ ��A<�N���������.ZJ�����L~\g]D`b��8��s�ftm�+��ee7�B�OQ[�k	�ȼ-XQ���v;��,/-����.�~tɝm�L�-l��k!��i�����b�	B[�=r�����W 짜mE2#� �Y��l���R(��?d��-��e|��+�at�y6]nk;��e���L	H$�B�2IA�� <qUt��ԋͻ��N�\��0�ש�+��}��l��(��ϸS&+�/�~������%�+Z��(���Ze/����f��f�OB�5�J#�^'89��ϭ�<.¼��:N�vvJ��9xX��a�D.}�G��5���T@ė�K���N�r�ӑ��il_��R�.k�O�[2XY^/�u�esN���q�q=q}�9u��v�bLp��$��㾜��][un��ȫ������l�øUI�x��x�!\�5.�(=����Bj�
}%]7#�H���8,T��q��[d�Yxpٵ��E:j�\�k����B�sT{v~�X��Z����r�Y�G[��Q�B�&̧��=��\��+ʹďB����ZrA1����IrM	������u�����} ������G+p³���j��ྑ����l�YV)�gj�!����*v�g�X���A�ċ/UB��[��e�<6�>tHA�7�o�H�������^��K�]pYt��(�o5д�?��R��% �4�)D?��ԉ��j��F�0�G�66sS�+L�A�n�����gO�`Y.R���sb�N�zP�sP�[v��B+<��Q��[p���D���^�%U�Ա�su�j�y�V��㜜�m���:��K�}�PΑ�v<���l��(����z~t�;x@s���c�j�v	|��O�]SܫH��� X���[��ޓQbF�WH�q���BS|�֨�ENRԓ�5����Ȣ���D�ol��$�^h���Ӡ�^��朷��b����
��3����Y|x��{���5g��BT
<�bL'�n�ܲ����*b4���c�������3���ߢ5���k�Z�id�aB��8"_�X�
��|����R��ۤr��qpi������ދ�D��{?T�`k �MT�Ya&��tԊ[z��
��r��+��T~��J��F��!��8z�)d���h -���Z�	eG{n3�$�W��4��!v� @�#���Q�r��G����p�Ò����<�;��m�d�yN˓4�(ʥޡ��q0���MB���4���i|KE��������U�O����R�80j]ݣ�o�[FB�WK�O��l�r��^��)C3�J���G��u��yi"I;��9�o7�Ob�W"��4ݚ�a�n��:}��������"0\pM���]��9u�-��V�PT�p	��A9����ɀ����m�+x�%�}#7�l�L��~�LK��Y^�F����D����d'G��C���򙻷����Lo���� ƣ�R���7�HE�M
,	�<OV�(�+�)�w����D�mʕyXq���{����NW��U�b`�8 ��x��D��]*���m���ui�L�z�D]��'*����n4 EO�vЭC²��c'E�Ho�o�����ا�[
5��c�@K�_�0iptKЈ�]�'hn�XXCIv^�ߢ��z_��M�@,1(��Q�HJ��	�hv��5�!�̕�#J����>\I��u����7�����P/KQO2��p�s���QX�)f����[��2�P2q����'r��a�4���PT����\�=e���C�P��V#��T�!�������|�+
�<M�%�%��Q��,[2U���}oŲZ ���i
k���,�cpka�rG��d�,L�]Ս��'�L"Wۚ4k_Oά^B[{�λp:��0�{���X)��zX�}��X��'���,t�7bu���4��>�͑נ� ���DO���b�K;ɚ�Z��,u����eP3�?P�a�ހj.�Uo�8c˪�F���/z����Jgeڽxf��o��꽀0�����L�s�P�݈J�(�B_߾�("�s� �Ź4MP ,��.�WI~*��
A�|� @m&�C����n���Cq��N����N"!�<��*
��s��](�2˼���9�.番t�=d�j	M��Ŏ�Ş���h�
�Y�W�s`��9�5<�:��>=�2|�݈0}�󔣘a�*��7��x���ݨv� ��U�����]^�a�v�>�+�Z�w�(_XRe��"��D<����]�SѰs��=�S$�[)��;���W)&P"�2�Ho^��uGZI���>,Ȍ�c��i֋���,P?��#<�m�O�pd�b���� ���y��L��Z7�Z�k�fC�$�!�3�H���1;������*���gs\��p܊7�x��*�j�N%<�=�U�[���M�o@rzU0�����v{@|'�8$q.Z���ʈ#e��������o���*����R+