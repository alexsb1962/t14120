��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��]	h8��`��(	�t�3�����U���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍C95^T��#� _�_Ü�@�hF��W��`��q�©��ല���?�;��XC��(�R4�K��b1Ø^���#K���lӧIA�a�V��R�5K�yQb�I�����
J�'�دv)h�V~�$v�p��"}�vo7k2a��pP.S��*����طǪ�`DY��YH\��!���1R�_ߥ�]��4�:j�l�,9��)'��e�Ni�H�f���Zߧl4���0�?�1~�x�c�	�L}���i�m���w�*��O0���G�٘�*"��� B]�pE(���B��|�(����5�:n�|����Z=%�N
x��]Qu ���������	x]̍��;���J�7�_���0rÑ��W��s�!5�Edɲ�<a�r��Ҏt�6��HPW��es��^y)�k���J�ҳ&ƵY�h��Ώ�4N:w���.�t�^6~�@�����k�8���҆�|n����0ӵ�;r|@�b�؃��em�J�Й�m��JNu���]�ߏ��P�umSe��S�2�:,�nr#�9l$�/P��pO�c�c�ENk�lAc>b�G��8̀@��k.�"SӠ�|&��c���m�Rܙ#l�%q�M�4�}�����r�N�Þ��t�U�PD@��k.͇�@�L�v���0�Rc=���T�1�\�^6uk��~1f��t�jPP�K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s��e�IC�_�\H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���%	v3�t�  ",����%H�$��ī�o��<�)�G!�u�����!�M��Evl3����SO,F=d9�[l�&��q�©���H��JnXeS5H�j.F�6�Z��'iNؙbG�Jlf)@̲#�G%�&0ĳ]o��in�m��+o�Tku�����F�N~Y�����rYd�ea�;y� ����t����M��҇+:|8X����\�v�T?�7G|`�UxHj,��|��	��b9����pP�o�����\{F˯�+)�A ��E+���XP��Ȩ�wl��h�Vx�%L��ʐx�?�'n�^0op40�zɈ�����/�U��֜��3�b9����,����dj޽����3i�z6�웗���JU<o^.K�}�$;��션T}u��Q��L(\Ӧ�$�̎�)NC�lԇ�-{��E����F��j��\w��0]Y��
�iC!�`�(i3N�By3��<�]�!����M[��Ǣ�չ�Ad�!�`�(i3c��Et��q���U��ꢤ�Og>ݣK�6<o^��Hm��e.��xu	�n�-�6��
�jW��D���M��ҹf�f3'��$Ι��o;�¬pX��g��U-�e�,���6+�mj�B��V%@��4��c��Et�Y�{'%s�[�&B�踫g(�r� k�|6�8o�`�_f>&�&i�"j���b7|#9���{k�h�+|�c�$�t�Yl���#�]�!��M8���	D%��_�ͅ��/��=��K�q�?l�_���d�uY�ا�W��_�ړ8���/�I<��f��tN2s���(����5�:n�|����Z=%�<�/��욷NË�����8��z{��E�EYZ/�矘��-n��I�?g�f��u�H(�3$�����"�却G�(��]��JX/3�_Ge�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cULjaGkƊ~F˯�+)�"j���b7|#9�����)��� ͢'�����t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s�h�v��T�v��1���6��	���`y�����g�,P�n�BL�Jx��e�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cUL�f����Y>1�Z���=�"j���b7|#9�����\�I�N�_V�/�O�	McV�6IWJE�r���秹�3I^�v�V�jQ��gs �\1�Z���=�"j���b7���Øf}�
�?�?KYC'v��@B�IeI�#�h��/`�㎏qló��@d���/��=��K�R�hE!3�͸@����gG�DI߃�����]Y����`�)�	�%{�;����f�kN�ı&l����[}�@��L}�
�?�$���]׽�kvo�Apw�I�N�_V�ܔp�l
d�R�.��On��M��ҹf�f3'����q�f@[�=�5x�>ݣK�6<o�D �ks�#�h��/`�㎏qló��@d���/��=��K�R�hE!3�͸@����gG�DI߃��S�*;qܛ[�l\����	N^�U{xN��i>r�<Uee�,�Aٺ�H�L� s�j8�	�A��ԡe���b�kvo�Apw�I�N�_V��� ӌIE���`�z��GZ>.�02�0]�J�ȓ�iӚ/��i]��i7N�_������;��|BV�y}G�2ْ��4F��u�Y�KG�ξ������eiqb	��G��W+��W�'G�+R���o��_�Rv�䩲$���dS@Ɵ�od=��¾ȼ;�jmT�#bs��2[�a��o���H�RtV�^��TBd��pS�*;q��=<�6>e��0�U+�qbp@�!�`�(i3mj�B��Vh�EtC�<�b_X�XV�b�z'hۉ)��d�7�qļmJ�0�6��Ra])n#�璓�c�������t �[l;[�G���KlG%��`��ǚ��ظ
��@�U#;�jmT�#�,l����M?��y�!�`�(i3��TBd��pS�*;q܆QCj�4Z�_--���gz���M�~}!�`�(i3mj�B��Vh�EtC�<�8
l]]y�1hPR����p�@�VҒm�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ����PJw�R���y���,!�������[��M�����y48{���@2P�)�#�gm隦���W+��W��<��>���-vR���B��G���S,��!W����GS�*;q܋�DKY��,Bp��S��.�g3ZE��g�Hb �;������f�q,�'��	%�qȸ gWVbT+�,���XF:��GZ>.�0����ڀS��d���!iM) �D��U��)���Y;e�iKI/B޾PԐ#��go`(&�L�xjzӝ���I(͂��-����8��;Yv^�-w2M#-5�{_8�Y��=�}�Vݨ��}Dq�f��Ro�G/]%�z�-uͺ�s�η3G��Hb+�����;y��v��\���
^�ݚ�Н�y�}�6f&rG��HbSz����ʪ���l��1bx�cF�����Of[� ��2�]�<�!�`�(i3FwZNE�&tS�D�'���Xw�j�7���W�6?���_--���g|�m�ߕ�><���@��`.��53���w�@V[Z��.�~���Fz��	��x�ׇӭ��V�Ո��Ú�'nB��!���c�A�L'�ɻ�L�1p/-�������?�/5��"}P"G�wk�:�_q�pWS�*;q�=�9��tsȸ�"rR$f��_Ub�F�S�1 �-��ټs�  ����'�W�6?���_--���g|�m�ߕ�><���@��`.��53���w�@Vw��뱐�
�:qEp�;�P�t�5fĉ>99��A0ok�׹��7��~���-՝-xC�;��|B#���rM�J�̔�8{���@^�4���z��Xgjn3ԏ�W+��W���#� ���u�Y�KG�ξ������eiqb	��G��W+��W��u[i�>��W�.��A$�P������5d�`UNP�d=��¾ȼ!�`�(i3�'ž1�|�'����u��r���2��}��1�O��dN�<@Iv��nt=:��:5A��p�̢k���"��w6�0��ɗ��zi#Y)M���Fe���2+m�7m�T��Ʈ+ˀa��z��2�,;�jmT�#�,l����M?��y�!�`�(i3q�\E��0Z'pǘ���Z鎬�������(���fD=����e�:5A��pfĉ>99��A0ok��fĉ>99��A0ok��W?�;���⾰���Q$X��HN��R��?�d���&����s�iV��	��y�����]T�
�?B�F�-*<(6i��ƫg�T/)�ѹ�;��|B���MRо+�-���a��R'cf��w��/��=��K�E��{#6�a?�d���&�t�{#	�x�u�x{��̷_��yC��S8�f���g�&l�p�q,!�.�g3Zdj�t����9?�W�.�g3Zdj�t��FĮ�ͱ��Jƨ�Jt̫j(&
M�K;��%YM�	�v�3� k�|6�8��:�EB�Z5�O�%E#P#L�
�am$��	��#�|����m�I7��-55x|���MM
��,=?�d���&�t�{#	�x��_--���g�QF.��v{��lw	�����?QZ���>��,H/������,�ǰ�������Z���zh�#L�
�am$�Z�^��h�@^4KT�v��1�5x|���MM
��,=?�d���&���=����t 7�J�[> a��M����DKY�������?QZ���>ś���k�����,�ǰ�������m2�
��E����,�ǰu!�OO��
}Z8/��RU��H��<�C�Ar��� ��иܖ��A�.u�r;��|B
y�3~;�>g��4� �㎿���o����E��C��5�%]����8�B���ow_;O
�J��:����{k�h�+*J�X�$��+�nj�a�0r�uzZa�U2X��������,�ǰ�������� 7�G�Yw�R���yWp�K#J���.�U �3Ah	)ޟ-�b�+�