��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����k�8�%j���'ex�c��F�WYڊ��^�z�D���)��8[�� ���;h���hPI]F<o&�~0������t~ ?z"z��iwik�a���Ha\T��Lo�	�o���7�]�|$0��
�Dۖ�t<A>����9�""�>/��Y�5��6��%���(dmO�賩�ҫV�4!�Tb\�Ⱥ���_�g7h�)���ҵKh����8�*0���"�ކ���Hi�_��J�l_�k�����,���v��Fb$��rЄC��){��(�ϝ� !
��Tk62,�.v3����rzu��ώ�]L��l��~S~M+ډN�	#5jZ G�:[�j��_jB�m�.����ӓ20�S�|�Oݠ|��c�,;���JQ1zL�WK���͹��e_� ~�r���ڵ�x'�;'�������\:�pcT&���m=�rû�{ؒ����[����
]+%#G�|�N#F�\O>����&h����Y�q���Bkb:��9m| d�ֻT`��#�7�n~����ZH��O�~�,���I��F�/�2H�9��b�5���?Iy�a��ԹimŔ6�{�,�nb��P��J� �֝i��t���;�t�����>u?8=J̱�B�?i2Bĉ{�q����@ǝ���r�߂
/�'���IJ��4��� ���؂6�U���j Vf�W�o�v=� C�Q
�Ax�>��t�H�>�/�_��?�} �"[���xv��/�q��3#٦.��1]wf��b͑5ׯ�@�b���/����x�X�t�65� �OY��SO�l��:� И��X>h�����z@��=��I5ᓂa�xBޮNM$�bc�w��*9� �_x1D� ;«PD�鸶|�W�q�����E�>a�-�yԓl�zW���="G�o���)q
�mhN���~>��vx�*nC�g�,.P['
�a96ņ��Z�EZ���;�t�~`�S�o.�PQ�\�uQ�Cz�%	�L��])���6���!��d(s�������b�=�1�b�D��>�%#1�4�x���јc�P&� �ti�͎�|�f9�8�̌k����O��]��;4f�;(#1��"��c΄��z�i���q�e��2��x��4��n@7m�?���C�E���q���[W���&�1F���#M�Y��[�����c��G�ٹ(/8��vSp|�\>u6��d$�k0PiD��<A�&z�&a���P�tʩ�UW-�[������/-@�{]T�(�yZK�'y����!�԰���4%&�DDQE��/~��VU��h�dLz���;�Ν�v�e�_Du43jU�^;4�=<F�z�<kW�"�3'p�8�bs��%��*\*���aq�������:��V�9���4�'��$�WmDM%�S��D֗<>�e%���(t��Ⴥ Y�IX�}�m�n�I�%\�c[��c�z�2�1D�f@z�L�Rj�z���g{���i�h���!.�t�����M�.|���˄�����d�9k�}rqx��߱U���90�3��A=�#B����G�"�@�'Tr�g��E���"{�Fr�
�s�֯~۽��i,�yE��;v�9��mM ��XR?�c�~Q�����D�?�dK�1���Ȓ���h���!�lO*x�w_�m��	�g�gy�k���N����IM����)���Uz��(��^|���b*�fcC��	��"z�kE���W�B�˟
DV�s�����봦��
����*�biQ����w�Z9��_75�;�V
p\���0���V��ih��ΥE�r�]LR�p����#������X���4���5��`n���S�!Z�m?lsV��x�[��
n#ad��x��%5ʑ��c�2Р�����D�%���X�3iٯ��d��T�T�b���tB��/��'�}ȭ�ɆI��!X�� ���2r�4��g���;=b�y���|r��6���N/F�ɵkb�y�U�d����N���;,ʓ���%��E�Yנ)��H.Ҋ�9�@VD/~�`��O���
|[���9П�ݷ?�'��8�����T�~�%�jN�<Y���^��x���б�c�7\��yj����G�3,S�JN�/.�8��~�LI^���|)C?>����r�ׄ
0]���p��5�o���O�Q ��thL�ֲx��S���Z�m/��RNtY%ia�Sc��Yj9K�.$P�M�g���K�?0�j�ofs�-8{���O�x�.�F�蕗L͸2�m@��;M��&���=*��O'!Y�} M�:	�8��Ȝ��y���	�� �<�W��La^���]��Z:G��۔E�Ct}])ubwP�f��W#��%B�˂KB�K��:Ó�֨�F���I��mme����A���آub�����(Y�����NM�2	���6$�#'T=
eP������R�N:Zo��x�V�Z�z@�"V�����o[zZ�"����yC$����W7��l6Sir:���|�6��g����%K˗�[�0�A8ʴx�@���Q�TK�5����w�w�	����v�G�(�d1�j�%^˔:O�d��+v&�V�G�bG0fG2�j ���1M�߰�Ս�V_�斮I����8��7�M�*Nj�:(0�A�϶�v�CAv���={�"@u�~��D�_W�_�r>x��a��W��m�L� �	�qim� y1��Al#�\H�J�ɜy����zQ�W@7�֫�n+ڐ�)�˙T-G������CӨ�������b�J$�F�́x�������ނ�׽u*������Mғ�q����7;ې`�0����4	�+S�JA����H&��d�ш4*���O�2�8l;c(TDG�f̪��c���<=�$��	E�C���E�������W�/�cͽ�[BQ���kX�^������Q�%Տ<|/#�1%��d�U*�ֻ,��c^�9�x���o�<rtDc�����C�������t�0���h��l���c ��2u���n~����Eko.P ���H3��w�J�r����"U�`��+M^���VCc����J�G�q���䄨[���S�lO�a]80L��<U^�#)<���g?��~�bx�ɔ.N���0ܨ?(���T�/ش�-ebde/�RV�g�p�Y�2�B�8|�x���q+g=�;I�W�U�+/���0n��@Jq�������D@1�r����q{�$���*c���Xk
�]/	��- 	�o��P`QB/.��B5�w�\�5�Ur�� ,Z|^�L�l�)M@";����J��EvN�?��@qV���C�����o��kD �+����:���S�%�
ާo�5k�
�vBkZme��y�E}ȣ��B?G�J]c��C�7ݻq���a�If����QO�; a�x3ʋ��ƫ�����Eub��c֫�g�\�K��H5��Y$�e����twW;穹����'c��|�y�F�B8�d���}d��Iǰ�J%MNi��}����������9uy/��Q���Ӭ�
#4�� P��վ�����*J@�ez|�v���{���%���l=Q�>��\re�7�=5��h�`��郴UB`��vrL "��Ov�ZksT�/�=�8���:�V���"H�9����7���r��=�ِI��	0��Nm(1�h�aQ���(�%	e^��>l�7��K�`��N6n����R;һ��#�:�6 ,�i�}&k�-�g���]J�]��T�x6����`K��>��|���Vg�G����k�v���g�܈Y?��vpa�.��|��\k�v��؅@- �Q������� '2c�D�q�����j�W����_	-���FE|��Xll��y9��ݜ�6�C�O�m?�zň�P�����߭!���>Q��-��8�"�H��wgmP��-�BH����2���(}��4�=��"}׆	��ռ1�S"����U��>"��|阯�];{n������q�z�pf�{f��类�!���0v�����^���'����Z�Y���t�7Ur�2љ�y�^�kO>���25�;���f��çU��.E�t����b0��?�g�[�Φ�W~A.b�����gʆ9�ځA
g)#�;6�ԩ�.D7 r����vZ	C~�X�W&N�?|ޮ�F� rǔ@��$|0n\I��Zl*R�}��ܑ{��a/���5j�
eK��X�r7,���U�,>D�^r[s^����5@t�!���'Ol���V�j��X�O�v��~fEl�y����B6��-4���k��E�kT��R&]���ֹ^�2$�����r�/l��,S/�4+d*K���0<|#D��j>��	��c�1�ߍ|�qJ�[�+_`tU�:��2�c�=����.��vxL�� �$R����<�w�e�+�`�������=Qd�Va@e�6���?r'5�(��{~�!�'4$�k�)A^�=_�Y�-�1���Uo���Ekz������cخ?
��{�I����f�ڑW�G��5}]Ku�b8x,�p:.p�gb��l*GW0	o�����U� ��e����LP����8�t�x�ë���t'���<%ᗥ���~�]6İRD9 ھc���G���I�0<�r����ja�^�!�<;4�<�|\m�z���֢�'�B�!Ӥ�k�ؘ�$S�5e�Zi���)�.2Lq-��@�L���w�JX��#"��O0�NUm��q�*7�=q)��J��m�i���mW���+쬲�C7�t|
<1�m ��gz|r��|�=�"�iPu-Rp����wZ�p��WdTM_�c9ք�T"����p�{��߉�{]Q
�\��Rj�%'���S�]h�k�zt���}��/KC�f˂�.�JJ9�-_��mt�1M�ul�,���t��!���`KmnioN����ZT���������/�?`Yau��/��އ��:x��ɮ�S ;�g:�f�����u� <�����
C~ˁ	��ʦ��R�d�j���W��FT.��;x��fp��YzP��E���c��<�Bvē������r�]䏥~:���3� =3B���8�wu�f�.�`�c���}��vsM�����(C�T�ۨp+��܁�)iXg��츆�o�=���`䏵��Q;��!�m����&"K6�0|X��t�P[, %=Xĩ�J�1%�׋�3����)۾$�e�xS�k�9�U�1e���gW-尐$ ��CZF��Ǒno��
�1ϿT.���;.����.$C���4.
���(���;�E��4�H\&������ƌ� z��}�~�r�!���s�w�! ԧ^��$d�o�bzEC,��3����G��P
/��1��兝;�4��̂#��
��M;�R^�0U��XLٜZ�B��B ��0�2b*�\Q/&� cRF��J�j=�Ac���+=R���p�����	�s� �f�:R�Q�!��۞Qqf�UŢx���ڃ�V�.�fECC���Q���A,�ࢌ-X)�)��ۗ�ӓ�T���(��<v�>��LmV͢H&�-F�.�Ӽ�9x�+���9 �'���*����ժ�Yi�I��e��,�_T"'��b<KcH��3���[�t��o҃��\D䢵���������^�����unJ�٘�{
p4�!���燏�a��.�M�G4ʇ(���])��<� ,.?+\�k����4��t�fUFm:ہu�Y�Yhٻ�3`#�d+�#yib��?d��G������!r��tY
|�%�NGF$܇k(�����}w����� F[�� �D(w��5��V�h/��B~�(w\c~���t
4u&@��v->��[��ƍ�r�=�<03��Ssp>h�Q|��+�����m!=�������/�p�3h9�Q����y����,BNi�� �M�.H�e���o�^���<���M���{�[��g�~e�C����h'Q�M;O�/�vK�%p�~���u4=�w�R�^_!|t�K?+-��F�EZ��A �
OI�\wn^��o�	$���B(�#��j�x���x7��i�������>:��N�a	��@O�0������ˆ۔���X͂_�JVHЭ_V3��~�q�C�m	��^h��+��TԂʻx!�B;p�PF<b�T��Qm��й	�#����-�t�#Nn@��I�pa�Z�g���3�P�[^W��>I'��;�ѲGlXEL�%�(�y�b�C� ��I�?���c|�LRF���R�Te۟9PW_`2�ńϋ+��3`G�t'��DN?	�Z� ���_�F���fX���=7�Ve@���>��^,�a`%�G��9�d��4�@dl��3�pP��_�Z�_��cƻ�#������[�����L�bl���X�ns픯zm�6?'6�����#[�@�ŕ�[��]:��h�s��rZV�![k�r .��}f�X�ߍ������=t	j��fJ	�<��:$(F5]"���7\^�# ��������S�0d��8�4	�vS����ˆ���ϝڋ�H�_��͒P-AM#��I_�w����؋H����}�N���0����$(V�1�|Y�� H��o!l�*�j�`��hP�E*�A��A�[�w��A"��Ğ�nu�s�O�� �2}7�%m����nR
���(��F�����!_�E݉e�H��:�9�S:B��CLm���b�-��c��0��
�7�����И����T 
9�9�j�o�_�B  �A�m"a����\X�~YwIVK0Q�M�|�S�%�"6���J��*�}K���͡�:��-�7�3���ȁ��Ȕ�ЋM�$;�y�+���y)c밋�[��C"y�������^���Z+�r�-r��=:%,��3.�]�n9�\ei���E�ۋ�O�1�F�a�CV�uAx�C��㉌S���w@�n���:D��E�f͍��G��p��Z��b���Z�,>iԛ)����u��;�Gʀ�Nm����gĽW�'�u�8�!�8-���R�N[H��o1ai��Dd��&C�����Y���{�k����_�q*���Mr}.���k����u
h �4�Ǆ�)��Љ���&���A����Yڗ�]oX�07��Ҩҋ����45{�����J��Q}�~ѯ��C6}j ؐcz�n�h��~:�C
���.�+s�s[{���wZF6�3��Y�:]�&�&_
�(�R�:�#S�-Ѥ��So�Ȫa�+�6���,&:�P����!�k�ܤ��|�|d��dD�
�tMu"Qb��P��&$-�d��\]�r��%�.[�ʰ��UkQ��.o{�����_������Y��8��6p���I�����/x�W�:�LyD`qD�p�8̱��<dKxI�r�Y�Ff���"���C7O����V�RP�����#�Ԁw��V��j���ܰ��:@��|d��w�S9ί_��ۙ^��Tl�a#\���^Jt�ldoB��HnfZO�	�=)�3mrٵ(�I��1�s����]��A��r�D ��qJFm¹E�����y�B!qne"��W��������I����n�0�Y�����K�*�hT��r�UX*� O��)Nգo� �@�8�n{�!���1��T`� ]�K�G���h�޹�X9ȿ+��<�e�Գ�:��(Ok�^e#(�|U��������&y�������a~��ڮ	���YK[���h�4�X
q7\��&�C�b���Xa�R(�e�ԏ��8��Y�8�	�P�Q��Ǣ���������U����� _Ѵrn�X�9)ihZ���i��O��PC���vQ�4TV��z*
s�%�ߘ��pd]��K��ڼ����j��
�\���@0�'���빍CTs��ņ}�aQ���Ϳz��5�l�` :�H��Ը������<�k���;��L,��+F����_�@~J�3&�oל�M��۱pwN�ɥy@�P�y�d	&���_�n��'S��&�}�J��� v"�.���z��vNvMn)����t��R�6��ޅ���@�4�� �F���C������muX�N��S����¢��г�'�v
��HlT�-DQ��^�I��^3�SٌVK� F"�[��3*&�uV�Xuc$��r	!��lA��|�r��l�V
�]�$@����@'*:q��@�S�n�nj¶ad��,�=8+];����~���X�\Nc`�h�nHZwY��j$�	H���9��]\��^c��|ߚ�k�֮=}�ʤ�|��B�rj���JT}�-ۀ�q�K��۲�au�0�N�/��]���;a�{�����fyǬ�r�n����� .�i��n�}�g����6k�A�!�����V	���Ήh,zNj���q���s�A
��Gj����$Gi�u��@��[G?74�M����k������?�)k�J�kڎ�+�C�����������%wL���uNT 3�A5�;A5�_���xo���U����Sa"�ѱ�v��� ���\�~�Dz��;aإ͙"�~7��3F���x�^ɳn�#�_h�.����S��qP����"�s��({�`��Ƽ�̐�ly� �v�I e\�->�����~p�̉�**��S�7ԕ����S��<�n��]`8J���X �Z�-+yN[����vGk}�P_u������Ѷ30�`z(s�W s���rS�h���~����[*�o�O�Wz�F�USjb��#�N5E�0�9t��3�*-��Tj��H��@�� ��w�=��lkeD��+4/�`K@f�N�
|�����fr�鰝�V�u�.*i�-{Jk_��'��Vcy�a�=\o�gd�y�Ň����c�ԍe\h4,��Q�9Ӗ�
�#��&p�Yaq{{�qP9��I_�8�.���KV�_��-/��R��l���i�����C=�ޣ��t�B�M