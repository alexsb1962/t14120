��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����F.��^KN|{�H����k,_��۪T�?L���v�����f�G��LE�� _00��~���]�B>5V
�D����4m[���G:������H/���͞2Zk{�^!�8���Y�p�6��A����D)6�LK�C3U��m��U��/�� ���R�[��kP,+�u|��C�]V���q�B�Z�Nv�Cq��E����h>}F�s�ߝ-冻�����WO���vp6a:.A �0�0�[���:�#䥓`�wE�����v|1?}�!2��J)������<�L�0�'��{��>�L�y�M�s_A&.4��˱�kW��z���*���7	0��Ѓ��8Bwn�dS��&%��Uҫ8�nh<I��K����^�F�l��W�jw$��A�&=Smdzd������b9�/���|���p����6��w����/�QH����H�|���9��������c��y$f(4v�?��Ix�x��u�.�6�_�B��9�<T.?0��l���唇]� Z����sR�{�6u�C�)d~R� �Fx8dq�g/�A��''`S�]����ڬ���b�Ӻ=��zՙz�MB�N�b@��ю�����e����#�-��������@��мk3$�UՋ�jя,�}�'-3�ǰ����.K��_�;w�����.z�$�z����"+(_و���&�A����M����&1VwՔQ��h��b�hFqF�	jH����z��#*[��r)c�	Y�1n�\�h)�a�t��Y��\�|��!F��O$�Ӻ;�9:/�w�`]XXD����"3I#�@9��h	c&	������]9;1
c��{&�1����t6���}�f�jC�J.�Q�%�b&@���o8�Ʃ9�Yk۲�P�\�P��_す���2R_�d��x?�3ܧ�)��_T0iҠ�K�7o�V�2��:�XF�/�eԮ�؛�[����?������Y68NqM,Ŏ��
'�"zt��&���k��0��L�����	f��]���0��l��V�c�q�����#ti�7�Ld�D�_9������5��7�Kq�F��{�C:�~��=���R����R��R�V�w��Z��S��%��>��&LG�#ꠓ��7�F�:ۻiH&_ڕ3s��� t��]}[�n�l����EEs����W��5^.Cuܙ������p/u��d7��<����&��i(�◮>�i}]�?* �(�8�/��z	�uܡ巤޻GO��^�w_������ ����R�S�u����_�qZWZ<X�� ���bے�#;�ܣ�I+��}J�g;@� ��k#c��(�֪$1��dw���l�-�O��Z�a��2�����S�1h�Z���1�JN�����8pH)9�m��*���<ӥ�]t}1\��4���7�5���i��ij��6�����a��"/5�UˇP)��bB:+~U+2ě�8�W�B����X(�1�[[#_ڠt�eeG6�DS��±�@,��Bp�g�Uȁ>�iO��O�A�^���
`�k~@�Fsd(��T�������Dj���!�L��}T�4��7aBN6���m��
��[d��Y�8>���|��NY�:�����q��]#e�p[Ҩ�=��Ҥ�.-��],������%�o3���x �H�&�²�v7ؾ����N�Ǹ�h�����PL������>MvY �� ��x(�t�uS8�������f/F�v9�a����������w�s�>�Y0ɳhS�V������^���n�c��J@#C�����B�yT6�w7|L>
�u��w)l��S	"S�I֘���B�Ȣϒ�*_��ТAZ��z�5G�l�is��K����:TT�W{`�-̖C��D��,��������k(�7%5���ـ�@�q�/X~�c}ѱa=a��%C�gL�:8�|䉹T�=��Q�~Թ-��i�{�F���9{��Ik�-TWV�ۺ[�	T[���4~�^H#�Wl=F��O�/��eF����r�T �v/S�Hn0�o�vU� @��UXR[Q��Zt�v��g��?kW��bP��S�:��Y�p�Q�,4�U��$�>Fe��k�/;qJ^��=	���oU(&�_�#68���S�}{V����Ţ:W�'�|���Q9*(�We���1�����5�O<���a�bקS�f�71�9?8CJ��-���7ٍ;4V+I�3斱U�W�.;<�Nq��%P�͝a�j�i����JG"O�7�Z���6�0;
���) <�E]�=�� d<�B�yo^=�ڴX������sZ@)oR���!�.+_�wb���-�.L���f����bX$'�w����HQ�#s���=UB@=5X/{u5,h4�ƫriI�Y*罇Uqn��,���ie�y&�#̍-��s�,z������`<�&\h���RM�Kf9]sS��݊?��������1��j$���*8�pMJ�F�.hh�e����$�I��6�mP	潊�;��G_�Z�i�񇀫��WL��o$����R*��h-�
���~W���K�:$5c� ƫ<�Pnݧc�
	�/�m��ޯ�%�|�-d�W���(�:�f������1�YS�.н�j'�k ���'��q�#�+��o�oޤM�^dL-)��Y2���ɞr�J�>�{�x3�SɊ���S�����b_�� ��N	U{HO���=�/k�;��� ,P�q��%�R���de�!�r�jjN�J⍥?���'o��-8'j�x� [�gn3�^��OvIa��T��`�	�.O��N?� �7���%|�a�)+�v�R�7����4�����/����9�s��m��]���%�*���7(��AY� �R8�SF�A��Qa�6_]§���G6���gA�3l�l�QkY��s��C~ j�"7�c��`(���
b�屐����x�d��S�*�6�͋jc�\.B_iCUq~K[	�}*��Tؾ?�d�K�ú�٠�}�IT���}ޑ\A�x���I8Hs�J�!f���,� �Sq���g΃�$
kӎ�1%�6��]�T���1�b�Y��sq��?��)+�eC%��1�ܧ&�Ǎ�'DN4�i���]r([��f�X*ǐ�:�/*�@�x�J?�*��k9����8�Ln�
��-�|�������j���D+���>��>F]�O1�ك�m���{�9܎D�X=�GMa`G-<�'}���O#�8�l�(�/�*� k��ʵk��â���*���f�$��u����
�׋��#q!|y��){&���r�F�5����7q7u�(����ky �ƾ�Q�C�-�"�Z1�i��pX��$'���>I��mbxm�3��Sgb{E���2vs���
s��ɩH�4��G(̺~4��ʲ�Sn_�H�1
2���ҭ虆�S��o��6]�S|0 Z�P��Y;M\��O�~��N��n<q �K'gBw8�;��FIϤ#�� ����V����'��ܶ�����'�|i@���C�����' ������YFE=O�קU,�㉊�Y DR�U[Tpϔ��B�BS"n҆�*���Q�$��.��ZP�cmV|���u�f��L֯�t�f�>w�*� ���л���O�a�q���D�������PTn��pCvom�A!�G��+,�����CXߗ���7ʃ��Rt"~'�M�C��T���%ԗA��ωzo^�=����Y��E_N���,_h��l{˙G`h�`����"�3u��\��Y��4�Ĳ���M�A�p���m���N��ҡ���3��=} *�[��ѿ)̶��xz 2�OM�S�[RvT��X���5T�nmޓ����t�=qҬ'
d�[��!7��6o�!�屴��"�L�0E��P���h -���1�R�Q��	a*3$�Kԛ�w��&��x,�g���9~�1U.�Ǟ�# e�?]�׫�[���4J�&��������+�K*�
��ٿ�rT*�"R��V;��;�A!+@ dׇ��7�<y4����sKT����a�{K�VF�o`��U�P�E)ķ����]}5���V_`�T@��Ȯ�����F�lM˔�c��`�H�p6�P�toj�; 
P%��I% I8�$�*�~]��n� 0DۮP���ޡAM�!�M��]惓��_#�y�M��2#GPW����>"��oi�@����;���y�$eE�4���]�O��S�V�h�����!U�bG�*o�!����8�� wn�F� C�b08K����e�CAB.��?��\݈��M��3���*�H��k��Z�}in�1�7Cw�����R���j�h��q纃��G�-�Á-��=_��_���S)���#�yk��r��Ӣ}EL�����9�R�:Ϧ[h��x���`�4�|"T�w��3�J���yO���*H3�^p%���_=X��g��4��x$ Q�MQ�Ӝ�Θ��)�j�@#m���Q�uj7Z)
�����O������q9ɋ<������E��-^xB&⻄縷<�JwѤk�ぺ����,��y���1����Oܢ&[�6��^�Vu��HLEX� N� ��5jY�E�f{�]-,6�J���6V��v�h]��ԙ�?�[�#��RJp�&W��S�*�ߙQ�	��&?�qd���
NOr1iƨ�o텲��GPo�:&��s)�<�.O0��U"�-��+Q"Xy��nnW 9/�S�~h�u锜��g���
%��^�������J�����N#!���i�� s�T���|�eA�GH�Dg s��7�\i�=��y�"|a|��|�/������`O	�?���	�W�Xdm�a��Rk�Xg����6��W��[p{��-ݰ ��2!"�fl�q��;�I"&��=�o�>�s��B�|��Qe~�*���+�Ipd�~ ���Y%��U,�h�`,�Z5m�Va�
'#%ֳXX���>V��&�k��U`�^=����5�!�����_'�U6�ۆ��M���(�Z��1��u�z��U[���] �Ux��D���cV"���[���x,��QDUzE�跸��*��)@/��a
�C�_EǜL@�z�:!�Y��[��@+l�ċ�����Hv~-AR��u�H�MC���#�?��'��b����X�^}�c�
�FǤ��q2iz�.��-��@.�r��"�h�M��!�ٱ���i	_X:��C�S�9`�o�-ՠ�4jeV�S����^��\:��q�%�C/����{���Ja�u�1 h�� eb��$)@�ɹ���������|'`�!0�L˥8ih��h�F����5��T�u]������:�S�*A�-\���S�q�=���56L��[mټ���
8bʆ#ɭ�a�g�����&���Y@��1:���ʢ���l���J��9$��^(&j�+�x����|q}3x8��\�zSY�z�6_iԆ�O������Y��)z����	N��<���v*�������4y�u�����ih�Pq��זּ�qȡ���t����"�|s0I�X�.��֟��:�T'9�h��0���d���̀Q��T?O� ��J�����2��o��᝹?�͋�33�>H���,�]#w�<mF��N���<�\1P�7�15)R��Nmr�����Ë�!�����L��]��2#*�HMKS�l�����OKw}�
�+M�ѝ�9����}�y� T�CzH9>����3� ����31?k5M�y,�EB�j��3���U,�1Xop f��BJg�5��r�LD�5�ۼ��r!4����;�!Q�]�P�4�1kP�B�� L\�3ۇ��v�8�<�;
��%t"W�����
(I�ѹb��Pa%l��
������N�[C&�;Z(�z�Ƽ�g� :�d*KI!�(E���0���j�A@����zL�����L�jm��c� ��РZ	']ü��sU�ooߚ˯	���ښ�/�o���N�S �}�:�