��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������f(�7�u3�Oq�yW�ul�e�8�Jy��Au�*$-�������Nƍ���'&+���b5�m��X��{\1L*�]�%)����R�����aW���k�)x�&J���X�r9�M/l����q�3Ƙ$F,�\�I���"�����>$�S�Z�d������7Y�QaD���0Tsn��|j0�m��B�t.Oc�Ie-���G_v�|�Rڡu�S�
��n蝴E�FP�1�%	ר�h�~�d&�0��5!��&� v��n$^�`#�?���Eo��%�c�y[����7
&U� �Y 6Þ���]_���5Nv%���"I��ͥ;�Yl��a���Щʷ]D`���x��<�j���
q��LP��$�v�)�*U�\�R7i��	�ـRB��r�F�.���1�#���ٶ��^����΁����D�Ř���nK0�>��,�X�ۦ(E\U��Hdld�P����c�\pY�p��Α����M=���A0Ϫ��C6)�5��x����h���官�D̞��0 �SGUs��∬*�� ����K���*�������]���sw@c(�������:������n[w�ɵ��ݭ��r����rPx�!�d����P�}l���Y�# V�^������-�+����S�>B��������)�~��v���8�t ����~��F��@��W��ͬ�r0v�R�1d������J�B�!|�g��t~�a�5��d+	��Պ�D���xZ'uh����K��E�JmО�v�3K6�������X�Wr�X^A���x��H'����Æp[�LlD��Fq|F�\!¢y�#Yd���w,��~��
��SRpL��u�YWd4�vOs�,�э���2�����M�#\�鎟j�7ki�W����#��Y�MJ�os\+m�4�B#�����+���p$یq�*��|�B 
i�e;Ia5���p������2�.�ގ̮+Q�btR}��G�(4�{6��)�w?�o��I�h�$@@u���#�FO�s�jڋEc�)@�I�Z�}�!1��-6�ZF��W��v���01{��X� ^I�GMLg�\�#�V�<s�|�ݠk�(�h��Q�<���&����e�����yn��'V���� .�R�����sZ�rL#fT	������X+��40"�"w&hT�-��,^��&���fj�t�����[v��TM=.MԚ���-"c(�c��C�d�wYnse�d�&v'�Lj�z%���q֩?�\hT����`�����Gb� T�s�j�pP:�TJqؒaZ��(���Y�-�D}��$9Ϸ�l��p��'�5F�H
��QO����P6�'(k(�s]��y�Q4���;F(� �2i������.�bᢲj�2"Y�xq�ʘ�e��RdT�������+�WƗ1�6�5�-����pKۑ,�z7tbd�(9%u���s�Y����G�Poć�!�1�0��L��{]G^��SH�>B������iA���޲k��*���������*'�����Ǌdu�TC"�&���/��B�C��J �鰕I �\�gn��m6��+>���l�B�1���{l��ٱyԷ뮢�ƫ��]�<IL�U1���z��nX&e�D �L���{d Z�}*�����e��
r9X+�!Ϙ~Ƈ��73���C�l	�T�	��ƀ��Y���tg�Oq� �m��6���p��(���;����j `��@�[���!���P0��);m�J8'�A�:��Ibs5"�������h��^���*����d75���G��J��Ä�B���f˪6fc����L����&qm���<�%4����Ҟ �&S�2=L������1�!�#$iKXI1��"����U}�ﯨ,�o�!Q*��O�\���=���:�ԆM���{�)F�ĲһO����⒰R�I��uk�I�A�l�-e(�;D���|r�g�8W,���w���� *��fKG���%11���cc�����0X\KI ���no�)S��W+d�{����$w�g �#��_�m�+	)M>�3�(�#�۔�0d7��3o�PF��sf��z�\�wM}D����n��0 dAg]g���|o��'��0L>���Ŝ0���T]2|�gm�Ǩ!���YK[�N��n������<��$��m�|o��N�p]�;RUFD-�_���/2�	��<�e弊�a�`D�Ț�5m�t�GJ��|���ɻ�8h!�0�������a��V"4F,�
���ʩä#�ȷ5�gy�'+�{V�4�D�'�����F�o�+ز�%���ܴ��!a�6��\ee}A�E%ѳ���l6.��
��+���w���R���R�Vh�u�$�����^6 )]-�>�H��J�ݗ��p�F�������k�B�0]����4u0�R�R�+�MSR�1r�;�]�_�H�4��
�f3�	��a	�"�#Q�%�W�Ha�*�M0�����3Q�XG����Ζ��/|��x�ӔK+�`]��@��q�J�C���߲��3�>�}d���#��޽�"��؏I)����,�x�|��=S���oo��k��5�5{�"X'���\5|�]��R���Z�%��2(e����_5�e{%�T�M�8�gyp�1���+^ݟ�}����5�꧀�g_c�6�U �a/E�)�qg��U�V�|�&S�2+5lPQ��"��D���ܨ}�lA��	��4˵�o��f�	e_oy�����������X��Е͋�q���g�yCȀw���Lg���2�M�.Y��©*ϒ��P��\5��6<Y�8hg�B��[��/]���^PZW�A7"\;��ҷ�HEs�ٹ�Ň<�q�C��W�u��Ռ*��{��u�)��|�#��t��i�����i(�����!i�A�7+)I��9\��=E�|����l-�C������"p� �nRy1�z#���*�tI0��C�j�Ɲ�\�2��II����{�$�x}Ѻ���L��N�IhN:����bDL_sTo:��%��r�.N9�຃*$�I��+D�5\��E!c�y���EW�����0.@&�?� �Tz�&e�s���'Y���_#���hE��(Z���O��'o2[a�}Qi����� !�PW���f��0��V>(�b��6c*c�g*�RD�56Sơ߰�D;���dcc{&�ɧ��k�w��r�ӕ�^Q��ӷF9B�̿��ߠǃ��:N��-G��������&!��X$�*�2:k$��!H{\����e�B)������]uƐ�5�W�¶wi��j,#�>�>f�˪���Jq�r^�_5�~R8�[�O�ɑ�J���Y�"=��#�
�,���'�Z�gja/.��߶�V�fS��*s��Tuge��T�Ǿw�Xy.���h�
[f���cz�e. �{͹����|�Z��x �Puh<y1����f1��ו�u��/*@Y�#�;�~?��x�GDA���9���uD�#Juj[�ND-��\mRFn4����2�#a<�%p�s�,c5�����X-vX��F���:�H�k�6��o�.Q�=
vB-��.����X�D�Bs~_�#�׬�17�w�C�:�5pں�����Y�ƍlz1 &�;~U��y�L�O�}�.F�фV1<��hۥ�IM3���[/4��^e�7G������� �����V�&���/�X���� 4a�)�p�XK�q��a�W�g�����q�^	����E�!Xeܰ�h����<`=��pʚn6��,�K|n)CHY|*���.�uʋ�
J�#4��^a��>�L��n.jπJ+�y�]	;����� �Վ:W�����_,�]��6��ɴ�m�uN����{J��%~���BaA��^��8��@�*�P�U�i�6���p�>.�	�_����f�P.?Um;���$�"7��(��])�3j��%ӷֱ�h58�RϔP+x_K�pM�L�n8��e֔�����o�r=
�z�L=-?���w��#Z[߃��9k�$O|g��0���" �6���Yq��k���ۮ��	fuƩ5��*����9r���1�*S��O���������Kx�ߴ]�܀�")�4��г�8U��K*��o��q�w9@9�b)��&�r՟"���J���3@�d��s Ɗ�ׅ�xE�Uܘ�o�D}��_����~��J@�y���u��3jYj��.P��iJ\�;���Πz�3�	�w�5�&|]m�<�
w�<��R��%*i����Z�H�у�YK��&C�o�	ʞմo�fӹ{�2*����LuV�?m-��[�.6�/��ӳ�S��r��V�]@J(H�$�#x�3j�;���"3��Ns�O�U��!��7�bQ'��_��ԗ���� ����T,|���ݩ])��#�Ix��׳�WAv��l`�<C��V�J�N��t?0c�̧.������p$kضx� j��D��򺱤��*0�H8�2d����Qx%ulA�Q\h�I|3���"ḙC��Ң��L�$у�Α�}ѓ��-�oTb�4�J�M�o�7Jh��"5jY(��o�����S>$]�%HA;��ѱl{�"����	�����������*w:�g&�3�Y�V�A��2жS��#�)�7�T"�m3��֟ȱ��S���A`0j�Za�͋�Gx���O>����0�CX�T�`�&ht�,�2x��K3��J���(�=}�ZG��Ł��5�X �g�o�0��.*���<� ��+�ƞ9���bM�������ha�E�6d���r�s/Eׂ�Iݾ�%�4�e(A�?�o�jS>��~H5~C�I`�89�EEڱ�j	3��n�B<�靂���
kB�i�b�oy]�
���la�.#�Z\rc�S�"6�K�zsY��ޭȳ��2�7g�N�d9���+]�9`{(�*�E�X�Ħ�
�2��W�.sIA�Ԟx�rtȁ+~j\��
�}'�~R�U��u�	�n�.@gb����~��QZD��F�N�p�+��}�m�qg�2�K	�2<�D�������Jb4����5R�o��6��WʩP0Eu�S�U��aeB��De���_������=�����X�M�`A"���.��U��.N�qGO7��Ԝ�5N2P@Rњ"*-w$��S5��? T�~�����zީxu�<Z��9i���}�|��Dk���š̚���)=���;�!�P�1}��������W�RǁG����x��G��+Ղv��K��z�5 ������������]?�5!u���'cǁ��9*��@�<�����w9ǵ^�@xmW��[qN�qq�N�A+X|��?���cwCE7=��f{�ү��h|�����wX ?g�Ǹ�z5��q�W�:�"��mCx1�d�M�0�_U�吩/�;MG }js;w'��8��Gq*�2zW1���4q�����Ɍnw�G�C��cU���`���̂r��=L	�P����Ə܎z���4�R�	?$.[M1��l}B;F�pk~^�B���=���p���ۡZ�9L�<ۍA� ���X���� #�̴_LY28s _V.�C����
ct�K����,�V�1�̲L�ڪݧX�Mo�%)�[q���I�I��:�P�ו��:gv��Cb-:�o���Knc��>XXa>��I�1>��*��9�r(7볤�(W���%?�Sa��ޖ� �f%��9�I���E��'4L�:Fr�8���"�z�a#�d��*�I�%�C���x�z�����ij�9�k8�qz�S�4K�0�/���g����_x� �AF������o�Ra.�F�����9b�1��=�c/+��r��,n�<(5�Y���6����F����B��[j��v�WQ����IDI�fv_9eGĺS��z�ݩ�͒��Lսb纆i�|���Je��b���n����R5�<�e�Ofn�~N�	�B'0���6BUOji0ۍ������P��+�WQrk*��Y����>���^�dkv8^��²�cN���ŭ�:���/@����']�3���uzF^��\����`qb
�d��RmWH�d-��>�^-IL��5C�R�00�XXH���{��^�d{!�)k`g�v�(5�ޢ!U�"c�3�T�@����i��wĩ�7���Me}�8e�=�*r���7�F,$��M��qA�=����������r�PK�q�s�V&~Z�j-�>N�>��k����>�&ܭ~b��'���t+�l�z��O��SV�|�}]T������}Ï�?3-O�S*jM
<�¯�
^{T�(z"��0�)1?�?_H⡋��c ��wO��"�u���>���yN��!��mi��~�ے�ß��� ԝ�\����(�{���	&	'�������F��CU%�ۤ�xgF��q4$����NV����q���t��$#,���u�i�����Nײ�.[v��t��6��uwuL���A��V�u�:g�n�i!���y:��+9��HF~7���L���|���Y ��v�	�n|۲��n +�' ��eQn\�Y)�[x�@-��HW���:�U}fʁUa�����#�ιD]-���$&��>�9l�F�n.�1�6�yr����㹽[���U���0�\p#E