��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U��w�|��l���&Ϗ\g��G���-�ta1� 3���w6���><���e[�XtXB2���ɼ�m�H܆)T\��u�;���V�EN�d�K��3�J�M�3|�Nq`���c��t���푠k�D��>�ʯ����cx>i}�6��0���q\+�� <�#�o#��R�t	D ��<��2Z�)xO�_��-2ӡ>uMľ��ѭ���dF�(_O��M�lӨ�a?����aB�`������WM��mV�|lȐ�Gs��+�����4�����qx(�%J~�x�3�ڐ�8��`��x�|�#���Q��_�a�I�p�	�ub؈�[���xcIA�~޴;4��m�.q}�w��)-v�4�-&�ZO^/����$�ɏ-�7>X���	ǅD�g�e���b��q�#��&&��iΊ�T����0m�:��Z��>�A��c��t0�T�y����)��durj�*:��$8u�EhMac��ۻ������٠�S�[�Y��ïs���@��w�������$@�����������~�]K�q��?d3Xzwq�>/AZ^��+3/ӓ���`��`��_�fiiE~,*���z�LE�@n&O�Z�;؞h�θYl_��+�.A�GH;'��a��@H��7V�iY~<��1H��%�U�Y�j7����p��[���s�~.]�#�f{1�;j�TF���q/w�$39@��`Φ�dA��#�H����x~:x���s+f�Nv�e���߆�������T�-�:��yn.��#zŞ�P�i���{a���nq�n8
9�/9�1�э,�u~N��wJx�0&L����T�L�y���~W���.x���q�ԟo~W��6Ӟ3�vx[<*�j�"�x�F�� 0�fY���̶+�5c�r8o�d'1~�G.���Xj�i�{|�kƲv��L.k�zG�:�����a�A��8�-��l�>8k�� .����(Z��m�y)���m)Ǜ����՘��巜
��~[�S���&L/��&���M?�/��'���!zN��/)x�'�A=���a^/��b�T��ͭ�@ �$u�H����;�4�j[#���1�j��e�T��&�3�BM*���oӽ�4!\l(��a�ʠVi�������$!N���Mt����mJI�ش�0l�E)��+�h�Y���E��g����zM��K'P��
,�]SR�����MX�D2�U�)�q�
I�Ҫ��4����������P7�Q�P���Ձ �Ǫ�ݝ*.	J�l.��\�iĤ�}��^����ۆ���\�|Ï�ܣz_\��7���Ĭt�수��ռf!5�pt����ty\��Q�A|�٢R[}y)ù�&[<���0!���	Dq�U�);P>�y�W�Q||c���(4��%5'�g�'���C,#��FK�30��l�a��+!u��-������6o�����%�?QD�?Ʋ�b�Ԙ�yAM��*��m�8uKjU�2�F{w&�+�Jޗ+TP\�d�h�C8��~�\9M�m�$�f]C��hW�H�U_2��Y��4-1QJ>.�qyPK������0oy7�d�׉C�-'aN��8�|J�i�ʲd��/g�7�0H��k;�L�BՉF�J��T8���Ŵeκu�&.�H~�E��<|/5����2+�x� �}+�i����v���u<����56��ټv�	�\vohg�G����S�rF���ʀ��D��'C�����qw�i+�#�P� �6-s��&��x��+�k��B�>с᳸������2�)C�Q��)��My�q#2_{y𮎆y��7`�n����&{�<�@���Т��z9]�64g�Ɖ���*�Ѥb�����\���EGҔ�u���N�x[���\yD
t�ksA�>;��?1���,j�=�Dk���w�~6���F�%��W�y��wY��#��q�w$V=���o�ߒ��ty��V��M��^�����~�SY���6Xk=���xg^z/-8�qQZ�AC%٬���M����^[]̲��,Fa�s�Sb��~v6HŜ��n����n���[�I�>�������g:�K���d���P��=+tmm!	�kSbe��O��|�͉���2�[w(h���1���N6B]c�Z��b�<x�`�1���Vn��ͣ���9j��4���ݴ~�o!E
4(��$y	๹uQL�53w*j3@�٘�}�,"���Q��aJ >C��.�6@齪�Q?xlO� ��M��L�
~0�!Ҹ<WS�7d���k���!�L�-��,�V.�j~-��q]�������y<�'"g�$���璉�ǃY�ltBJ���=����uh����xh"�y�˒����u �����@2G���/[ w�~u��W����T�ΡY>��8,WJ;F=��ZO+/��5B;3瑐���j�� ~;��䝎+|��e���
H_���u�9N�t���V����U��$m3������BHlFOO�>]�Q��L�1ۜC�c�K�����<:	Rׯyi^��7UE�ɵ�Nkj�m��Fe�;�P�N-����Lǒv��m&��_	/��k�b��H ��m��n��;���נ ��?������(BgЧ���c�o�����	��-�[ˮiL���}�'j,��r�]��'i�w[�lN�l�6G~��x�KO�sB�E!؁ɚ
2"���}�&�pzi�����=�xo5����7L!r-�I0���'� `�/�iV�<=����vs�5��e��3�!�6T�q{�������,�.�dH��ȇ���������Pg�A:F���ã �ˏ��_��z^8<�G_���r�|�%�����\�6S�DG$^#���}|��� �k5���x�Cj2Ւ,X�%���<�cIB�y��侁��LDca�{�N�"���.&"(Im�F1���1�Ӈ��_j�I�D�O�R3��4������3�R�����ȯA�0�b�\��Z�61��d-�ܿ!*�;�g�c��?y>Tx.����ѣ������X;�l����Y1���PA��.;%W��|Y�Es�o�ZN�]OJ�YK	��(���A.�3'��Χ���}��h�sy4 ����v�`Q[�|O�3�P����P����r�(	!pz�r��w��RxQ$�EfqH�!�)g�jV�k��:�j��8��=�5c��.wSjLY}F�Cw��.��Wd�O����z �:�]�fMR�q�����.�*_ ]��u½�� ���P��k��}$u&l��T�R,K��Z��ђ��a����*��|�Β��<N�|[�a$� N2$L�n]�;JhY��;�=yb��O>J�������!�[t*�i㊵�&U���r:�y�v�[@��0�S`3?g�&�F�KfIۆuV�g�����u׋�ʫ'����=�o���G3���z�(
����^
��{Y��M[����DWX��L%�$;�<��&OAyA	� ����I� �$�}<��g=
��	���qp(��$��b�
�����.����SZ�UJ�b�[ÅkV���Ő���XVf��tD���t!y�kËA���Eܺ�۰�\d^���td߉�%��Z�k���H�Fx0G����.�#�����HFd���������fL���W�`�M���GF ��E��R�)RM+�ju�g��V.���9o[1�j��|��}Qb�D��7�2�W��y\X�
�=����X��A�{���#h��i��V3N��$=K"{�� ����6V���֥$/���OĆ��"7�§�\�P}���KYs���|�Ӧ�J�C�)����0�$ɇ��~-ٿ����˭"���)<�RG�L�5F��7�@����MJq�9-�\3ͭ�i�nw�{���͏۴��������%���l��Cx}9*h�R)���p���KP��bZ�N$�5�3���w�m��P�B��M���'k��{��B��`V�*@���
I����!�~��Ǆ:�ߦx���P�ʑ�c����t��{��85��[�m��MZ���n�.�������>*����n����QS��Ͳ%IC�����tO�/nG)�(:)�Vl�M� r���&YwR���/��U�B��7P&�_r̔�G�S�,���O;
�^a����T� rl����Iq!���Ԃgu\�C����.E�+Q
s�E�lQ�z���СV�β�P�yL�|���Y�:�?��pA�ʸ)X7�$"�-	?��2��-[���
�oK����FP+�����;��~�>ܚ��ghs��XAY Ub�	�(4Ҕ9F{��G�x#����׍{|\w��S��+��f��~�c=[R�e�	�{{�d-��s�'o臂b
WP�'9}�� yL�<&^�� ?P�����q���!]l�Y�[�����ؒ<��c����u�z�o F�Lw����ŝ�~Cv�� ��K^��"B�!G�U��7qj����`�"&���"IPJmpԨrN(� �t@�Zo�(r�9��Z�K��U�BJc'1�<
/�~#�����Ī�
���ڼb3p���jw�s�b;�q�#���~��;��;e��ޞ�=݇,�WNJ���7�9�H���B�٤[R�����;���K׽�T�l�=�/���߆���o�I�Y�&�� �ܸ���"��E\�)d7s%,m�㩴��<>e��H��;!a��!����e�?\��#��nz<�{���PV�b��e����lOb@�xY�6��C�r �՞���#���GX��J����Ⱥ�
u��߀����'e�iL	�5|3��-@QjF���T}W���	Wa�H�z�0G�����.a��&��T=�Eٻ$8_��Zo	�Ū��b��ʻ�ܗH}aX$n�[)�>�d|u-R�s[o[��Ws+G��oz��6�!U�@�9��Ǟ2+������c���ob��
YЩi���F<�s�;.�<g���Z/�+����=���"h�`ԍ�oD�G)��O�e0�� ��������'Q��؁��e�M�K���/Lm�H�����Hdkɉ��������t����P�`��o��\аVȄ�|޷���3�����γѰR^CBr`f)�r��xwn-�>���1U��g�B��7��wO��
��r*����r�V���J���Rij+�m�����ߡ�dL���Xm4� �VB�#Lִb5��ds����W;���GF�)ݱ��"����J$/ޛ-�y�����]c�L�����̵��V�k�����:����kOQ�U�p_��+�M+��x�ݜ��f�����;>]�_��Ƞ��XY�=wVf	t�P� �'��\H���	ۡ�	�H���%�Y���uT)�S暠������)w><������2'�ʾ��-��`+Ju]�K��R<s�MlO{N
���D�_]Rx�=��G�}���%�'�vj5�:H#==̥�������D1�'�"PO�^�kҏ�D1�`59� 8"�h�"�������iG�5ѐ��E�s|*��gG-�+k�Bf{� ���ٷ��4������=����no���� >�i@�B3��%a���?EI� +v���
������I�'�2��ࠇP�cy$7UH5@�$��c�&�?TFn�J�OYE��ŷ�a�-��m����v;�����ܥU�`Cg���s��C{bPh�b�p{X� ���O8SU'�j1���������V��ʍ��V������n��/#ra��{�rܔ�dPz��ٶ�[�O���IcWz\C�L0 � ��P�/����F�g�`��ꀌaH ɕ�i&�	��MN����l Ȏ�W�W�Va�2p���P��8+�_�ˊëw�zj����[SvN@�./c��N�	�d����)�E)��V$x���a��S?��������d߄:�q��8��)%����'q�vR6��r;�K%�ٞv�eЂ�'qB(>W�\p�VÉ�|��6*=m���H��E�[C��c�\��9��2���{j����=;�;�����S��A�C:�R.��h�P���7�ǃ~�q�[�����/�ه�ՉDk��T
���"�4��b �Ƥ���o�ʏ�$ 4��� �/��"��_�XO�Z��̔�������c�rٛ=aN�����Ӡ[a��� �����
�YG�z;7?8}WS�gg����:�=�e�$�<����l��.���t�EB�\FRw>�uU�>5�{�`2��^k���d�v>m��k0��:YRl?֪���-�O!�!�b�]�%)Q���..�O)�m�j�N�}?�Aè�1}z��eV�B,�N���|3�c�_V�h4z�uu��Eb�#�6X��1+�F.{�E�z�wg�Y�l�')� �ȿ#�Dl���� 8 Y�D�y̙0h��p��@�z#��[��S�4F�"���a r���To�Z˓�:|��+`�� ?��?׍!�/�2����d��S0��pFM9W���XL���,�	4G6ׁtPd$fi����eLʛ� ��b|W�!�� ={;&b�~\Ǽa�4��O�3c�4�K��.��j�._���9�D-0	r�	���>u������YLN�B�xb���ßò,a�d0�A��ʸ�I����_��0��d��jq�m��*e�>�x���x��E ����[C#	zo�a�s�����tA<�	��<�A�I��ϏA���O˲���i�~Q��{�o!+��'�%�[��2��GbPm���Z�zs�[)|ƛ?vT*l����\�U�A(�(�^�u��;	3>�<Y족�{�!W��!������;�`\�����������N�S!���w��j�'�R��H�P�?I#Ӵ��.sw})[&]`�1.�l�X�~D��6�9��(�ݑ�u�܆/����fXu��"�6b|�w���!:���k��Z�U�Q% ���Wɽm=�d[f}y�1�CFmO�!����釽�
�_В��PS�U�D�\�.C4���N^l�"#��>��c�}�A��9y�9�A��[Y�I�Go�.SV��1���iެS��.P5�5'��d_�86���W�k�u�0MF�f�n�X�ޟQ�Dq#����2P��E�U�Eh�`!�P���e��B�Ti� 4?�7�D�V�zm\n��0[D �X搝;�k ��|n$�r&u�w��2N�P+)�����|�J��v�����!��20���(���qB�0�4���8�S��;�#��)t�C�u���K%];隬(�ƹ�ٰ�pS�~��1���L�.]��~H�֍���ݤV<�{���C��dܟ�*8qN7�4H7"���̈́W�L[�^����-=�$-4ˆ<j�ݢ�����ݞrY���q��,�V�v�{ؖ��
x�sR��Q9N�w2 D��1����q��.A4[����	�9����Ty�H�X������uM�?�F|(�ٽ��^���.6E�z����w�!=�-ƷE�?k�2�-.*;���l_��ۧ���X���/�@������	zI�y˕Qx\���`�~�w�j�il���VӪ�;^u	��[��ϛN'[��d�@���C�>�JSG�E�� �zK���<���/�r�ꄥ�
D���h
d=�zGn�$76l�S���ܝ!Y�T���1=��,�CmE�Ka0������۷�]��j�z�p!bQz�tK�7�_m���С��D��<E�	�� �x�=��E&�n7F��Ԧ�
qM�Sk�vn�R�1��?(Q��x^�u
�}�NG�%ǗF߫�2��Z��p;\��.�ӱx"��P6�Es*�!�%^7e������1�mZ��ׇ--�?�/�cM)h�Չ��G��В�ݝ����M�o����9��^�*�gΔ��J	��g�4��F�:p(��;�e��"f@(�B*h��@��s����\��pK0	t�+��o'�Z�˳m[Zˎkr���F ���ʖ���U}�K���w,�gh��W]<[>d
��|O?�����Z�A���3�������a�F.�������~=����UBu8ީ�&hԬ7��<�X#�vn�e(Q���_���kX1�~l�����E�I<���ƙq�߆����59,al�4䒴�[#�^.��R�% �:yؕ�< ��
��E�����=��6��љT���l)ӜF�4�8�s�5��3��N�ɋ��MX�g.�d(�w-L�V��_AIM9�9j�ڙ��)R �ѷ���$]�[��F���������/�*NH�����c��	o�Y�7i����=���0ު����D8�+�_�j"�[�Q��*�\���W�Γ���܋��y���\\F6=�B�Ģx�{s��LD	M�h�T����_g��Bf�Y�H�!�{������5��?�b�[�0Z`U�Z�ߎn�(�6��VZ��y����r��o���*����g���E4V;��N�(�����)�'Ƅ
t����1����C^�BYm�W0���u/���*a�p�%ď�_k��է�	@,r� W�4+�\W�׈,��>�zM!��K ��J+n�U���N< #U��\�*��%�tM^2*ͺ���-��P���	e A�����%'�o�=�����,ewlh;%��(�S��ᱝN���{쇑��	�z�[t�A�^+AAΦ������h��^��j�5��(�r�[��+��ה�3
ڨ�� �mĨ)#���)N�fag�i5��Ze�'x}̌��p;>YsM�ۿ�DJ,.�a��H��'Ԝ?�dxȒ�$g����3 ��ׅ������@��Be7R`� �?f��;�ܔ�eX+��tT尰ѝ��#�]�}R�_KChƾ�S�Z�av��V�,��I��d6(��'��ڰW���&�7����fО%�e������\�ؿx�&�\��)�� � �Q��2r����4��%MB�ut�Y
P9�����1*!�2�0t|ٛ@R��Yaڰ��;��9[�;� o��:�?�6}>q	��1����-�F��q�1)��Mi�%8�| �Ȍ�.N �[�h쌕�/�h5+@�o���+���lĐ����w��Y�ʺH����r��`���D�Y������Ne��C%>hF��	�6@knlkj,�&g&�D}x4SN�JSڧe���e���~�#Fn?���ڑ����
��Vd}��x�.+9)������q^�h*��Ɏt-G�Ƚe����Ι�Sɔ�N�z�UC�Cǃ�0�ʅ�un:Ύ/s���C q:��\{��{�f�����wϵ��O7�������w_P�D�;�g�g�@��5-8��2H	��Y���(v��=����u<������#H��{O�U����̇G�}���=A�����٣�ս��ҷ�qe�����LI�$?.�2������N/)��nn�.�E���Vg�tV��ݠ�dFed�O}fD� ��Q=R�S�G_A�����W�(���+�� �
�V��1��6D휲5�L>J9�����@��b��˼�z&�������-;� �H� H؛���'}�?�=D�-��3�>|��6�~��M(]���C�{󜵀�|��}�=;i���s��S�]�U�5��z�2���X�1�\њ*�@�h=�k���]]к!���x�٧l�)ɩ9_�yN�5W�h���0��"�!1W��;|�1�B����Fa9N��i6ht,Md��Eo3v�L�-Rb+l����RA�C�;c@*��a������#~�M��KtT(�s�U����q݌�q��+���\W�����q��������,�����0�f���H5��/m�4�s�۽��G�fpLd.���2�(S?��J�����bϬY�Y:��n���kH39�Ͱ��ؠ��L
.j�)k�+#c��9�8T�x��n���s`<����bxz9,C;b�W;��������Wo�p��s�?��,���CJN���ҧܴ3o*H �{k;��o�"5Ԩ-��~��4�	[����DV:B��W�w�s���i�ķ��:R2�� SmƟ��M��>��W���b�	��e�Y����{�:n&�e��G�8N
-\W7�>l�vi�b CZyDn�$�X�rw`�u�z��\��BR���v�8�<��.�;Y�0G3₿��� Cm$<#t���+�V��1^Cj��}�[۟�.�������#�u�ͷ�4������L�۷X`M���4m�p��o�5O�����UdE�o@|,X�g�Q��Kem�[F���*���,�6K���\�.00@ �&���2ج�=��
\�ʜ^���_{�+�[MH7Y-J�آk̋�yn9J��r`9�Ao���n�6�ƪ��X�n����!s�Q�Ǭ��5<@n����M a��4����n(��.�"ifd�I�!�?Z՚��*�ǥ�x�+���.�Qq
)?�4 ~ �燀�\E�N)Kz"� ��\�#׌����Z7컌��ּ0e�6?Y6"�Mɯ"��	
�dD�x��������9N�t��~Y'~@�0
��2��"�. �P�~��ܵ}�������K�)�i������+w8o�е!Ř�߳���� E��<���%)��_��Y�?�Ra0a��m���D]W���)C*�l'��Y��[Ƚi���m��x*-uV�W�Ai�h�|T^�]��,����Ql�lL��9V8�O���3�бl�r�x�jg�{s��Κ��k�4?�S��J8�����S�q:�Qoz�/�2���*��m:"���홢դ۬�S���HHrWՒ��:�@)� 	��sc%F��\��0�}!����I[�¼�K�a�k�t/?#��g�g��;j�
�1���2ac����j-��:YP����l9S�������gz�|J��dH̑M�Md����k�D�{�,�/TQ����Ώ��/�攧5�:�&e�<��>֢�Υ�U�->�-9wW��č=(i�U���͒!6@W.�ë�̨�ƈݼ�����7h�dն2o���<��J|���遰K;n))R-�D��Fs�E��Ww=���A�w>���b�hwo���� �?��9+�Vw=�#oZ����LM�|�V?�����J����K0K�N����=MBg�RRtq80�+EZ��U!��!.��8S�z�۴O�81���i��L��{p�ĒVA	b�ch�`1��h*�I]p }������cPtk����Jo�^7�P:s%��Q@���U��KӍX��iչjǫY��|R��jP��;£}f��3��w��u��,2�����?�ɕ��+S�#�N�2�t3��L =mWP{��������EZf�1t������҃�ۯN�,$��TL��a�FHg�~�.j-<y�Z���\��a�W�|I�E%�b��vm�n�;�q����\�����JN]l�Sc�ȁ]-�7rò��AR��1s��B�r�foσ̧��P���{���|�BS�\���i9���9t�ݿ�@H���XE���5\���N��(nI�,>���>��LZ����I�7�-F�ǽ���R��U#m+��P쓏�Y{�!|w��%_�(��1L��b���ػ����ʌ%����L�A�Wb9H�1:-C/���t�.nީUs��7�»A�� PM�Ja��@9�09yNpwZc&�y��;5Qg��(U�>�41%@�"�3 ��¤Đ���t�4��"w�PF+�eI ���O��h��

prM(�.�a�/��
r�%��Ni9�o��s��t�d@z:����扦C �?3c�K��hL���	�]���ְ�}f�2Pd��a��}o��a��p�g��1#��)��zK/.�I*��3�yH�M��J��F"�\��D��u�L�y`N/i��#�N�v�K;u|��Yn����٨��}S��1C�潞�f���J{���	���:u�����%QO1|�s�T�1���}�HFn�,B$��1�3�_�;�X�7��]�3��9z�ChA��n���:V���AI��l���$���ps �uIR@w�~�qy�崭�b�Nۺ��x�S��{l_]�]Jd�:K��<I|;��f�}Ҕ��p#z@�US�dsT�S�v����
/���#����7��N_�y��VO������BVtOM�|�u��[��f5���D_�,E�	����n]� ���gPA�σ$�>�*q��e�x��5�'ׄ���Z�٭��\�փg-�ဵ[SV�t��-l_Y�]��e����h³mMı3������`Y*��|i���'�� ���7q�x��tq�,g�>����;w�rOWҪUA��$�3,Y�[4R���뀔�S�g;���yò�W��K�1RU����l^��*
�Uqf�;��ô ��@�U{�j�����2m0A���$����yY}�:��Ф���u#�7��',`��?7B�z�:욣^���)���b.,�[��$��>���:�V��E�&S�;���xnWf��M�*G�f��ש�ˌ���1�<̻�|���U���z�R�۶�22}==�Z�+΋�������zsc<��X�/tj�7m��G!nh�Vנ �*�~7 C�� ,�>�r��+�Ł���Aީ����Y0�~A���P�|�4�0��l��z��'�X�����������E\��� H������]��T��Z�)�A���^6�r��U�=���"��4H�o������_I@jKJ]�������~�z��T0�H�w�8i|M�3�a!1��O`*�G�4<o����_˳��I9{���@H�z&y����
��C��i��#0h7jK��a�	:��"�"3ÿҩ���}oi��$�$��(%T~���/�� ��Y�6�=�8405ּ	���ma�⦺��/��~��a��(�:>���3%�_��zbS|1�7x���Qv$�*}��ٲ�p��,m�;3Ej����fw|
�����pF�xȥ;��j����-��3Z��Q�G`�PReWoe�����C�I���@s\�`����Mс�U6�A>nj�i�ҵ2x�^�Ku_���I�)�V8�#}a��x�;�+S�FN�й�<�gj�־��?܀	Q�'E4��ǟs��@�X����>}z+9
ގ�ZP��r���1�.��a1nZ	G�0���J�k�.���>O�0+���3 l�X&.�&8xW�qr�F��V�]۵ ��v�X��K�hs����ق�[�?��4��{����"Ru����/YZ�:���*�&�;��xǱ���8|�vx�����5v����N���I��r$��H~F��(���a�#��9Vڳ�D�{���⟡꟩�a�zL��ݏ��:�^���w�%y%� e�M�zߖv7���ݝ���%;�����N��ۅY��c3���}�N�3P��N.�hZ�{P��P��n�D!�6��
�Q<E8������B�(�XG�6��]�"��7��ݒ6�צFcr��6�LȮ,�V�N�qC��O�YKȥ#�"Zgcu`�<KE�y��s�S�����S�jߚ�%�'jҫt;0T��-�����Ł���}�'b�������ä!�XO�<٘�-�N�����ʔRyK�ʗ� ��6�%��Tta����"c�������,H�%���� �K��t<��l瀍��x�'Ď���jc�JK�y@�	[��PU4�5��kF�j�b$�X��ul �K�k��:�l�*��n���i�=�m3W��'f,|��>G���T��K�up���m�h��Q�����T���9�QOgH��6	�.��ھ-�x�]���}�E����,X.����C�y�ɡ��>ˬ/�^��a>,(}���*�z<��p���r眍�����
p�l�Ҝ���E��2����c�H��0��a���X��8��ML��`�r����usO(p�$���|�����F�10�0�z�v�����[{rD[�����Z7�Щ����MO��j��8��`FN��h��Ф	S7V�x
�'���^��Z��� ��黔i�*tu[y��O�p����|2��:���5}��j��0W�S�����G��:�mn���