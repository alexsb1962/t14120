��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L�����I&V~u~[rR�C�XT���o����۟�V/]�@�!ӁUټ��)����؊������I�Xa-�w�H}�T0�me��|_��������M��)��H�BK���G֓�r`6��Lg�6�ދ��׌�ŵ�G�0�2�!�J��c]Mw(�C�����Af=�Эh�c��I+ݎ���O�� ��^1��0s���=9�߸K�V}9��^��*!�S�����p�QtVx]�����S`�)|e�_R ���bd���_63Y��UgN��l��"l�����I�Gɏ0�4��<vT�5���m�༇�µ�U��H��z�4�n]����-R������ބ��I>��L�� 4):E���V!����Q##^W`(�
�P�CI[q���Y�ӕ��Cp�5뿳�p�3� �agD oa��EčgF:K�=/��R��MV�ٳ P�"�:����Zk�Y �{��W��ϗ��ݟ)m�F0�XFk5 ����V�ӹ���:>�H�A_!��K�� pxH���КϿ''���H���%��?H�} VL�Wj��	[��WUt��6(2�"��M�2��d�)��*>\o�䝮6g̍�u&���;AV�{joНgl�z�-{@��oߕ�����W�S���i�f��5+��l�u�Q�vdy�-u��D�d�~�W��QX,_�_�IZ��E�]���v,Ik�5R̅<	�{�B�v�ū݄8��Nf�x�L��_��amY�A�A"���g�.��0U�8W�Y5sgVu�e��s,�	Ә�׹�+�YŅԘ�v�N��&�%��a�v���5@x�=
s�V����e��}�������Y�7��5�N���sе�>�1mN,I;+ev%3UӻP�d�����Y+���d��/��:e���(X�Jܿć��zY�<0b<L�Je��u(�Q�A;q��7	�|�e�	{<a�Dߍ��M������5ؾ�v�7�te�~E��
t�'=^/i^����:F}�B��6<
�����,�O�%�5��x`��� (/�l�#�����OLdgH�At�e����y��nQ�we��C��I�vq�S���L�0��.���s��&�q/��՟O(�.���G��3 �� �ѦK<p����ݿ��6�E�z�g�	ASQ�#�����V�r�0��GQ	�P]Жy��EeHH�.�T{r�ɬiX��;�	e��)��rq�N�E�-cPA�P�"@�6hޚ��Ӹ�vW�jg��#� G�0n�������0�653uV���l{�MU5��8�O�A	�(�ZՏW)�%�r$"��)M���.���ơ���L��cQi,��r�R.�xVmj���Na}@�������w�E�h��8�/<�4���<9mء>��։�����&F&��:܊y�Kۢ��;���E�Zx��Y��!��9f�2&�濩,�Ձ�����
�$�Ezy>�]��}_�_�����c��ʝ��CqT��������3c�GE��[Qy�9Jڳ,5�i;nn��bH��q�E� �.[� ��-��5����U=�=CR�?��;����`�bo:���V�ώ��\A��t	#�>��>�o=��7���F�o���c?��Ro��Ob4L ȃdͦ�9t3)�I�BJ�0���7�IJ�gl6���F�$=�{�����R�����[�Cx�m"RoyWb'�ߪ4FjU{?1ȧc��j�'�e���aQX\A�Y����K�*���������])�%��[������"/�+C�x'�Y�A�b�O�z�VM��Dv�qx�-l��j��d��ӣ�D1˴#m�3�#�4����Ѱh��hQ�A�my��/��X��<�y���/�2s;���zT��q�K�2JH|���\�#�7IFۺȲ���	�~�-���aq)�܅��pÒ��n:M([#_��jC
�����`{�G��\��SڔI�j_�E����ʴ�tz>��--�Qw:E��IT{�B�����,2=MXm��y���p�:��T��8w:��+��5l.yQ�°/z�R �l6l"�i� ۩�۪a�U�+E^E�fP�T;a��K(־�C�������\-F�xF�J�As!���
&�]`��i}7���<�w*��u&O��N$~II�>ɜ8�L�ad�C�[�y���_L��1�g�,�iSH%|���)^�z�}|Q+I}�E�=�ᢷz��㽧M{+i��NM����Bh��H���ż��+��@��,���_��|�K�F�nIF
ZO�[�u`��r#*IZ(2)��
��KJ���y B����wOl �K�
��ԉp�)���3��9VC�Z�F1i�9��\z.��-�B�)����fk=���\�`���+��y?��߮�q����sE�6 ��7�s��}�Srn9*�~ɶ�$�/�:~��$I���6�&A��<��jB��K�y���D��O��y���ڢ���̔��.��Ee'�'A�V���W����boTK(�x�d$�BJٔG�@n5<s?y��s�2�A�
���R@��#�4�y��!?(�^��%���H��1��3�Ch�A��EF�}����Jښ9�1�'!��Xn�hA���~l��o ���&����ST?pr-94t�|�&9�Y��)]`l��"ᾫ[x�A�2=S�� ���l
`���Q�GE�N�`����(4�^�j�!�|�˼Y�a:L�,R/E�H';@Ϸ>	�=MN0p��*�L��2�o�f0��_Ƿ�J�u�6p)V��-/��sec�^�1�c��}b&1[��o�4�z�-�q�!}���(]_�)P����Z�Ֆ�@Zq/�QL	C(u�D	Z���'��ʉ��R�\W��>N��s�lX�<��4zԜz����)g�'�r��YU2U\Tem��e�U�I�v�]�*l}���f�4j�ت�Q,c�+�/3�O�1;?X�2p�bog�o0t��z��m�2��f����H�*�h�S�N~�I�Lo%�^���s��)<�3-��\-�21���J:}/�%�;�E��)d�_0 �a2���>�3�S��;1��.�W�v�ڭ�b�UN��{?�����|���R	�.ˊ.f���)�F�Zl���I<��}	���]V�ڤm���K���+l@-��*�t��ö�#k̼5��,.�S*�;�����El�È�d�oL��xh��ލ46^� �|)�[���Ԕ�p�z��zf�,}(�v~���W=^�j�T��S�mP�mbI=)ҳ�G��nRķ'�M�kX��<ovmg˲�sY.v9��TdZ4���$,�o�߂<4�������Ri��=�̷�)����!��w�G{59R���%��y�֬Z�