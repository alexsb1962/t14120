��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^(Q�`QԤ9��<8��IϾ�} ��P�,X%��d^|�������6��X���@N�ykl[!�IҌ�x�*_Y#Fx�[����Iu���?2�F�r������[���_��ͳ��Ϭ�#G�G%$v��]]�(��$�f���;��ǘ�xgT0���S��{�.�k�q���j7����dK,�ۭgѩ��t���h!��'�3�x8��Ϡ���j��N]��1]���Rt��<��ۯ�7&?$�0���d�L�T�?�M���F���.�W�EnV��0KF��3��ᆜ͠Ϛ:a{�6��/��Kkl��,�;%C�)�L�~
 #��X�ǧ'�0��q��`��L�L M��v���b�	��#M�
u�;�^QK��'�����}�/�@��Ś1�`�)�ƌ����t��a����Ʋظy�!ϑ�>��.�W�gIu�`��N)����e��1i �VQ���?��Dn٦�F�-�Վ �u<t�7��� �PlY;��°��l�����P�&��dw�Д���L�j�{5�*��~V�C�}5�
�tAv��)]o4��_R�T��?�˟1#�>e�ҝ�So�*4g��/�Ǵ�ͻJt�@������"}8Uc��9�-�Q����j_kb/�=��G�Yǵl\y4o^D�5d���h��M��2|���ܓ ��?�8���$Ǉ�K���Y�h"2�)]o7��v�`>/�q�'�ǻ�k;HAg%E�4G#��1�Z��Habf!Y�V�yʎ`�+��sy�M|<(�+g�.�"=`�&�Cٝw0�ao6L:wo9�F�du
w9������gْ��.��z��/J��$�1������k���Z�6�H�*���=�$�����ݷ�@Ϥ�rJ��[&�&ж����cd���bU�t�䢧�aizci聯(�w<������'1\%,?�a��:w��.�#��p{�����c��a|g�N�˂�>���}���б���~�{��2���%A������S��0�2m�_� ���9o�ޠq�<�����h~(Tw��wVŐ������/'�E��N��H�RW&%�����h;&K`���>щ�d=rK�J.�ꔈnm�l�b�� ���.^��#�~�I�=쏵&$1Q¬�V���i�ǿ����x����vB<�6|��0nI?��P�Je�g;*���igz+�G������x�$���{28�?(��4�Ǒ��fJ�&������^̠CQ��J�\�/tcC?�h#>��J����
�� \!��}�V���7����~0 �:'~:���]v2�����V�R��d�n$��ͻ~�����Ɛ^w��<�?q�Gqf��(OoM�65���_�]����&�� �Vi|�73;S8��ݜ��z�#c�n�cL��+�c~�a���`���R�X��Y�K��M�ߗ���$�TMGɎFL����*�U�S��OJ1�>m�	�Ý����g��fKb+Ѝ���V�Gk �����D�"�$����'%ΘR��؆ ����c�_�#��r�x�ȵ�M���S]*	����>�C3�������d����'�T��؀ �1�:ӻ�A�B{���/�U�������]L��pf}mmӍ`�#�>��O�M �$����U�=�kf���-.O_�h���2��H�']P���(��C'z=�i�|�3��$��ŧ�f�o��BB����Z�F=W��'��~b�z��2�����0�nX4\�x����<!<�, B�� �`A��](Ǻ�VڃPO�K���k�zDW.	b�Q4ڴ�m�N�G�8ѡF�%*]�	�ۨ��pC���~�=�������+�)3XR(Y+'�w-�B���&P4�[%]�����K���c;����~sZ��n��������}Ĥ'q�!A8@������X���HsUf�VP��4&�֚a}�t����Cԍ���Be:���f	3ßh��|S��ʘwvX�f��t�;�B�4�ˋL��z���L�˯��J��c�{b��6��o��=��2%�Y����mF�����LdF��e��F���6a�6͎����ᎈ;��	B��$�Sw�LW���S���mc,)O�{m'�01��W4E�|�7�e��c�4}ni
pw�aa���s�^{����z�9]x��>QF�l�"+SL�~���RO0�ks䕰�
u�6� �#y��=���bz���-o{1 
>f6�J�D��g�9��S_��^�\������$�jr��z�����#�i�^��U�ڻu�$d���$�����7S��S��ר9�a��]���ֵќ�LO���l2�>���L��b~�V9�w�|�W���; ����L0�ZT8X��L�ҳu�-{���6�qWD�R��pB�*���o��^iY�z��PG�}Y�+�X�>+���/YǺ+��ѽ�&���6j��!�3�?�m�1�U�'���-����ֿ�^}�ĉ��-S��0��-������m��)�AN{�,��	+%Ֆ��vKռ >�Y?�(>_ ����0̆\�dŰMsW�dw'�Ah�bqN|E��2f�ٮ���k����s�;Bt�3x<*=,���:9=��ni&9�z�; �����y� ;Տ���h�Q��5 V����$;�]�3����u(�/8��3���b��KX\�Wg�(;��Ϊ���^�;�l�2��_�k(XڵZ���c����C��?����g�p1��<���=�Z�`60��7�5I��M�Ka�$�
,`���ff��u[@��.�ON�5��9�s�ptC��8��iֈ���ܣ�nz�ο�%�ZS�Q�uC0n>��Z��B���y�U`�;�N$���t�h�&LE�i^�a�H��L+�I�������e�x�)u�寏�^ԥ���HT�t�o�K$!�
����pǧ�,�r���ڌ�T#�2��<��2z�}u=�|xZN9p���R�Edc��.ե�Ml����<�䧊ڝWT�������˄h�!f���M�&�d #x	A|�Ӧ�Y�� i���
�9s5�ʃ[�.�n�\ŕ�e��U��ym�!f�N�I�. ^N���uS���܈�2}6R[-=�n���v)�Q�X^��al�,��{N�{��jw�}��x���a���=�H&�ԩ �y\E"��,�����'ņ��3�Q�Ot�W~���! �=gz�TJ���p�\���q'���)����K@	{�ia8-2��뿈e�8s��y�z ;k]+=�FO�]v+Y�W�ձxl���+��X˰=��G�,�c��򻣕T�`��4��/ɜ�ș-K]%y��L�O���E&�����F�]��i��vk�9�Nهh__��j}��l�W�����Z��RQ/"�/`�q� �w}���g���̪})�a�X�)�[!�������o"��XN��`+���<��ꛥ^wm��a\���!!�
E��k@�F�Ȼ[�WP
�J%45U�;T�Z��k5$�'Y둒 ���	�iu@�n�{�]+�#C�-Z��Ey�V3� Pa|h�����y��껋ß�6�чv�N�K�=>7![
���4�,�1L��S�6�G�#S|�j�W|x�\�qy�^(��#&
8�vZ��Q�N�;��^�wY\�	)����	�s���^���J4@��5�bs �Z\�Pr�{L{�-��9@*���bp]C���+��zI���Q��=`�yΔ�W�E��H�:R`Z�R����{u��D�荇��q�@�?�t�xC7���W����:S�z��;Ř>�Gc  a������j{z�DdX��[�� ��Y�b~N���	FE�@�d/\[Bx}�EE�2�/KiM$��t=���x���݊�xw\z���ǝu\-��2a�M.n��DfMqGAM�Con��dT}!U�/���څ������z�yr��K�4C�y���q1�C檾�yǸ�r\�i��	lgJ~qښ.��Z6�Y�;�����Îr�P~����	k͟�O��36A'D���������-r�ei#���V�(��+���ws�1!����G�<�b!|�c���۴4chj��Jur�B4�����z�,���U�ㅳH
�'�p@��x�4	ǫ�NH��:�Jo7�B�}P����1���QI*�R�,��V�ώ|���;V��ױ�9����1�b �b��ۧf����@�}�8@;�s�n�Oƻ;����듽~�`���""��sV�%@w��!R��-�(O�=]��Ŏ(��er�=;�#�.��A�ʒ���Ҭ`�t ��yFu�o����l�H^���5z-�_�T%MM��xAE96�����0��o�/��x���T����eMmId$L�*K����������tii)y3����	�c���q14���O#�C�@B����e�q*7tmQ�L��S��Zy���ߨ�y˝H��CK�9���<����	E�[8=�7��&7��t]?W�<G�R*���i-]�:K�c����O�7u��t*Q��@�Բ�c�l��O����Ê���6� !������ߨ��A`"	��X���vDi�u<=�c��:�����]� �L��7�:�Z-���,J ��g�^���A��ק� W���S͝�H��l��/�������pw!��/G�/.B��i�������d��s����^DR󆮻����z�c�@ǣ�T�v�V��ve���*��������b�$��Ei��FycKxhKg/��8�XK��NV�7#������EH�ĢBSĎ����8N�UA*ǧ����p�­0�X�s��$��^M�Ę���k�?���S殘�T��}�$<���,i��h����5Q�8d:�U�R��: d��u2+%ꯦ3k����.��Y۩
��j�ц��"��� r	��6p�]x0�z�s�v����b��k��D�UȢ�{/��v+iO�$�}���=7�<	�2_d�KM�}��8F�?9�b���^��{�,iLK(%%:�f����n�b����ٹ&��
�Z��%���$��������mp5>����e�Oz��5��XZ�i�������{�i�`�Pr��cc�N} P2��FRg�c�n�u�,uG���`���y�:W���$,jܲƑM�T�a�e����?)��zpM�0�0ϟK�w;e�)��<��R��X��`Ji	�-�����z�/ƸUIy^n�]G��N�w�4���o>#'_!{2h��"c��J�^�^d��5�d~t�z�3�R���:������x��`��b�}<�3@w��FbXk���1oD��G5F��\��s>8�U5�UI��~���]M�[���7'5)�2P�g��[Y�T���S l�B�箴�`%��q��7�Yj�|Ԯ��]s�Ƣ�
+�ܔy`�[E��K3ν[���G�H/���v�n�wD5]z:� 9h;TY������%𽢲�2�MI��jd�9h�(�Gk*�!F������߆�ޱ��].B�J�5���ū󳘅�[��׎ߑ�2��+��˽D��9�!��V&��t�>"�4�x�\���\�P8�|C�V�$���:��+Lu���\Ǵas����⦣�)��9:'<~�h�)N�t�l �2(�;�����'$?�G�%�A ���g���Ü*����1�����B݇8�&;� u�8 ��6�w���;��Đ���u�&6&�Ǝ�\�YGFU�B*��q��kC�-fM��v��%��='�8S��O;/s���)��Q���`y�;ê�j��?��p��jL�w����imGf�������Ͼ��p�K�� k�Q�UH�C��<MŅL�9��v�C%gȲ��^�ImEu@�xRz{2�1�Q��$n��J�]#R!�>�k?�<����
WN��7�E߃QƋ��r�Q�F~����>�G�5��j��Ɉ4k�9��yӢ}�Cd����%��P�����/C�������6�Ǝ��+h�j/���)���uN����@3�ν�zE�Ae�V�f�?��
G�K��\9`�}!��pi�F(:�f��$P�8��\Ԯj���6�3!0�����8 ��S��ΌC \�E�[����;:�ad���f H�;�B�f�Z�n�c
���������.*㗾�Q�=�e���`QpH�Ǵx�)�Kf�"ƐV|gE�����g�'� |�4�)��W�̑��3& /:Ob<z.��:�#�w�'ϟM@�;)Z �=�jl!�6y���t4]]�E�T�^9W=bC�yEA��|q���a�H�"��}��x�9�I��:Flsǝ��i¨���%��9�8ı7\|(�Z�����XR����M���5;T�ulÐA���1!�pA��b�,��In2!�0Ivk�iH��8�I���>ͱ{΀�g5o�nχƯǧ�˷g�;{>�v���j��x�dM��m=q,=�p[�lO�b)Y��Q=Uf98m���_X����])��O���gDi���k{�7�}B,�H~,�bo"@��]/w"������ĭ���l ��E��Z�����m��N�����PecH��P-��<*UG�7���I�����i��K�k�L��4|sos�&0��FV��,��D��Y�_�-�o�Ȱ	��]���=�]��Xu^H����S�o��ŕ�P%l��Ė��W�K*T���MP��W�苻��>��������p���]2�GC��/�{���ˑQAx+}��j���Nl����C��F�᧨�/�ѷ{��rD ��m�.���uX����v'�AZ�O��W�5����ڕ6aq�Z���ާ����)]AK����S�d6�9¿�oH�CojQk>R{��Z�!œ$��Q�6��t�?6M;�s��'���T�&�X��ʝ��������;��]��G�+;�(�����VLҨ>�*�Q�:��W�n�6!Qqd���i�B�/��-T�5�Y�*f��_�oV�9�
��ߟ� $�(/��Z�E��`P#�5( �W�S���EB@-ڸC�6Gi�.Td9�ش���%�߯gߒGG�ӕps���VD����ad����O5�%�Wph]��}���.���!>Ed�_9�6�v���L)˘^����FX7$h�1���FD.|Y�X&��ҝ"�B�B|�|oK���W`������Mi�7 `s_�^�ON�-�8���K企T<E�û2�^�H��<2
�7��܄�HX�>�6�U�V����Ϸ��� YM�Q��!.��z�?n���jT�O����:Q@	�_��D���&-%V���!��eV��?*��2�o~x ukpPp��(�O�[�4��Y��x����A49RL�e�TM��r�$�i�ař]��&e�~�N>��V�|.��6�н�ݭ4��zY��h%I�1�/Q�(�v��-�Z>�V�dx�G&���蜷c�f]�Z��a]���.	�?	��O�<Ԝ6}y�J̄��ふk�^p��e"G���P���v�	���jK��@��>�@�hU*�����F�e����_I�:��:��9o���ґ���1��Za~���#�J� ߜnУFzӭ����vB��]Q��=t�b.G�o��K��au���h0�Xl �FO��]�N睆��������r�������$M?8�p��A�P3�;*N�kR�uiX��T�=Ƌ�r w�W��,�?�ro݉"x��è�Q��0߬�YV�3�*n�ĵ:-��uĜ��_U�I�>�u�Ĥ��q�Y�k%�8/�_��I��Fe�*柞ɔR��I���z �_�{Z��+�����Ӿ謺j������䨚Ec}hI�iƙj7{C<Þ�^�W���c0��y�Po ����g�+~4Kɏ�bm��r�![��*b�3}��1%j�a�[��`;��fQT��9����}� �_k�����~�c�B�l{��?�.G��(�Op쌛;W�>~)�C
�*��OI�fS���m�Ou\��Ć���0,l")�\��
Bt�Z�_���਒��W�����
��K1B�5˫e����-XOS�Wh��{�%�u��㵒��B�W�\�P<��w�Ox�4�z����?�Վ�F�F��K|��g�֩�̽�@�w#�I7�M_�Z��g���j]����z��Of��ٜ��>d���Ϥ>*(�`�z]�a6Z /��k�'QS;���(C��g�QM����!ogj;U- I_�C�e�C�o��,��#)��Xe�ٖSD Q�g���Q;����2���
�ҟ�bd=�ϛ`K뗘,��fN�����sOIn���u�+��É\��(�Q������	0�x�b!��0��,$ݲ�^l �<������S�v�k��e���,�7L�f��k~d/G#���zy@�5�`�{�ّ(2=�j!=/�v�Ϋ��G�Yv�^��|�C��OV�5��Ѓ"�	@/75���q�� c]��6sp��ۊ5���1���ic�b�y�1~�R���8y�G0�s,���O�G�5*����YK��r)�W��^��m�6ς]�9+HK���?¹���W��߀y #��փJ�H�W!��E/
XqBL����t�	n�����P��
d��J�sc:%z��g jm��D�z[(v���*�����r3��3�!���r4K�:`c�%E �@U� ����Gj�I:�aD�� �3j�N���uN�"Y*5����D��2�R�K��P=?ݏ���I��45ڿJ� �_�Q�|��W����4�U	޽JL�e���Ĥ�tynp�,�Z�@�8��d�qgX���������*�v�VNj�(���FJ���S>�
�0ɶ�%�@Fh�x5�~�ڑ�Ö_Э��L��9At´!C����2|��� �k�=��Q���!̽�y�k_v���;�Y~i�wa:`�Vl�鉵Q/l{G�X�fU6#���=��Y�Z�1s�+���m{L�q��zϣ���,���! l�HkI����{[6��<��ǡ�������p������ޜ/�9FI�TK'��ڱS<m������E�����,�Ie ����&��>�J(q㿱�(��X��_�ADXyW>��c=5���)�Pݻɖ�-L3�̪����Ǝ��e�+� �!l���kk �2� ��0�Zآ�x_,;-.��m�d[�X���9��8����n��6l�}�2�~9%G������S �X�;���J�������F��.M�������g�>J��i���� ��G�-�=�5����7sN�j����큁[�3��n����4i�T�I^n����/{���m��l�\�C`��k?&�7��,��_��:�k+"��!��e��:/��������d���m�_��g��>��.Fj_�A��������J�1�A`���Abj��ϓ��>{0�'��v�\(��L��0��
�3���BDg����&$!G��H�	���7�YU��'��ِ+��V��n{GzA��(��P�csE�7nYۆ��ge���sװb���m$�@�\��x�K�&&U�D��*��A�ܕ��z���#��,<_s��(�:���:�E� ��	��k�^�A�9�"���Kz��.�jdY4���v�c ��r��P7��$�|F�@�j�w����ˊ{|��f��٩��� �R.�1��ZQ^��>�$<���>MY쩡�H< ��Z?��t!_1������yI�d/���X�?p%������x�l3H�@S���w�,��"��V���/n��N_��,S���	�`�X�yJ���"�E�*��K7;^:RJ�jf[F��Ec�]��;��9�%b�Cib{�y���� ����A�Pz���b��B�i�o��z�+"Fi�MH$�&!^�ӿ!�5C�p�/�&�������K7�#�N��C�Ż�c��t ��"i���HQL�U��#T�2I�RhLj{dૈF�5�&;A,/"H��4j��$5���B�h�e����{��'/�F�f>܌=)�0����"�ڥ�Y퍻����4������1ʍ ��*B�C���@� ]��u���Hq��V�(�Ω�-yli��o4�����g7%�NǼ��)?T̳��z�_��}��C�y�wM�Ev}%#��/d�;��r��@�J���Uo���Z��ԏRt�Y	vy�~J�����db������b��@�m�U�ٰ�6�K=j��D�#�B�!O�Oa"f4b�,���i-��d���b{����u����$?96����	S�1�^		|���M`t���dsh�h�(I��ߘe�,z�ͦ�#�Fl��(��T�v�[��s_��G�n^���U���*0��/��|�:��ִHO�mm �e���ZL�0ƞ�P���!���K[2���8����������7i�ȣG�^L�nE�7jSӣ@$A
b�m'daJ;w�����g���7�i�~�A�쾀�Q)n�����5��S}`4ԃ_ib�l��9c�.dy�h�ٮ\�<Eu�0�����'��9�1�(��-�>ō)k�{u���^��9ˈ�t��i�a��^�L�T:3�:�'�]������8c��܎\eAY"p��ߗ�v�� [���-6��6	t��oN�@�^�R���~8�yVv�*d���֯�ڝ�@�!/~+<�.�%./����f�H�WN�H�U�f� :�k��ngćg�����'�Nc �h2�#@���U�Xa����,0ɸ���-��]ڳ6�q����l�柵ڷt���O(IO�a"��w�(qq=�ꨙ��z}�5E�7�-��'����f��@ip���0�RK�վ[?��B�1�2� w.=�BC��nK��t��(�e��ݕ��K�B��e:�y�I(��P>D�(���R䤻�x)l���to&ҧ.�%�Hp��uɏ�-��f���������`#����6 �M������P:X����g|�y��vOW>��0~�'���"Z�� �?��t�Z�o����1J�2��_s⁖��UP�c3�z,k���iN�s���@8�q7v̵�:���7b�	ӄ3x��L�TR���ș��.=��~�m火b�!hUj��A���<r�F]���up���MN����Xm�*��O����*�p�����aB!VƲ-r�%�g�LhjG�#2�n�^=�U���=ѡ�a��V��6��4;{
c�A���st	�=���ڞ�>�LK��	�����C0���h��3�[��@H�a��dB�Z���&�~�F�V^{�Ⱦ� ����N��?�r%�TFd��7o�����j�Ct>:+���|(�}*�ѷ�M&|ͫ�Z�:)����~�r <F"��K=0�׮^���hp,�_d�%�� B:�"���䬎<����@�+��Zfذ�{b�LNYV��upw���/	�?=l}\��ٟ �Z��|Yw�-tS`���A����B�l�Z��g�Q�m���;F 
��FU�~8,�ar�i0�W)Sv�-�g�a,:�X�o��]�!vT	jfl�
�6*�:����42ޞ��.��Z���c"���]D*��_��n�?�������i��8u�Q�K�=��*��۶Qy��{7ۿ��4��!�ټ�=#|��7���U�K�J>�ol�+g#��a���]t�- ��[�2� �h������ieFCkq�����gp����^B�M�����8L���M��W���	�@��L�5��si'��R񭤧K��)c�(ANRN�z��Q�c�M�Z�hv�V:��&J4��"g<I׭�}�!����t��$���ݻ�ae�E�k�"��e�n�ʴb	?�O٫����p�	����4�D�GR@}2�H�n�I�Fs2�+�#�2�Ee�d�3�U�[?���	�)c�4���xQ���&d�M��yz��;vev�=�(�[���9`��|y�����/F��Յ��WX��[�|�/R��k�A���쑭ϱm.��0�)�X&��_���o� �3=��>��Y�S�f�m��>���Pv��{ �	+̝��e`sk�H�V�vV[�\�'�plRSk�����#a�-]�ڞsh�j=���tQ���?�E��ު�7&�|/�$��
&��N��g!���8Q���U���n!��~%O���Ӝk��*"A���>dڷi�	��	��5�¸�;8�[5��sr��6a��������~���bP�N �<�u�F�����g9�DPզ٘�ÝY%A(�?I��>g�2 ��B�e�YyZx�~s0�e2u����3�x5�F�I��He@���z����F�_��]�#�u ��C0�
�t=�Rq낌)���-�l�{�.��"�����]
j��q���EB��M,�wO���Rm���R��V|�t&כ}�ֻf{3aM(1�*�k����WZ�%[e���j� )B�Hm��⡾R�	3Dì~����}�����O�`��x�N�܈����{ݞ��ۯ� ��0�ߓA�4p��X��qr��J�=x��̠-r_���,~��o	���-����U<�+���ݍE,�~-fu��["�7��T���pP���ygD-�d��o�y���0g��I�e�8_�؃���a�RA�Q�XP�x�$�x�;s}/u�/�����<	v�#|��<�{+�CF�>�1��䋝e�=���>262S\���?՜^��¤�� ����(G{TX.$]��0�1䧧�����L��N��$t���:�Aw���q�x��jb�J�-�(�%�����)�&wA�X&������&�Z'4�J����i�����@R�o�����	��a��D��`N���"�� :xd�8��q����i\��^�i�|�c9@�D�4w	A�O�o�bX[�&��?�,�+��uŷx��dg�v���da ��O&Y¬i�a�L�I��g;���_�D;N0\s?�A2�T��T!9(���k���7��%G$��I����Zj���R�>�����Ċ�# ��ݽ���p"'��%��ΌCJ���0ֲ��W�����XNw΃ � ��a�%�~�4�dC����d�U
w�]�o�̎�����C%���eʽ*��;�S�NQ��ڞ]�H.{��l�J1��~��uYz�;�I��=/�Efǅ��z�����V�`�j�r��q�u(C^>>�V
�)�[Up�p�w��W}ݕa��QS�0�d����m��� ��V���F#�1��|n�0%$r�Ш^�[��/��V�*F�x���c�k!����*���Ӹx�N��<�w�|�x�p���ohy]��t��J�'��(�_Z3�f>3�Z���RzZۈ7ڊ�!���@�'\��b�v���n��Ȧ��^S���$�m�"3'k���6��n��b���ͣo�x��*׍���]䁂^H�4�'k��@-&�l�kt�!��T)�/�:���ںf��r���Rd)���@��ɛEd�m%� ��,R�7PlA�7�Hu�z��Y��T�x��n��ҕc;U����u�8	G$qf$&�4��Q*t�s|������g��=�Fi�YL��f��<5=s��SP��9y��Ǧ�@���E�.#�Eg����=��{�3\�`ۢ�Z���=�g�kdi�����0��<��dq�z�^�F��s��`�nۭk@�n������`3��r6�[����K��Q(���)Ѝ�b�r��k�cEك�,aw����d �Č��ë�<u
,P�s�V��N�t�a���� ��ZguϠ[ ��t�{�ġ�d�l���ƚ��z�Y���/�JT+S5=*zK�����:ܳy�l,���>����� V��k���g��5��!�u���{�8=~��O]�u5������FS	��2I F��J6�PYpɉ��Zn�	�'���~6��_NGi'�bRnb�k�7\��2D-�u�ϐ�u��k�J��Hd����g��O䧹 [ʝ��(��:OY8"��4��? nA;��S�q��D�å���KJCzl��|�r�vu�MJ�X�g��a	"Br����(�ּ	�G]���R�71��a��P��Z"iS}��=�BV��Bf<����|�7���:�嵣L|B	�\0t�w����+qͦ ��Qߒ��\/�?о�h>zf�)��`��n���x������O1$:m��X�Gv���";����׊��͠�����ӄb�Т3�m=�-�\VM .<�U 쭚�)a�o	ͦ�hm�#v[d�G0wȸ~S�;��j����ȝ�":Ö�H*\�K�`H�,���Bs���<���-���D�������w���sQ�a��i���+��=�8+��޼�ob�����K.}]�O�&�0�\��x����"�yť�z��K��w㢣a	�n=G�a��.!��}e��u	�FY9�i��{��O�G9�θ^P-�� d_�}��EZ*�V�p�Y#�J�{���#7߱�����KWΝ�$����e8�I[7�Dϰ>aL9���EKb�X&oF�P�v��t(��/�i6
 d��;z�ˍNM ��gxF ���qS�f�y������;0�p�IrH��θ������~���ؾ\���W�v1#b��:�E�5���'��JT��I��!�	�-�p�N� fP��*M���x��H(�Y������!h��p����6o�0�9��n|�:j�)�4e@����#:�uW�#k��Ph�25���6>�4l~Y�y��`�V��|�ا�%+�����ژ/��0�b�b�i��UV�.k8!�苜�/L��������ƙ8y%f���?������u"��ʻ=Y
�\��T#D��P5����n85��D�����{0X�q��������ӃB��Ƕ��䈼���=n�X ��-���3��,~Z��.��'����E{c��������@
i�5[h����;�9�f�+�JN���2��N5�P��#ߊ���:o���C��~�$��#�I2e�s?�1A��0UK��}Z���dm��t����_�Ȓ?E��U(���D_�����R�}�XJd��m`-�d�UN��0��E��4�;���5Fg��U#����\���J�⋱��k����v�@���ߥ�_rzu��N�KxM>!Z�`���1[Ʉ�zKRB�}��,(&���� G=p��RÉ�,���+��$�`��wfg�ˣa���լ{G�=����%^sєܪ_��d��{�-�-:���a������ԓ�����io���:�-�-ӹ!=���p�ܐf���z��k�Zi��4�r�ء|pM`;���!�Z �Q|�I�2�Ƴ��<#ZH����Q��=VJG�$U�#��l呱\�\�����8)��a��	�9�F�&a��.;�q����<�E��nf����>�Xm�f��n�c��W����G���u�&2�t����_���'��'�6c*��i���a�67	fx��(�̅���9�J���0��t����)�w	��M���4�/9] 2%G�ʐ�@��v��WB�h�@!	n����Y�D��Kq�6���N��O���<�VB	��M��kQ�(��z����R�0́ ��c�ТA�c���,W �1����l�q
y��%��'
�j�'�s��s�d����WP�$
Wr��ro
�dhѢ���j3M7GԣP�}��?j�c>��H^��O�m�<D�G�j�h]���S���n�6�����$K�z��,@d���Z�O̙�����,�F�pvf�wW�ya���72+��,��rr��1؀�i�L���.�G/́�Z��:ҥ�VE�U�T�Sź�q�����p�k����� G��`g�j��k���)�X�8��?/��9�P�T �WuK��m[�?���V=H*'cjXv����{�2��f���$;�a���
��x���t;e����os���jm#�{�#��7����bB��ƺ7c��9д�([�IF�"0����I�`ΒC�#m���n˱/��J�3
ؙJ�ْ�U����(��kHQ�=Q8)�;�1`�~5~z���f��@�e�K��ȏU�����NdѦ�?8�k����e�ԯ
�^zt����/�)��Y�_꼠��u��N�w����K)Ck�w����o��\Fg!��yp��\(��t��;�*�݆���A�M�øT�i\��d����鯸�I��^�4��W�ppkG���F�f�#���.e[ߑ��[p����j���Qo��]��!Hkwײ�B��L�T3*���	�5���V��� C�����hJ)7�k�.��H:��ȎV~#�OI@�1H������/2��\x�1Q�FXw��'��Q����5[�gY���m��; ª�PuZ���W��3v�z"���,}��߾/�w������R�^jD� ������>5I�I�S@ŋM�����[�6���7eS��`�/J/cV/���Q��_ �����#q���, 
�O�5*�,`��(Hx4\�>$t/�K�nѶПwPI��+�E�x�J�kh���+���C�.�RP=}DP������0�d������*�t����l7����_!i�n��*a�Yg��2�񻲫u�c��)��XՐ�q�+�L����6�q����:��I�V�1�l�t�-T*Bcnoe�Γnv�WUW�����Қ��W�?Rz����s3�h�t�k���kyWl)t�)ף�f�-sn�B�?���� ���P,�K*��On� ����]�����|��mÞ?n�$=x���:;�������N�6��0l�����C��nHa-��͒�鈖)�ew����Y*`�$+�NL�^���GY�i�I���9��C�����[�U��{�ǚ�яxq\%>
j�~��nn�ȏ&���56���D�n���x�Trl�)�j!��-�G�E'e�T��$���<ݍ>>���,���3x"4��*�ޒh�cz�|�k/��ÿ�@,�����ds>��ᯱ��bC�e����ʂ@�
�k�e�*p���8��b�9[%馵[���J�&� \,�NI��n~�����p_�[p�i�3��Մ!�g����\Q�pTf҂K��	GW����zq��A!S�MSp�i/%��K╧cNu9̙�
fG��7�c��K*�'��h$�/=o����)Mm�h�r?ؐÞ�xCbe��a��m;yMv�P����/�}��l�.�(bh��P�F�W���R�?!
��O�����:a&�9���Ʋ�W�4�[oR����(�ߠ|qiڭ�qG���ȯ�^�8����:���x"-�UӶ�E�,���!�ǂi�%"����a���`2�֦v���{���*	U�,�$��a9gchau��[���|'�U �^#�H��L�4�+%�%H_P�$����yJp"��(�|��3W�
��aW��G@�3Ɓ+�]-ׄͣV_L~JX:����������<ܾ�7���|y~�5�F7�ǌ0�+�3/��F��+� ��0�)׃���Z	�:�yGV1����L�{V�z��,$�g�� �g�|����#�.�2��h�
�H�CP�&6� �s�,�_|����̤	rj�^#jm����K��Ǒ���۴�	o"�������sd��6�>[	4�uHHU{lMի�P�]�PG�Ɗ�V���XN�Aʐ��R�Maou�"�|�7b���ڌ�S����f-��F*�'������'T!�F<	#*�!��;�uҳ�w{�yJ��G�\�	��ݝ�o��1��`0���]�w
� 4B�IO���3W���R�(rG)EFE��Hm�@��y#��{*Tv�����-#߷WԢ	�L��b��X�*�"��7�`N:��Q��͞<j�z���3%���vx$���[����~���>���� <���Ƿ�vl�!�%���{�Y
�Z�U|9+m|�Y����W�R�x��!n��ܚF�
��.��$����+�/�'[��׾#M�r���+f%�>"x[�e�ؐ���	��\�#���<��L�	R��Ji�U;A'��_{�//�$��z��F��)���Iw�<�����W-�&�б*ܞ���t����l�`D�Ӈ 9�����q �v��bw����p��崮����<���pkX��p�����ƕ� �Ѻ�ݡP+n�9��4*��� SE���N����BV�J\��6ov�p��uxpQ*8Ț� ��+��樥~]n�k,�l��u^wQn��|"@eaɜ�|`��T�i����g�XT'�A3j����z�.����7�?��N0����Ȥّ�.���0�����޹� ƭϝ�����˫egT*茖m��=uf-���&j�?�7�MfV"0�HE;+m^\bP�װ�)6]��.��`�-����XjS���=�R�݊��� @�5�P"'R#�@]�,*���GRC���=z<��Կ���q�@>�o�c6��rU�^�� ���sm!T�@�^-8��_����y�;�ɗE�Q��`|8v�Q�-���;(�G&o��?��+D�l������zS�c�ߧ��3�4����9�_D�~��T�2����&���k4G.a�\I��w���3[��H��C��;�}�������N�}�Cz7��@_h�&+�_B�Ү��Eu�����Քp�W��h�͕��}#�����_��m�~*�%w1����_m�Mv>+)�H�dv�W�r�0��Zϑa���W�v��4D�O1ZՂ�k� �n�"�h3�-O��iK�\���6V//ot�F��}�H��HG#d��C$Tn���B�(���t��	>]�I���C�����KN���D1zm�@�H�d��:���1p�^��#���x��|�3@ܻ<�bN�!_E���"�ul��Ra�Τ��@C��i�7{u�F*ug6�[��(��P2,?�X�H��=B�s���i��*	�;�Nù�T���s#��X�!d�^��V|��o�@vz�x��N��q�� &B��t���r��
��� ��n��t��[��m�g�9!
's��+[����2�Oci�E���QZ���M���a%��;5�BFv�|$���-˧�k�~�Mmޥ�L#�����X�M��I�n=�O�t+/t$��]���%�s���ݱ`�p���Ɨ�������{�F��4���eZ�}�7W��H
qV5�	=+�۫TǊa�hJ��_j�D2M�;nm\�8b~�b����f�>s��m)~ȧ���N�6�U�oU'��|����{g�)wD�����Zl��Xe�j�����&�N�-�4vb�,D��Y���͖n��`��P������֐\�_fZGB<W:���2㪇p�*Ȩ����ɱP[���)"�9)?�r*$ZC�}��&}����8�B�w͹��?�Y�h�u���E�3�g7-'
�_Q�:Fetu|��*1H
DYD��/J�@��|j0��s�ͩ�䍓YA���~KU������o�<��JP�"tb\o˜�=}'IC��|� �.�е�	��}3�~�$rb���]��?��6����˘̎��T��3"8�s�xo�����ꉂ�8���ψܯ��R'��C
�7������ȸ`�����L���Pj�%�χH�̣Z�*e�ZđV����V�������J4�Mނvx �� ���^=��%}+���cF�����B����!���ߙ�ѱ~<���\g8��bQ=@��_��|��#? �Ϗ�W:�{�MRc�C���Ʌ�S��ͫ�����i�F�1���릵�x��5��U��P��{E�N���LA���ɦ����� �Tsĩq�E���a6�`#�;�C�� mQ��#E�W5�0��O�\	�)Ǩ�P����FP?������[�ކ31
C��9⸛gN��^���?�y�=t�>���۳C�U.����-��h��B5cmgbF�i"�^�n��8��|�E���:ͻ�����&Ow�/���R -=������^��K��\j����(A޿d�X�_�0�6^e��:��D|Iٛ31;�2�u�G�L/Z�NiZ@�XT��
��b�4���+t:����hLS�4y���v�$T��Mw��,G��,��l��t^g�S��Q��ˏ��:2K��4/�a�k}��p�Ud��Vj���Q`�1��~cjW���$骺`\&w���R��1m�ƻf��  �`�m2�9����`�(Vj(�tڭ1u����J��!-�A�t;a嗟�����1&u�`A~����6M^�6�d���,wj`K�]����
�8y=A��#��S�S�qFV�kSٍwM|C��k�
��\���+5�u�n�ҫ_qO�Eu�U2���dWx�kb��a��	�"s%1���>㶥�I���S�ٮAC0=	�>�2�A��ߤ���U����8v��'"��@	����?*Ҩ��� TTg�]�#;�wT!����,�t�hz8H�%�E_\����_UDU�85���}\��,N�k0�P<�oJ�>1�}D��|���Wwg��o�������Ӡ�.�M|I���1	�?AK,U�b�am�ډ�q;:��।\�[��MW������6�c�
���Ų��M��e�]�8d�|��B4�<cK1����fUᨓ6��$���o���q�a�48I���qbM�2�B�?�)I