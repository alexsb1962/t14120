��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������V�Ud2�	5�M�\RE�X9�wy��æ���<��tXW�St<h��V]����[����K�5���?h��д�W ��[�DZ� �Z7a���S	��\X[�S.0!�82ј�p�B!����m��P��z f�YW�I/�t���C�Bh�h���t��P��I:#tv��M)�"�#�O����)�M��T�Y0�g8�E ?ig5���"��j^�L�RP�I���H_N���*�*��'��9F�9�Ht���J"��NWZ\���aj�E��w ���϶:d�S�L'N ��d�)ڴ�v����lZ�Ue۞��(�mQ��V|Ճ<�\ ��`�ߢO\S��*��"�0��
����pz�7��k�1|���2Vkϫ�����N7���@ܷ�����?{���D.@!�Zu}�,�6i�kbM.�����S���9�5Z+7�0�[��`��3=�d+j������˅W��?B�\A��x�S`tk"��3���k����Pz�ۀz9s
�C�.$��ձ8��6�X4�$����,ϲː��K�yG�!��>�`.��W��7EQ�jY��ep�@0GZCkf�w�Twy�燰:���8�2���lxI����=� �hT�.�A3�
�9�t<���O�h��L�w.�0�h��?/���R�N�Xd���K�δ��h����c/���fosu04&U�0�:C��\z#�y2�&���O����LZ�?C_���L(�r�#R��h&��U�\e�C=G*��9rO�z�.aDrDW��_�><�V�-n�S���V{�9Z��<��`
�2��KF
x��Ҁ�nܧr'��u�'[�	�49�Y�����[�����(��	�ř{Z�=���.��t;A��P�phw��X��Ԟ��k�9C���%~�p#�G���I�(EK_��ё4����-�E��m���X��eQK�ڷV"����T%)@,d�fo�����i���q�+;���@����+�iJ���]<�R>��=�ZͮF������!g��M@�t!�X3� 7�ቱ{�_h����M���/K��ȒA-s	|����� ���Ź��?� S���<4�$M�;vH��	��V���x�]����췫�W����
��>$V��&���i���q������Ηb��!!�[�ǿ���,š����G��1R���G<N�1{�<�Q#��N���\u)TЛ;�C/���c�ȝÿ�z���
C!1x]�Rˠ	�k(�(�\��}p�L�=���xLӊ&����e����8���
MK�x�=J����=&����b��	��o1�V���y�Ͻ��?�F�����H{���Y��TtcnP���v/���-W���FsRl8aǛ ��<��h�7i�Vm��o�5��3���l�H%<{D�i�UVz�ݟ���磋4�U�(����-A���������7)�t�%v�G=.����[��SBu���j��I 0dՂm�ƻ��P
�6�kň��f��o����Dȣ�n���mT����	Ym8���>�CKIGL�b�Y����S�&9גβ ��4P1.p�W'D�M��.���B���{�G؄�4n���(���nc7?KɽU1Ґ��(�:X��.G8�r�޵�yÐD��uO��Fer�����'�5�-rXT3\�0i�TI#8ʐ8�"�K,=K2����=��31s��h3�̝*-�v��� �N��SW�X8�_�ǈ�ʼB`R�I�+w���Q���̐r�#yH�Hf8�w'��fu'���;�?���F�(!h��*�`[Njs!���I�Z^��:�DH��
��mctUވ�5���7_D�llYգ�>Ƀ`�e�\�`ГRz��wQ:ڜ`�J��U�AÝ��J�IV�6"��l"mܚ�D�v�n`S���/�ر�2;uG�L�4)<�}7t��5`X�a?\�|1��(�u��ԕ �n��@�Bɶn���:d�1�/�hM
��X����(�n9��b�6��j�����/�k�AC�w����v�����(�A��6���z廒�ۧ����N��h*;U�q�C���$�~}�p��ǣy��I��)U3�Ǫ�l-�;Z�Ij�9��t2�f��*4c�I��qSu>��"~ܸv���/���yU�B�Lg���^%y6�$�%2ȁ#���o�O#�p�*�dB�H�qP�N�8)�;k�g9=�XK�Q�bw���G���Ww�M������k�)�VW^��>�GZ��`�K*���%�E0HTO֍��+�
,�:z����lF,�9�x�5��V�gz����i=]�d��P�>�",_/=uOB�5s�j��.v~����3.�p�F��r��չ�C׳�IgI�Ӏ5�\yr�H(����Զ��)46�K���;s*��`6q�:k;�:�Lۖ��)c��>ώ����WJ� �\�;9�8IB���Y~�:^�Z�N4�{��T�\e��j5��x�I��2�v�?�{��m@�����LӈTܼ[�����);d!n
.�E���0��\�׶�
�����!����S���_N�u��.��\ W����(�]-���X3F�KƋf�M�,/�|Y��DU�|���">̈���EׯQ�(�JAŤV�u�fv�-0�(��g�ɓh�K�X��	T�������aH������O\4�{�h�@�h���42n��F:b�\6>a�EFS3F|��f�3�	�Z$p�Q �	mKr��8%o�_"�#�7�3��yC���.�,_~w����H7î��ک�ĳ�0��{��J*��|@8)�Vg?� �\���]�\m�������RY����ϕ��n��r�U��H`x��<�;�#;ʦ��)�,&�Q��B�_��ݚ]�*UPq�R�n�c�0o�V64[i��6Ү;���eR��-�4���o���"M�Η�H�R��'O�7d�hiQ����ȢH&j)��,:+%�K-��,���	-A���)#>��ς�y;��7D�3di	��^��gg)оO�&!�v�ԛK��r`�����Zs>7��fۼ��J�^�8?���e�f��38�-q(�wzX����o�>$�A1�ɳP�Ҿ^xQ#}|6�]��9�{�N�zs{~Tb�Үw�|1:n�(6��l� e��c�ʑ�d�=䦢cp�zD�Ě"N P�sP�z�t�%m,�(va���ጚ����!����̟@Sx��OnW���X�H�*M���L�4����s�ҨuZ�=�y���c˞�T;J@��m�>9���|�@kE?41��E�G
^��r߲�2\,�q����(UB�q��Cr�<X<G�}7�f�FD��l�A�H���B��AG[Ü�/�(�2�F���dFZCyT�䅛t?��M���N��7�)C�?��E�@�&�e.�9)�wE���m�����U�a��`�����9aP_�ɛQׂܸX�H����s�w��9�����QWYU@�~����0j�u���_����O�*F���I�>����"?|��{�͕?���2C�� A#��5��D&"^ߩ���N�κ����-�_�=v�Ϥٰk>{���g�+TsAɂ�"jAƬ��8m���ޣ[�& �Y[Hv]ӛB R|}Z����@�tk@k�ǒu�khT�loc���*Si���;cf6N�7$�۵��ҳ9d4������RH%G�Q9���g�17̈U���ݦy�t%,5�g���J%�sոw�BUS��>�I��W��YdŞ�hΎm{�A�.3bƹ+7q���Qof��u��}6[����������Py$iA�@ɽ2�T����f���HC���� q�-WO:	�P95��y�/p��*QJ?��`Aܛ��d=��×Nq��8��h�a�c���X�;��[�dsa�I��4:�".�#�*�ܨ�ǁ���v#�{E�~Mg�F�P�u��C��<?c��� ,���1!M{��gD��CNPpA��B���FW�s+m���Z�S�B�Fx�4[��f��^=������A��ۜ�:�q%��v����x��0��-�p���L!Y��A��: ��3�74���L#��>�'-L�3w��^�2ؘZd�>��f�;���ND>iS�Ѽ/�]
s"���BDᐾ�Z	�1�@�R�8�<!O�^��%蛠ڜ�,��$�Cu����e�VSy�7�t�掜�'���.p[{�pUwR�W��9;��J�VgҠ��w�Ue�[����4����m�4�Ҷ��do��_9�4���a��&�����*<���o���یt_��	���ׂ�e�}��/�g�����'���A��-a�������t-e;۰*�7;�Bn�݆w�ǔ0�Q��2���TRZ�j�N�V�w6�;~�>t��#ط��HzJ�EpCu���L	���\o������e�5:��X�ٶ�P~!��~{�������/�H�z��b^��W����H�����rw� aJD�]+n<^�;Z��i5�����o�����˺�x�J��6�d?���B�îG��A��zt�}E-�ﮋB}/q�V[���«���BI��K�:��/�%��'�����PBG���횆B�v[�W_2;�����}��R%Y�W��}Xz�1���)���e��iK�� �%FD%(�,�M���HSq�Bd�b���u�|�����x;��O͏~R��8���i��Nq@C�
>0:����&��I�4��!ň�WVu�RXz�m�:�/�����AcQ������V� i�R:}��3���ŵY��Z�+g��Ê.h��o�b���I��F��h�%��+���JB+�j��'k܇�b=�������%���@$A�Dza�b͙���|��in��+o�mf�
n�3��DC1������X�7T��Č���7œD��CgX�:��>XQ�g��`��������Tz���D�W��m�V�Td��#C�4]��f�	�YnA�EI�u[A�`s@K�/`�{�[r��)!��D�t2D�͠�;��>H�HY��>grM=u+sZ_תĪZ]�-��f���-���:S?B��y��X5Q�Q����@Ow�����)��]~A��xp@����kp�� �a[����_�4�����4��.O,(%̰B%�0��`�3\�s/d��F�\&w���m�5��25�<N!�����/��S�@��"����my�y�<���2�4��:��c�t&	�Ȥ���`�X�a;[�8!@��`$�_"�z��ʛ����	�|�3'�5�"�<54j܁"��q�E��2Q
���}9�#j�ɷpƆ�H����|��MEs��+G�POo�)L�cZ�PD_���!��t�d���7o�G�h�K�Y{�|����HqԴ�ښ �;��ݸ ���(jw�J����!����H�6����3�Zo�������ש!~������D	S�����N���ݻ��L�z�[���M)]󕥈	�kZ���Gy3�+]W��Ai[?;[��0R�3�<��Q��۹)���kh&`m��p��y>X6r��L���/���,6W�W��fʖ��R�����<�0E*�A��\����Q[�1IR릁\��������l�F���ɩI��+"\B<x���+p�/EsBX���?HQ��Ժ,A������\
 �S�X�m
p�2c�`Ƴ���&�٬c���`�ik�y�)!�����}�&��X��V����J�BCZ�dx45�16.�Z�����ob�!YP��^U\��ݰU��>�&�/Q> у�Q��.��8�Юt:]xn[�u8��$i	&��Ē����}����O6c��U��ޛj ��bJ����u�NXuZ�L��d�5i3��6��{�w}��H�I�RNAYW�����<=�j���Ol����B>;LxV�8(�X`� ������η��@��l�˧<*
���p*�zYe�<��lRJ������k�uTf�������]�"���_9�:�fb����Ì���$�H9�y��G���,]b����ًK.�:ф%J]�K�Q'0�=��6���T��j��������_��i�"�tfu�������0q`��N}
��V��d� <b���� 8vg=���<��z�+��FE�'S鍶�}#���Pm������S����(������)2 �7�}О
~��rB���8A_�4=|3n�z�*gXUW�A�T���c�{Q�r�{�����UeEq����|�TQ e��6r�4�۶�@&��/1����v�>�|�q����I(y_�:�Plf2M�*,���)��)&�e]�K�&w�����dw�����!#'b�,&,��ݚ�k�W�
�퐴_Ғ�ec�3%=��(uz���aU�M�T~ECȃy>0Y8���9>�wSO�-[� ����]�� ���i�	��i�җF<����]Z�h䴗�h��gQ*�`��JX�/^���J( �� s�0�7��]��� M�����ƕ�F���R*1�L�ֺ���9�t#����k�S+"r��$m��G(nsQ�A-F�t�'�o"������C8Ջ�X�j�	�W�㘂�؋`������U�����
͕�G��=��	�Ff'�K8W�u�R�|������C}�;@�b���k����I�?���uR��</�N�E��ݳ��V�������͢�uYb��z�my�o|:�/ǆ���(�����@�H��\^�T��i�=��@R����Jps�b�8Do������b�}�|]+rd(t��s9��B�V`C����C�w�#.�=Ѹ�g���&�Y$�_s��5�"�A���(�Z�w�Q���R�����+sSL���dxWw������C8�H5�ٿ@܋c�-��jt�ߜS��t.!n�Q�Q�o�W�ϔ�Q��G��d�-�)kv��^NЭ�DG���G�$�ϱ����p甗xQ�4��!&��HhMR�W���*<}ߗd\$HS�?F�5�C0_��(؅��L'��3eZ���v�3�����07g�f�1����P*��&��d�r*�pы��M����MY\�)y��ڌ��U���M���.�����8�����#C=d�=�k�?���T�����8�N�"��%z�恇$��x�N�u���<e���jV��<q[�,~����8�_�$wl%�2�HM@���6�Ԧ9p۪p:�2|�c)�6%����g��m4�W:<�Qu�n�[y�3<d���{���� ����t���r���s.9IԹ<�!9{t�x:oz_KW��Ȳ���AǗ���+5��1%�?a�[��kz<w��h{%���F�$fx{��ܥEȎ=�a-�U)b�WG�!�6[2:���`Ӫ�wG����W�+@�{���^�-�α�<� 06��Hqܲ�Jn>��"��`�R �����'k&�O1�v�C��[�ۧ���Uʼ���.G��A(T�9=��	�=sj��%<�#Yx����"�����&�]�F'V��n%PA��r��S�D2��\u���3'�;�&�H@�
g)�?p�d��/�?�@�Gs|O��D%�+֚4���(i2�}�n�"�)�-ЄP�L��0G���N��Z-Z�퓗��p��S�9Ӑ�R�w;�t���L�3r�J�)6�07'J<1���;��`g�a ʻg��س�Y�*����G�n79m4��E��}�S�
����oJ�e����[�9��sz���7�(��,�J��6���w��y"��ЫzMi ;YB�sv+88�9��>�p�a�l�g.c�5�^�oO���ʥV6����uW[��P�·福7��b��ܺqj|��H�l���sU�Nz�V�N��r���l�c+���;Q�ˬ���4�R���pR=8m��5D�U�5��������-Z@x@�9�;�>�\*N�`����O��P����	�%R��K��Y+��k�)��W0_ܕ��E���oJ��9���i�ξ�P�$2��H�U4ZJ��Viw�4�n4ļ�f�aZ�ʓ�b�����_3R���?��}��p�e�	�odt�����U�[3l@�m�灱�}��j�AToe#� T�`�X���}��)s	b��J�Qm���}�|�[�6��Վ#җ��:�u"��>�o�'9���?��~�?�n��1f8a�+����A�l��r,�?`aت�����[��;���PԒu�����f����"/����End�.��ѫ�kˮ��_=����fU+��HK�W�Oc�q_5�P;����P2������}�Tl��ν��J3dW��r�
�x�	�5.my`?���ľ�l���GHv���*x��ذoFj���lvM�I�[#$��&|!�5y_�.E`����6�Ys��F���D�Kp����3~�Q�Ϛ�?�XI�tTC���~����Y<1BG�L�$QR�N��E̗�a_��(�,*�	=Hӥ�o���=��	���xc��}��?Y,O- N�d��~�[-�0��ƶɒ7�qJ���p�=�u[ZQ<_xr�-��u�����Nل��~_A5�<15�\�[Ӑu�Ei��@k�h��{����\d�{��m����T����jPz�(�v�D�����` �"jPΟ+��5��U�[��Ryx9��!L��^!�.[?I���&�Z��_GغXW[��>�(���89@����I�T�^3�5�#�[��LӴ�c�b�b{�(}�	����p�)�� �p�S$C�}e��;�{�|[�f��,:O��
�,.��4h�;p��9":�i�í<:�1@�2S�[�P*�rӞ�������]!���F=4ا���y������ay�&�]�n8���:9QW���*�c4+�>R���ݰ�`�= ���2N	��P�1����	�Y j�gE�-�nQ �Ȁ ��
�j�zc�GNeF|G�`PnQ4b�-wn~��<!�C#0j���=��<0��:n{؈���Z�w^�߯?�p���7��M�ˤ���b /FH�}	b�$�*��˳YRݢE�n�8��ن&����E|Y�Sn�K޻w%�ç�P���C<E�+��Fͭ�;~,\4`M�r����_���&/%Ӄ�f��rVʂ/�l�/��D{��d�5� F���?�(W��V���0lw8vʄh��s�*���0�!��a�j��:�*�K!(�S��H� ���^++M}16��\��9�؃w�  sT70��N\��G���2	�ɐ{����@�\�YP�ZE��è�\!�=���B}[�Oբ�d3�����LƋAv<����4���[+�f�\}�r�q�{�6��Ҫj�w�@�/#<Sp��n��*�b示��~����'��#��K ��C�ڄ��m���_h�� ���:���D?�W�~__<� Ԑ�[��尝�
�}e������.��iR`Ɯ	`@GQ�7�q�8iEX�2�U[
ժy���=I�;Dp�aƷ�G-?w��,�Fۖ���6�o���2�w�����4s�7�ϲ�/:z����&x��F"WHj���Sd�`#���p�?������ ��6��;#���Dn8@�嫮��B�~��h��r�����V�_nL�Y����P"Y*;6ŷ)@Ů|�C+A=[�����o��`5�@�>%���1���)�w�%��|�=T�m���e�|D���.���T�qߵ�G��8[3�4D_)D+�����ɃΦ�)
��.�ɯpq�\I�rn�I���U�����%2K3�ȷ�;Q=�gY:�U���\7��`��c�e'�j���sTU�@�c�r��܌f�l�V���v8�v�P$���ǮV���NhҮ`?bp,�����o>T��U�z�nq��)'��ʻ6�Fh�g)�� ��՜�x�s��/J+�U��� Y8j�*�A��E��7�Rϑ�ii��o�:��ƣw�b�jᛱ8z��~�Y/]-��(����n����"r&2n1o?F�S�b���c�e]�,��G��h(�qrٱf,����Ƥ!{��<�,=��Yq:�f��	z3�k����87NZ�����c%I��쟠���]��g�TS̡��9�7x~=(�6[&����w��w:� ���z����Ç|�)�+d�?�1ڪ�[�L-�v�J���qZ�x��]bH���e�'�M�K����La���_�v0Ժ�z��¡�:�X��vcc�;�x�X!;��� �溆�z��{r?�M�չm�v��Zd�A$d}+�-��h���@�7B��(��Mw��k7�ȋ�A2��VGf�Qc���^W�^���ҽ���R�G���]�L{��{Ȗ��W�]%���朐�ڒ� ?��_²��B��.ՎH꫔:9�]�f�1��^AǄ�`�����@p�D���ߦh�_�`jB�ar<-��z�M� ZD���$�,f\�C�b-���Z��#.���w�m��@�y&((!�rL���\'j{Jƕ�� ։\�s��1�ŶB�Htuhi�	�V������۔���؅�8���$ַ�g*!a�>�h5��+:.��8쏜]��zR��rD��e6��q�\�E�#pX��5����y�
�1�3Wo�N3�+�/��"Cy���L���R��ܺZ�>���r�nڔ���%d��7��/���1���Žd ߥ�edĳ�[55h���Њ1�������wXE��h �P5���f ;�wu��+y���.I���|^~c�{ Kz��v�*&��ck�%d�勌�}%���f�OV�'���J�!��a�ZmE�Y��I�i�*и5h�YV�+'.wFb�n8j�\?.�S�P����N��"y�k�5��Sv�k!KX0���U�?"�I�;���QW���z�ZR #\��5P(K�B�*����?��`��.-�w�ص�R��Ʀ=�h�\Lf@?�
Uzd�%���<��5~�Q�:#Pb���-zЊz�7 P�-��M�HF�X��-�V�*j��˧.�U[����+G�}�]��) ������M��΄GU{��S!Uh6_�$�T̎�[�MǡTL��eIaL	�=�V�!Yҵs�b���� ��L��z'�Z���fH�PS(����O *`{	�)��<3������p�zea/��Q��g��-�����`q%��CJ��Z.�ɗhB7r?�Aم��u�vF"��:��Mǐ��(�o��d�+,�E�8����GQ�BD��KiF��(t+k��IʳZ�Z����;NHIb�[e�P4
Y�����DZc�PZ"�ƐF{��C?�k��vBr��q�y�U�+1[4���9$;V��(/���Ͼ_������	!��&���'��lLM�'3F-���+��@��o��p���X��-ą̗`���#2���%�foh#'��)wq��0�=�v#�����=�dBG�"w>�Ɨ��f�5��]�I���F���nӪq�G��0�[!$�]��f�y���O36�P��8��!?=�I�-9kOH�6����dl��͓�
�����2��n�9�侽L�w.���q��$#)�>��X�"�!��z�Wqi�j$�ͅ�#Q2`�{>�b�������F�{Y����PA"��M��r�k��ֲ ����/��>!I�kzö]������6��s���;Ҝ�b��š���}�W�k�8l0�0��'�駄�])M�*�p]w�l�~����Ȗ�����Q"�*����o��[�^s����¤�	UFH�a"jC���2G)l� �-�?JX|�^J/(�}����*{������-z���=�ȕ����y���hh�
�u����xM)g8�|�;�s/;\�A��ąt��uuMb���|��J�Nh�i����4�j|-�q�?��Y:x=M89�6�eC
�z�%ύm��~�O�%bnИ�;A��U(��aC"���yvt��s����~�y�룖{r�̉휟"�x�h��!Ϧ�
|��7#��_��<4��v۝sP�B��?ՙ
P16���'*�@�p�}�l�ʌ��f|�@X-�چ#9xB��yT]��m����?�kǚx��nX	�+�X��Rprc��r6CnwNS���
�	���/BY���C����+=K�ѱ����n��H�C"�2�^>$*:�@Ǣ�ط|[�կQ��_d�;E�/D߸�Z��A�:HfU��W^ݟc�)�Aٺ�{|�_O�R��*ȭX�"��D�.�,.VV��m=�DvX|��(ux��ԧ)L[�|[��cW�IV�A��, ���̞4Lvu�~7&eV�����ШE��;
	��"R�(�;�������w\e�*�/<�
�ʗQ��8�,:��e�ca��p�{Z��6]���VR����"�JNl'���*���������E�ƭǗ|J�n��\��X"���U��@K�~��u��}����;�����]�A�S��$���M*���M���Co�����U�]��*���W��c�m�T�f�R3=e���)u1�5�N���y8X ��@�(�����c��߼b�����]q-j"�]�	�!s_��:��Lÿ׮�����oj���K���� �ģ��e>�I[�lV��h�+ M���}O��ߊc� v��.��%�.���r�0`���8)?[�g�KR��V�반��i�/�.�>��c�#��x��F�R?�9�f�f[�9�I-��äs�N�-ꪉH����S� Y+�����
�&�6��<p�9*xԵ]�O~)c��Qt�bt
hs��_��k�ld��WhC���O��Ǣ�I�Oo���2��h�����ɸ8[�G}��Sa	z[�U6��X��6-
�u��d�~�>��)1�����U��O�0��gR3��Q�;�/��ȥ����fa` ($]['�����-�8u��wy��Ď�S�7��y	�[Ou�wlr�_ZJ�����!�7.�bA�At<�[�/�
�{��Pyim���ð�a%u1�����D޼��Tu#Ur�~�r |�Yτ#�odN+��\a����ϐ�{����_��'���?�r�R*Z���f�i�S2c���ȟ������k��o�:��ry�5�D
�e�SSY������^TS�]F��&AQho�y�;�XL�E��q�9԰!�6�M��s��\���0�rI;N�F���h��K��O��܄�*j_��5H�e�^��*���.�%�(��Y��V��1>��صs�9�����Ny�J��a�k��ŧ_��.]��݁��tn��<:���Q��ӗ��$�����I�YI� ���4�`DW��t9 �)5�6o(�t�B�@���KJ�P�k�|@��M��:d�#�|t�9�3�� i�BΜ�> ����fװPD���|��ª�n�B*�ZZZ7�^{����ژ�HP��n���b����
��L9�#Ǟ�S�<0b><��T'a�O͊��s�cxY��0n���:��1�&�zV�$��>�)B�(CUq�*oOP���l}�䣪A,>�婡�5���kv
K�+d�Q�[ׅ��>N���p��s�ُ��U6�h���L���e���-����@a�!1k1z�[�]
h"��3�`��.��Z�Q)���e�0ػ�qC�!!P\��n�)ώc!$�r?bh]�b�Ԧz�4e��壝�MYX�_�a}.t�b��&ǖ�����e���_øG#c�n��@�ډT)���\xh�졸�֔�Ai��Hy*a/e������w�@8X������ܬ�%�w��F�O��xhX㸸Z�T�&�]h)A(�&C
���F�>qHg���A�mo��+˸�� ��Peޠ�kR�j7���hMl���m��z��f�­���u�`u�b�^
C�K|�o��=c�����>�l0ۘ��F�y�B��5���@7n�$ �z\ꨦΓ��B�?��LyEV挓��s�)5����*��A���]&N������� �챳��j>��!��H2���|V~�MI�,' ף&�+C(�5��avT ׇ��⍩er��Q���b~˟��)�������m��v!���Z��^oZ�:��!I�ͥ����D�A�"١)���|�l�%�o�����>���gm����A���^>��oIX�ٚ�
(WX���$x�s����;�y5��|��G�Ͽ�۴]-�����EJ�p(��n��B
k�-�o;I�G�H{k><ORT��߫b�v��0���� ����wy_�M��C7{��hp۰�u�����yu �Kuf�A��6Ε	��O��8K2���I,L꒎84憑��1b�Ra8	��Jt+���!c���~���f�}k�	]�{��0�����g��qK7�H��X:L�(�7�t�Y����zO)@���7G^ۊv"k��c�K�_?��%Ɓڱ #�g�|�0�(��H�qY�Qx�:��iL������	C8Xe�)����<��}a�RI�Q�ӛ� !��B8�B�?�ih�I�	&�m���T�i
�%l^�s�g��ج��]�o������$���L���f��c��$�^U61�6��Bls⫼��`��V��B ��N)+��̨��ט���r�s�d��	Ƣ[�=~
�?g�QN���ֿnf𞭛�d��fRK��ҷ�w�믱{A�j����~�ݠ��H�m�O ���ǻR����1�u�`��h(��7����HP������s�A�հRP�>�� +��l���e�fX
�,S��hPd�@�Yx�2��pT�=V�	r�ԅ�6�y 'c�<�� ;ң4Z�\��&�<�mq7t���/!Чby�		ƩUNB	�م�o�^�p#tK�q�W���s~�6�3E�s�� �v���[>�Y�F�tќs��r��
X,=Ea9F6|�}�ߣ��WB���,��l�m�+fSr�X�u0
�B������H�>@��ɫXMt� \c�d�R�IA<�V)uU��0�:������7<u����Θ��$n��S�l���غ���e�j�pv�7���'A\�kw�6s�i$(�֔�g[�\�x�7u������pZc)��>kY}���|I���S��d��Rp���l����+ɟ��A3mM� �8}���GWqc^D\�d<[j��� =�}<��\�d�"�[�%K��T~XK��`����v�6�j�e7���,/0ș��|. 5DnOW_w�[�x�jH0s�n��#�h�p���#j"����gV5y�(�4�u+��Y���!�c/��9y����Px��	�]�6����(��7<g�؀ѻ�
Z���Ye�3������h�Eh<����k;�Ѷ�E�S�j{��4Ǻü8D��.�u79��lD�L��[s�!-:���6�	>�\�A��J�g+U+;�� i�}n��Mv�U��kY����/x4L��h�A�b�6�ן�9t�.�^yx�����ǧϧڇ�3]
�H{i$�sYԀ���N�OD�Nb�L�ҤB�mo�Y�� �^f7�,ґ��I�5ޤ���Յۼ��M����]�#o\�5�-(s3���o9_
�T�*h=�;)���F�w�!���`���s֓��1��_��-7M�9yYʦ�'�S��^1o��Op��W�Eea�1�l
*���%W=!ҭ�Rիǵb�^�Y_.Od�����EQ��|��2��K2�NݶG��,К<п���{&&S���V��U��:Ԃ�u���I�\�ưcq��ڍ�R��I�D��mL,�B1��k[�V
-e/8�']��S��B�:i
�޻��ھ���@{]�	T$�	)�}���'`�D� ��ߍ�ƻK�yu
�z�#4��X��P�����>�֟�ҽ��f*�� �:1�t��?gC���%���G���
��^�����ɞr<��2֚�m�Z����5㚧 ��2���C�w��`�o�=�ԝ���DZ�GX�� �zoB�0��#=#.�����&���t]���ӈ�+�@6�*q��\�T�m�;���~�wS�c����͓~ m���2��ߛ��*�o��y�震w�t;�)�m�,����us�F$���}T�n�!ZQ� �\�P^Ii��>Z3�������8��G4�8�z�n�oʟJ��c�H��������]1���@Vˆ�P`���<�� )��O?C�a~����	�>w�cCMԷ:T��������"q�K/|�X�I��̓u����C''�+Z.{��̘izvj�~&�  �&Q�﮴�����5�gGM���j��$�K6+e�k�4
�j���(�ۗ�8�_�u���A�#8��/#����XN,��Kd~M�+5��-�ΆD��OA��?n���G��6�q�P�k� �@�2_�+⇌���Hjahc{��i�i�u,�`3rP�F�h�(�H0���ࣁ�6�-"�9�K�V�����t��݋��bE��N�`�x��I��T��S�)�	���^tg&��@�����4@y�����O\ �Ϩ�V^M�zЊ�w�?�|w���d�X��WU�-�l0���~_M�pH�.����R������w�S�����=3�T�i�3O�����@�F�x]�X���Ot?f����6z[��8o[A��G��iĘS�C��E�h����1$nݦϗ����k�x�D��,��W-M)4l���?��P�=^%^������}�n�e67��tC�>ǁ����7XﮀMN�����<Z�beL�A���`�D�@'�0-����Zc�{&��,J��R�W���)��V~�-Q�(A�؃=sͩ��t7�3I�e��,��bBX�S����t@���~�_~n�b�K��l�eT�ʗ�4&�����tZ8}�@ݧP ��xf"Z&�pu��N�E5�\t�웂i�	XKgi �OAL*�=��Ŀ�+�ݮ^iLeM_��P����E�ZZ
��o6(G��R��yn�) n���c`�s&�(���(�����_x+q���s*ͫ��NSB�N�Y2wy[V\�%Q��ײ
�z�e�B*���d	:�N>�S�0���^
¹q���Hݑ���(��o�N��_d],�=4_	o��7�8 �wJ�Q�D�ٝD�� �v�'�Z�f�\��Npt2�"#KB�d��J�!�"�`�tH�k,���5�7_�L�����G�0���BR�N����$.����Wd�	 {��Ęi�FɈQ����2ͅo$k��F�K�X�-�t��?Xg;r���@�WT-�R\	�}D�͌d4��j��DO���5����o����LK�ŝu�V�,3��5_N�$�����e��9՚F2�I~�'J�Q�0}�.+�^Q#��Za�cX�/5��X��Myt����X֭y �u�T<���� 4�0��W!���T���>(j�	�*�Xd'����v8�f �&�Ud�"U}�K/{8�����Q��O8����㲫�g�y�����>G2ӵ�KXG���H?���n�Zk!�
�)a��=����^�K�5}՛���MW{�.��v� v��u 7�%�[�t�_��pK,��⨏Ry�FI�S�$��&*m5��~�D樊e�^a%��&�K|0�>��SY�kXc����AjKIX�:w#-)�^���1�$J��ӚH����P�v9_zÝ�2;�)m��^��3��������wl
�._��G�����&;�7�P��f�Ŋw��C&�;{����B��1��8�v�d��<��|��p��Z��H�"܀�螩���ʲP�93?0|rUZBq��y�ߩ�2uz6H����gk��=t:}���q
N��n+M�q��[�|�N�����1z������;��A�e9;�����vH�ٽ���Qq��=6Q72:B��&��(������Q~*Ú-/�K����$�Oe�(��2}�M�U9��W���xؤ��^"�.�ph/��z$�k x�fOT��yP��H�v��SQs;Շ�f�'�WB v+�S�1����k��B�"���Ѧ#̲dt�O��R�l}c�m��,��[1�C6��!eE�ŸI`�ňI�{��B�F��3J��k?^VK���'ónV�X�ȶ������w
<��Q��R����ZSȧx���y��r&!�|gRQʥ0����0�m^UX��;x����>՜*5Ϡٿ�8<{������Y��623˗c_��Ѫ �M�ѡb�䊴��r��*��GV����In9�PZx�6!�GF��B��I���%�܆5�F���F�2��LNV0v�F�SG���pӂ�G�X�������p�"��~�HSW�y9/X��1�=�*�T�;u��Xh�k�oo�r/5�ܥK#�Xk����(�Br�1%V8��a]�u�Tj쎎L EJDzyO���u���m��N���h��̵@�;>ߎ�N3�62�I���.o�����%�	V�6��gJ����j�+�:�Ei>�����f�6�j�6{_���l�����"�s$JJ3�Y�v91!�(�oE��5�?$�ly���x������ЖV��XgT���7냞��}�/�\��n]p��/G�%'[2^evՏɀ^���a��NT�r����/��֗r�m�-��u�{�a" Ü/,2[���$+�Va^oP̿h�XՎ��,��$[�E��_��5��*7I6d����[Ԝ6���޲t�Q	�s(�7�*'�P~� N��6r���׸6��'���o�&��m�s��7���͝�X�W1M+{�z`��^��hU��߉���<�og"���XS���fCe���u'�:�ژ����ܯr���Ύ�u���
췿�݌�#�(n�e$=&n�v\��S����3j�V	N�'U�)�+zL3l>�G�+�e��w��/�5���v�G4���`��!��9��Ϡ����G������8y�9p���)���l��<���=��Ɓ��
�)��oI�&c)RaB⛴��l�t������_�,�v��Z��������g���q����h\����U9�*k�Z&I�Zp��h�hI��l��~�'��	k��i��s�_���W�.�����T���t�ږzLV�-+k ���XS�G��<�`Dc!x
����A)��a��E���jp"o�)	r9�7:�g�c��>���w��b�f�
$3ץ	�/����h�A(.�Sǹ���L�}D蜶@^3n~�&�0L[��e�l%��Bޑo�5hT)]�ZPKD*�Z�N+���e���`��QQ��y#|HN-�u~%��'���`e	ܮ	K4ݯf�UhMg�GD��w!Q��Us���X䧠�G��g����_M���^��D��9l퓑���`Ov���t����a�ؔx�2noY �~��`}>[�"�)e͂�}���ۉ
���d\u���O��	Յ�J~!�����ori�-H���zJ�o�^���_A �<z��I;#����kG76��(4C�Jp�.�)�x����a��s5P&q�m��LB�3����e�������l�� ИYf�eЛy��V��vK;3�c�\�)�%\jn7����ceL2uƤ�/�0���\{K�Jn�^; �&{n�r��I�\	�_'\x�H�Ě�VT
�
��1��Ft}�<aR�:�f⥐� �fh!��w��h��ڷ�U�+mx(��c-H%����C�l�^���5o���e@��몲4H �&tHB*@�Y":w���(]����S���I��_xM�8�?jó��¹J>����L �X����|K�ce kK��?( �˾�ar.���u�7ғ�b��;�����O�u��Z��<&[dި�~s��) ���2�VX�W�m9D���M�4�#A=��;��L7���Ce�Y�&�z��<�K��pՠ���)mHM�iX����%�5�D�����ڭ3U��
r��s^��s���_�=���M����{	��LsR�%v�8a�ޕ����P�ydF�� �:Ϯ� �Sk���0RCW@ے�\V�G���ھe�V׈!7���x�3u8�ن��XW�l����L �������k5�>���ur�{TtFbȈ=Q g��	ߧ��P}��T�U����h���@>��$��?�:�oLB�o��<#Y�os69�==^�<�Dr,	�Z]��qU�H�-�J	E��j���P6B�.{��+7���u�( qm�9vV"�#�?����ίz7"�|�M� !��)�F_����@�(ZR��^n �C��M�uA�Gsf
*�7a	c �u�������6�w����NX�pE�2���G��?)���q�Hg|�o��������F
t��/Fn��(�D�uVa���=+j~YøM�����5T��/�}��aj�=Fx�����]��d
Y؛����� R���8�m2�J�;�g-j���1�ѹ����TSLr$n�^_�0OJ�t\Q'�R���((p�+7~��CsI6}ʪؔ��EF��P"3"{�q�nx�I�������t^��=G����������<ޡ�(���������1k�P���LkJ�b�(ê&��+'��f]wV┊"b8bt;�2vd}�O2��q�;0���Ӂ�g�l�UU��u���
>7J��7&���l�[Ñz��em$�b�c;�e5���zd�mT}���ݰ����a�_5�.[���"�40�#�_���>�/ƯF��$�yf8:��s��GI�Z��9Y� ��7����x�{�q�k��ѡ�S�bMZ�عQ��yy��f��o�˥΄��ȣ�����YUz�l^�Q#�x��[��c�CЌ6���Ҧ��vX��ŀM=�\�V�{y���uJ��c�K��ne#�N��"��W���lB�,��AV����+�OB��6���ĪN�_��/�87�u��C ���ei�RpX���!JA��a�E_4�o��aFv`!lI]�b.�N�a�Uc[��KPۀ��P�x!�n8t`	�����U`�bR��q� ��;��	Χx�=�E�#�?��\��2t�#��_�uLy�8��vCE���K%@dPA� w�ό�k+�1|��;�-Z�9H�<n&Yw'�=/>ȹ��l�L���ǩ�K�J�0�S�t>dtz���5ّ�Iy�"�t�����2ad���u����o�n����g��/[Xc�"�O&�u><����j����*�����=����_��a�KHbu�TS�}�4����2=l�,�괬oð�
�^��Xi�~����e;���#�Α���j}��"�S�����<��va��EY �C�	Èٱ_FӦC��m�����V��A��6޵혖�MV͔�?WbfC����1�����A�Oa�>������������={�˂8��4z"֍��pxg�k>ZLT ������}���F����F�<��}���r�v����!��x�rw2��Ջ�:��݇�˃J�,C�{jp��2Uh�%-�D:܆N"�:b��3B&a������f�]n���f�$�P��ŇT�[Y��W�<�afnU�n)�����%����5�-���4I�S++�I�A�hŷ���r:�E4Bh�c�$�m�7�tAWCB1�j	�)�	(�����H�a�߷��������Q`���}}�˽yӉ��X��=��7 �9�ϥ2�ZB�[�	E�zň
���h�I$���E��F��p#n5]�� �Nv!ö���)m���1���]�{⯽i���T��5j�(�Qi���P�L�K�ap��?27�ʝ��C�L��ݫ�6e"��?5�Ј����Wo�q��W��O]|���pq��F��U�Kd-BďV�+���ץ�lKwxҹK{'C�������MO��sUa�@�&�D�h{c�Wk�	�����Y˸�@�izS�g���?�C��)�ur���,Mg��{20N?l�_�"�0�̴��2��l8<]y6
r��G�����RY1'7X9��$l����N���jpɆD������?�à}�'�� o��C��Z+z��kkE[��zp8]��@�dz{���^NFV��]�����M��E���F��{v��L����
��	v^�R8r�ֵ�+�־��Y��%pV�h�<��@i�E���_ ���kv|NL}�۶���(�v�M�s�?��x�{�Rf�;��.3���_�(�܄U}�2�+y0Qk�{fj�yz��%D��dsނ|���?�xKJ�裘ǲs��}�W�t�آ�A����FWh��雩��bm�����+Ƃ��@�VG���Gk�>;u�;~��ؑu�����t���W�ls�R�����򦔫hH��q��
:c�@�׼�Vv��䗒�=��5��3u�.���j�_�p����.G�9�P���ޫ;i.l��vo߲{���ڷgl;+�[���'�q��:���u��--�q��*t*t��f�-E`���	-:S����ތ��-N&�aA⨾���Z����4��7��~� O��CD
�U?~(��a�0i9�-���(�dB�]ϳ�����S��0��+&���J�9;+K��}9�|v��zr��٥�Z&`l	��^U1h^`S�ߟV̵N@_o��V�e�_���cT	�ݩ���G�0d+m���J��ڗ٘�p�w�~�+7js�=����L{�bXxEVS��ͱm�c��5��k��&<�c����7�W�E�u�Pw�m�D �'1���A���<���Y�����=�Ê��	�0o���[�)���x$�V�����C��/�-��-��ǟP!�zd4	��L5	�km����E�`e ���U��5H����Fn9�EXt�j����S
͛�e��GQ(>����^�Z�Lc��嗉�X ��f�#�˝�*@v����W������wKjx�ٴ�$�S��'���j*�3*�;�"L���n�yS�C�j�Qה���E�3�zYr��k��8�T��?M}G��D[��h�(H��I�|��T�)�l_@5�q��ׯ�n�ab`��ʡ��q���)(�5?"<x�44�aBʱ��ls���l�Z~-�4�Ɵ�u�wm5���9D�ɗ���,>���m�z�!V�840V0j}à.Z#���Q/��i��{�=��&o�:�/�*�/,�}��`������Uep�z,�.l"�C��p�U����n_���%��7N���1g�`�ֵ�&;ś�Yl��Q_ j5��/�ad�B���8�ã"�$H��6���I|�f
�=��t���.l.˱BU&��9������\3l)J���>ҡ�41rh J��s���T�4�:�R�b# w��J�`��;$oT��g�bT��`�uU�	N���Q,���ҚفAȈ�?�����3|/ڧ��	����ct���mt�}�Kg���������:l���k����C�\;��:Ǡ�Rc(S�,��q�Ժ���m��9�ŧ_~��0�s���PfX�G�:�A�EV���ϸ=g��bɰkh�s
�q�	��am����?4U�����䈝��	����3`�mϟ��>O|��)M���~�Yt��4m����)|>;N�{O2�`y@��r\�@(���X��$�Z��	����V{cI7�O,l���Y�:���٩����M9�,�	�d<��"�8އ�֐��^W��FqF��C7uI��t<IމA91�W��"R�<k<J|a閫�l�3na5*�7E��
���'��P���x���q	4�d��!�c�%̺��$�X�f��� ���N]�bBf�**	<����F�/�&e�Ƙ��m �;ͺ�9S�z���m-wua0;�8���y"A�z��f�~2ф������)����g�"(�z�-����2�aX�MP�=��^p���6��[��~���4Z=�w�����91�������\��s�y���G��� ��ۍ;J�l�o����ϝ��-���Q��f*b2��"ON�sO�>b�(D��#�z:�'}�Q�v�9����+�r� ���K�D˂��,�X���䣂4�Fp8b���)k���M����;xH+M/x�#��]���E��I��Xs>���=�t")F�
,W�(�n
�$��C���"�q�w�*�Z?�j�}9��9�0W�Z�(�o.�޳��b�Ui��*��T�`�뼠��2B�A����K6����h��$VD"[�G�l���XYv2�i�ɸ�켓��H��U�L��]K���Ɗv9���t1��_��o)��IcI�k�n����T�Ŋ���\mw�鋅)RmK��J�ūW�#@.�5ǉ�������1#\]{�
�R��a��v��'�GT%M`��#~e�5�mʍAt"�n��ѾV��#4�Q׼dG�d���QI��|	����:�YH�ph%��پ�a]�<o��!?��2�r
���tOe�Pm����7!I�;/c�$��I�9k�Zf����(���DI
ֵ��2����m��x0"�-8C��xp����Ǣ�h�<�<M� ��3���&��L�]ڒ��|��K���CU��������۟�b�v�Z̯���E]p�t�v�9�bu��Ѐn���UZ�q�(�Y�ǥ�]������e���7u�<+A{��)�,�/� 9�NRZ�45G�G�	�I�_!�i|i#�z��P�-��5n��f���l>�
B��;=c,�+��H�횧�?�z;�dar�MG�k�JP�fu�3�`*z�?V| �G�tl��<4�Ȁ�I�R�e���
x��I�P�P�?��+�y�%mp�N%	wwf�Ԓ�9j�3�q,�? �[��x�D��gb��i����b�-�ow#[�e�q�֮L�W3�����3�Ԃ���v����o�Ғ�1�R"�xſ�����^c||�'�`ռDt
L�Y�ϴ��	_5>)e��i4`���ME^b'nO@;.��Y��d}�m�:���k0ދ[	�9Zd�C���&l���vϖ��	7���k:��=^H4l4�rݙ���kl����2��3�z��9`�1~8����T1Gt�����d�K%9��c��T�DK��^��E�,�t�7Oo�^Ӯ�?����'��4�f�a/zntq��4X�%��sX��Rk'���Q�qz�Z�B�:Iײ��C.�lj׀p�[��H�l����n���>0.xe���ԗ#�������!=��/�E�f��?��}<=h~�jb��{�dZ'KL��4�~|�N7��0w�uI�YlP,�nh5�Ӓbvi��پ��`�������Uyq~�7��t�Ѽ�Vf2��������]��]δ�H���s��e��C��;�qg�XK隫p���@��kg�*�cU�f����ѣ�!b�Gu�QG`3�KgZ�z��k�jpk��i�JOUs���*B�$��R��͓�o�Er�@h'o)7?�-�&P�s�.m:��*�?Ks���X	Y�4-,vs���@���^���~D�I��ϛ��+w?A؞���H��/�lG<`>z�Q��D& g]��H��� p�����N��N�<��t�x�V�jB0U)�؎�q@�~#	��vof[��z��|�ko�r���*��<-
���#
���0F}o�����&%����"�g#�Q'������_��ea��}����Ky��z���
X����Q���Tv�bm�����b��b�
������6�$B�>�zk^��s�+7��� �
볒�BLڮP������'�*�g��1���w<�eѝ�N�V&�{2H�u�����`Viѵ1D3�ZNM���!cU�s��B��Y���xp�hQ���K��N�
O?F:榥h:,۱.�RU��t�p�ֆ�M�g�ՅCi6�d�#�ǎZ��q��/�ēb��������U�H���'B�weoo�K�&}�B�P�)�ƺёg%>�ՑĿ��o��~�-�#2k�X�A��"Ӹ:���8�$�t">���vgb#"�P��&�gj�����l�
q�jX8�%�4FYk��7's��{�>U2��꼿�[qy3H���Z�:��Q���2�
��W�|��}۝'��t��I<64�ba��q��ԡ���S�_k8K��A�&�6�#q����?8��[����b��mh�#B�\�YXtl�
���D�ِR�@�'�5V�vٵn��(�y,������9��0eX������B��ӧ�E��`�eQh��5�d���7�Y�;�#��Uc�N���k>5�z�x�7w!����8���&�S2Πh�m3q1��Ӵը�R��K��F]f��ҟ�B;��X�4����Z����y�0	�Y���)F���8�L�z�?8*����� ��nz���	F�W�oT�g����r��`�ܜ$��/d<�CW<����[��(�9�Դ�4�:���	�OW��qI�qv�t����������dĀl|���Nć:s��t��ڿ[e�PnY��~��8m�������n�!�8�bV}�J�"ON���4lA�Q�0��e��~-�&`����ރ����� �2Fߠ�z�<���c�B뙴�8�$Z���*ME7�>N�[������
��^�_Y�v.H�ןٗ5�`��$�/ē^1!v;)y,-�u$�QeK��sT��q���#@�_�ȕ��0|�hYY�����9��ܬb6x;���%Ɔ���������+�ߋ��u��`C};Žb���w�1DAX>�/rX�Iެ�g�#ST[o���y�����V?� {=W��ŕ(����h�2��ם��<�<���a�nJmY�tګm)��i�j�	�\^�㫀5\SO�Ef�R%2��\{��0�s�\��3i�7��3��B���$��پ��$���UKu���ܻ���c�oe�����J�ⰾ��	z֓'&�g$e&Q�H�(5���t{V�BR��8r�	ҵYT����˭�X���(���D次-	�K��wA�r-ѠԮrv���r��qzZm�#�^��~��pyJ�.B���g��"�a�t��*��֯��AY�ڨ�O���0u�S�v��&P�������H�d�����9��ZT��8��x�-���(wY9J�l7� �7����z�7�.o��)8��%(������(���iͬ��$��]���o��3�ß���ؙ�?aR�{v�j��"��A�����yv��De5��x����yF�$@8;��S2����VVv���$�!vy�N��IO \r��d�#��s ��z�2��"s�&,�kg�|]���ɐ���	�XdL@�>괻H ��V�To��<���{�t� L`{�M����$eR�_�م!b���:78X�K��Z�G��F��8�o�������fܦ�浘9po�J���cv�X9k
���)�ů�m���<��PX��� ��2��}��0��߭7�б�}���C��bnk<��oR��B��U���*IC��a���ܝr�(��)Yh=�C�Ul������y`n;X~mA�����:L�bRa��w��l>5��*[::L{�UX�G�(F�>�ꀇev��@=T�e|&;���St��/�0�7�