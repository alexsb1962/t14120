��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������f(�7�u3臉C�Ӧ&�$�O/{�)���i"#���7���3��,�D������ Q\@�n�f$4e���vwP�S�g��A�NK����~=�/v��	P�-�=ѹύʉ���=X�1Ѿ�o���os�(�B6�h�8�F�S*��^�ߓ�PL�w��:r�d�s��3��*��� �=�z����_�ڜOr�bp���e|7��\�Tc�=0*5�<����cWa�<AD�gC���	��{x��~C>RW�j�N�d�n�g�����%� p�Z��ARd�S���=V���ě��+��믪�)O��7d�h����sK����s9���.3�Qh��`"_�$�]��B!����ud%��W�Xs�0��؛��pߒ\R3@�������Շ�Z9k��;)G��a�duy T���!fڵAt�8D���s�}"<M�8O���݋j�ӅE؈�~`���a_�����)hI�+Q8�:�q[Ig����
ĄHBm	���TJ���ɮ�����%fJ�2#+�	����O�"�e:�u~�/�����!�����Ю>����B*��2낆Oh�Y��+-� ������?�%|l����q�z��u|:�:b�ٕę3Q���a��X��L1y�w䁋��	r�[_�iFY�]_m��]�>O��@�e�����ҹ\[ԏ��8x/�˴n)ƻ�$��]����K|g>�y�Q�\�W
����Qq-Ԯ��t�(R�-�z�Ȅ���%�ʴ��C@�&�� :�}�������|�A��.��j�1��]dtay�~@���7�w[�~��y<
�NO8���B���	(�<��z�nG`M{0�y�'�A�]"
�X�-I��
�p�������n���bmB&?9uF��X%�ͯ������IX�����=���Ɇ�G��vOG%��wp��]� %�lV�E�%NZ��}�Q�a�AU��:�<��Hn_�uO���H'��A� 5�$���ja?�:��e!�`K�¬�-�!��o�`��?��*�qB>G.��z�1��%~" E�YX=N�8]ɨ��S�Lؔ��p�Qժ��HbZ��권r���������l]Ys^eA*�hmH�%���~�L�ţR!��r0��7���(��^e�Y����P2V+��_&�?�gٞ�]ꧏ���El9WUB 'B��W��;��O5���aP�cu�X�))"�fT�Im`��/�U �B��F��ޓ+�<�����.^��m�B��*��X	�K��_�*�����e�0�Hnp��7��g�R��Z�pM(��Z��hU/���$������B[*JV��)+�ՕJ�GЬ�T�5�m�N���h����EH��a���Z�K}�jo�{��' ���9��G�?.���@�P���Έ]�o,: �6Y�ƒ��$Ɯ2�ǧ��c�c�×T��=�u,�{RP�ٛ�PMz���������8#��)���$
��}�����RA:���U�C�aa�Y�����o��8��oaGb^D���5�U�@�Gԟj�m� �Zѕ\2����.a�(�ōJ5#�9]���6�ß��Y���*�2�zg���GՌ�J?�<4Y��^a�vol�|S]i�)%��BS�ܿH$2)oZ���m"h���7g���ۡ��pNF�F{���h�6�)D#��׍��x�����׉s5&q�V�'#���I����&A�q��(�~�ו���#?���v�1kK�yB�!^9]Sԩ���F�$\��f[
�*�62x�C����*F2�F����R}E4k�H��q���lM���q����a�|Ƶ�������-٠R`�]!����P�{�b�غ�zOD��<���ͤ��y����]o��俒I�U�r�<oc�$��E�$���8\F�^��P�0Ԅ�4{(��,��A��9��,��\p��d\��l=j�lQ��0��`?���R�e��x籢�9���J�nt�q�F����#w ���;���F�x��a}�"$vD\*\���;;���/�F��Fp�Ie�Y1�C��"�3>�ي?d�T�Z%�Z�e	�ɪ�E,CI���^B�����D�vD�m���}=m#S�TU1�Rc��w�
x�e�6�;";\����֨s��Зq	�WM����}"�*+�T�ha_������?��Cj���-���L�)>147;�V�'�|�,�t��<���/�;%rr���"�h����ݽ�c��ݮE� j�c�CRr!�]��ϧ�J-:���'wh�ҿ1��)2������\�;0�0�H|vN����d�ۚ�`}���R�:q�� 3��ZF2��3�\�M����v��0����x �]�X�j��� �_�*)��,�Niԯ��{;[�V�k�|&��Ü.3�0i�*�z�A��밡�Hz>�i�4��o&&*'`��0k"`Sm�Zi\���][5�ܔK�U'(S!3n����>r����}X�'�jL����y?�t�Raw��BR�Qe�ߍ}��*X���g���?�f��Z)���M�W�oWt�%Z��* B:���FQaN_�~"�����a2�oH�Yz�5Y3�Z�`~ұA	����f����g��
��vA�7�7̗�G�gWQ[���4E���B�m�'�]i�)������d����٢�����k)��H���'���f(چ���%6�hsFj:���s��WG����2a����H|��^`�S��ڐ���gC#	��SH�"k�S��:����D���2��5wdJxA}l!;��SZ�����edJP^'h��R|.�җ��_�پo�z
�;> bV��m����̔Wi��
�'��+�'P�hR��H�8~�`���;9��F�Nyk<�AG ��:���f́~ÇPw3��U٣��ɞ��ĳ	�I �0���8���Q*�kR
Np����(#(�/7[>R�R'�u�ڂ��\�����K�̺�^���U�sG�q۔*�@�'�B����;Cѿ��q��p� �ك�p��>a���xB�tQ>��2����d���$��G׾����g�#WԮa{�Ur�YQ׷J*%k�A�Ѧj���1��
`�l�D���Õ��-:2%��s�T���45uH]�4#�������n�n�<�9jngz[�g��<l�R DZ�g� � a
{eQa�<���B;y&f�x��Cu+��=���J��Hy.��r�ׄ�b��JX��)�x���p�u䏵ɱ�Q�Qa�@�����3/��J�p�����Ŏ~�1��ҴaSƑKR�޾2Hޫ�@��s���_�3a�}�[b1��w��]c��(����mS�a9��q�wN�?�&,�MRKt��� �F�n�u�ٶ>�E��^�So�nC��u�`$���#��� YLֆo��F�kcV?��-
^���1�d���i=���<�0�h@"�}8֥�ز3j����� �D֏�@��n�U���畄�ǈM���m]N'��\���#7�Y�˕\M�f��?OT��7$��
~=�6&@Q��h�=o�'S�OO��V�������!ʅ���/w�U����s�Z*ꁀ�$+0.��^���������פ����T���nE�aykt ��y�e��\�ߐ�X�d��u-�?)�i t�ܥU�v�>Ժ���KrK� �KS�M�g���T+rb��̖! /�Xe66Ԙ�З]��6=e}�Vh�s���r`]��H��˺Bl����k���)���ì-/�%*��@s�/<�� �`a��V�����v�s�ڹ늺���Z��ƀ(8P���$f$_y��s/,�:\9���7�����EA�G�|o��K4Q��a�7�E�g�-g ��Q�^>�9��u�����������x�4	x�m3�c�^������������$޾2���L)���fH��j�>��~��>EY��iL�Gz��������F�_f��S�gZ�4��ި{����'m��`it*���G�q��c~:H*�@3��3��N0�C�&���b�f��_����&�)Ԏ�8Ċ�f�,�� ����Rs%:k�2ʤ� cON��q�eM<�8�ǐH<���P%0��
��C\M:�����-zi�Ĵ�V(�>+��,d 5��M$qȕH�����ǻ�u��]ݿ����:$���{I,��W	�G���<��L��&�vy��c��� ��DBm����,D�Rh�3��goa��3���(�����X�B*�r��{ QPp���Y7>�n�D9˸�cK��e7w�绖(!~��D��� ����ǜ�B�ͺ�Mf�,S
$����=��Qy�e%q\E��R)T�iи�1IZ�?������ޝ72p��D�A����mVU
+�9��<sFI�>�I�'�Z��^ɵ�*{�L���!�b���/`�|r%:�B-�+8���\4�Aõ�fF�w@���NE����TS�5܇.����.�:�a����ݺ�꘯T\,CZ��@Mg�qԘ�C룷���@.E��:�Z�h3�C]����v���X���s�f��4(�#9x����._�"~U�w��@����&NNw�f)�`�fYu����pȺ�m�0E�k�"����i�p�!t۾7-���9���&�j#�����s�~��"� Kt���w���5А��&�S�ߧ|8�a������#��5�)DN�S�P_���#s�#߮��Ɛd�|�_���� �W��kB��|�{������+�l��A�S�U�eP�9�� ͹�ؕ�U7����*�4�S�OI���3ӷ�N}�� �"��)�C���{t���-��}����~�~�J닮�8�h5[Bt#�şL���߁[�����ڌƸ�=��(�q��;��Ո4	�[2#=>]'Hw�f��W.N�3'?�v) /}8R΅�DOke�P�'��Y᠑��l��@�!�>!����6d����be *@,�Ո-1����&`�^G�N� �!֧93`؉�~'��\�����{��k ���Uۮ���%�Em��n��x�Ql�@��S-;�f��$TI�|;z�s�^��e��vΑʕen�g�rX�5��n�����:m�mC��í��%����8�me��ɠk�Q�H6���^���Ӽ��3����M�&��]B�&ѰsS�����sw�<R�r� �s�kAp���O:�x�{
��J�C�A�IۼV��6�;�d��`����e+b����z,���3粟O��;�]懙�����T�2 x���D�����c����
�^[��-���o�e<<�E��P���?��C&�N DLs�:<Z�� {C�%���g��r��Ȕ(GǨ�V�D�w=�v�+g�?�tؖW����]�7Z����� �T!g�%۴��R�o�������J�C�F�_�8�.�3k?�Ո��R�@�$�S�|��~���i��C�EF�ܑ�d`���[�����ƥi�a�B�3L�a��t�m�l��SF���E�v��ݳ�2������ߟB��iS �o/�����I#v#�o�m��L5����� ��̼6��	�rgn���1(���	���zhˊ�j�^��V��'�Y0��;HO�-��)��v?㺠z祰(�WW2`��A��-���f��fe�g&�W9���e�����T>�ly��9�?
�Z�|�|�%�b�k�1[�2�J2\U�+ b��`�h=�.M&L�[��\�c����t]�@:�%2o�cX[��p�>b�(�Qv�4N�	�84�4b�:z��k���'dMR�?�l�Y���᫺Wa2i����L�;�y�~��P��;�)�ڎ#!��	(T�*���BF/��4�)Y*YLi��mD6?�Q��w+0�fq�u<]���=���<�7������4.޲���l�K�LUAH���Skl;c�mwz�aD��}͖Ϗ���Y����ն�a�8G3��[o�WXH��6.���oa������{Y�ed!�ӄ+�B��B]���_
eM���[9����3��nϻ�g�7���t�a�����[4Z�ઓ|Q$[�ظ�]�f�;�Vޕ���8��a0Ӷ�~�=`�"_�o4Q�G��(����p��zgp�)P��W[�-2�Zi�ˬ����l��z����î��B�7]X�g��`��L�����s/����8�P_�ڵ�X�m)
�u��8�,��kif/O�kvb�Z��!#\�=��J�7�R^���Z"���Ay��`+�J�*����H�y�/�CR�B�K����*ad'��w����A�{0�`�y�Aǌ&;H9.R�>�\��:�5�!�\bTǷ���,H&�I��Q-Cϟ
� �{c����6�ܖ�~���])�ݖ��6l�=��U>�����+;�~�@ K��uai|f�!9C�y�L�!|��rgH��Z��o��a����p+�Z*�	���8T`L��w���ۗ�b�Z��r�^-��r���pO�@�S\���L��\��;N����r��9]j�M���u�ք-�1u�4b��Á .~�_j.
/���C�A�)2�_8$�?M��?�B�{�b)���f�d�1�fuV/dw§V��q,�z�z ��Mb:r�p71�l}q�Me���g�%	��m���v-�>�<ѭ�d�
�I�͚)���� �1%�ov�=����DZ��4��{�;N?���|����`ci�h�x �e!��Z��Sn��}ƤKZv_��UU-c��]R�
���Ew�����4�>�%���Q��c��|�8≉j�Cx�GB��#�!�ٯ���te�6HǑt���ܨ}Z �Q�p$��!�t��3�ma6�q)&L_t�z<C��;�6�q�k	���1t��rp�$��ф��qscj�^cA��d��]�4�o�t����rp"&���U6���?E�F��*O�����̸r6Q���O�5>����(O�����؍$��l��Mo_��H�£� �T��T�����;�����)k��W@��e���ɗ^f��O��w/�X+�D�W��=���ڇ��x�S�		~W�έ�mUѪ���D��!	���׷�{)�2/a������c��1-f�tYNuI!�0#t�4G½����9�GdYf����'\�ܧ6�O��,��lDk@�o����$w$�*#�zR�R��љ�Kl/��ڄ)��ϼ�t.���*�F+>.�rS��s,�oa�;��{<����@u������y���C��k%#��KY,����\�=*��Os��˵��P��$�[��W5r|��N�X2wrȉ���3�3JH8��K��+�Y#%-/������|�7}U�By��݄�U�����q�H�4Ѝcz��Dz�|�%�'��w���������­|��t5��뇊fͿ֥�X��U/i)��vSʘ���W��]���f�"�?P��3ق��Q\��{��5Hv��_e-�A�i���H�*M������c�a�(��6���Ӈ㤣l��?c����
kEF�C|������֕�^�M	:�Sy�F9�(<����b��X�r>���K�$[
8��櫛�-63
��v�"op��m4���K��iy�~w�^}g�J��a{n(]�?�=DI�>�?��o��g�4�7��)\|d�IE�[�==�G ��ڒ��O`�)�ձE����z4���F)K��"m*��>F���q�S���d��/Ә��c/_��I��(����ɒ�x�na��y���P��1�$C=��r��w㠛e�x
t��ْ�p�?��KFTA�{��;E�`<�a(��>Gb	\�k<�	Q�y3e���w���ZeH���v,�˭�q��5g("q��Ɏ|��cAw��U�֖�j;���-Pz��z1.����ʶd�w!�&���x·m��t�#0�2����/��Y����^mGQ�״�|�>��~_qj<M޸"����&y�k���h��6�0 )�(���t_l�f�3�S��1D��3D%��1��A�y�0"�t�xu�l%|���/'Ǖ��$�Ux��DB�v��G.򃫫8��	�������`[�:Q;���2.�9;:?{b�$ ��<M�8�٠�E�=d�^Ӊ'�A����(��d�Jp�c���{��>����A�z���]�vL��[��:�R�	}!���i�aI{逅Wx.�c��J�ң�萩�dK��avD�4�6�mVƺՁSDl�������O<���>�;�J+�{�PV����������_L���e��B�g���mhA�3�����@D�Id7�p�+��F��LIs�����ѣ�vT[.#k�"9{B�ʯ�l�q�! ��ėǉ�_�%v�A5'_��t��{�P��>�4�%';�Q�@��tq�~��Mz�p]Ĝr�`�c �Z),R<���j��k %|R���5G��7姇��2]����cW�\�B h��Έ���l�0�d��҆w�}+�������Xy���� ��y>NE��AN��K�����Q��	�y��%YI�'��\!�_~EO��FM:ż�l���z�>M������%+=��H��R4D��6:Qq�Ե������M(`����|(��J��A%��"��ڟNN�ck��s�I�`��jZyM�^f�-ڴ�;]�%@��=���'� Ҏ[&uǱ�Ly	�pvo��(h(��EWE���D�=�W��]�9��s.����[����Oy[�H�>�^�|�	����[�nW�t=�Pt���S��/���!tWR�)�`�YY@Dg�VN#�C��A�Jm���Oa��N5֣���]��~�ޘi���.�a���L��2+�.}X
/�PZ�C_M�,4[�$�����s�	W�&�� '�W"_H��Y�-����Z$�v��%2��TJ��G�ּq%�C}�c�"���V�IH��٭v�`��0#��t)Oǘ�R�*������EK�-�XeJ��*�Ǥ�BTSMkB�4]������k	 s��K0+���%�ɼ� �I�R"��d׽~U��T�?i�}?�N���ύ�֞�VY���Xv�0A`s�{k���b[i(�%Y�9 I!�]��{��N�|9z�:/��Ls�q@7{Mdt~���y8�<'�D�Gr�^��͟�Q����>���pI3	"����7h�9#�=/XI1*[���
����A!� t>L��?#M��tA�K �N;]Ե�5A�>�����|��A��{���tSZ�v9��՞����k[��[���~�^�7n
1,~ڮC�-�j�����G�d����#;�`@0� ,Y�YV�h�RO��f>��[�n�3�"��(eT��"/�\�������jĨB�"g�X��1�ꑉ��"jc��WH�I�B!����|������ߌ,,��joe��������~=��r��[�K.=	S]��^:���N��Z:x�J��6��OL�ї!׮�\81p����o:����W���N�N��Ug3�Ic�c�cذ���8�߀2�򠉆��@�R��*�evʺ��ZɋR�$K]z�UC��Qءk�����-l�1�����zҠu�M��bH@�hq*zq^u�v>�m+C[���f��I�a�$x.������h�?#]V��"�_�%H��i�7G�.F����W�ʨ����K��V�ס�I���}�9_Qx.ʀGM:�+"F�l˱Ţ�M�$�6^v$��^P�
ZY(o�/J ��0�L�L�kB	�{��[r/{7q~�k&,�v1('׷V��$���|t��H��M"Iɨ��%�4��g42vq=Ӭ�F��7�Ғ�:w�jR��K9a��<h�(�E�[Qذʪ�
��Q{�U�Mm e =�i���ɝ�/3X؍����S�v�#��f�ڊ�l�+"�9�@�����$�lbZ|^��]�E�"*^����ɯ��Eה����4	8zr����_y+u�q�$�s�ϰ��\s_[�+K+�r�E��z�E��[39 �)��X?�w����Wkߵ��+=���N¤|�YE�n�:bΏ4�������x.�h�&��|~�Ԍ(����v�7і��	��M�;"E��A�Lm������p���&���=.���L����o�J��ݧF��1l�ždd7SQ���OO�}粸���dfPt��������:��]�m�b��5����,���/o֥w�U]��8��	���^8w����X��ʐ��o�0�����(x>��8�#�W���Ro`�~'�c�OTf+N�僜l�2WmDTo���(��r�se/�6�A�dQ�S�JX}��EW�����I�˶S�b������������z�5��#��˪\�@���v�{E��]�����xZ �+�p W<v	!�'ɻȏN:��n[����k�.�����)�Ci����O8V�]��pv��L���j���||��K*�:g��N4���4�!��AmR��0�I���]��A�!s�_�5KP��<�щ���S}r
��irj��5����%^�oAD�A~����1�kW�p�D쮪�����AbscNB����V&�l��6��{02�w����5+.6���n3;�_|�"`�����&�W��「���f�V��g�K�&m��R�޼[G?�x��{7	h�@H�Q���2� `�Xy!���/���d��]��,�I�K	�y�c��s�ɽ�� �v��s�rSY�I1��:��`����>d�.�����%t�޵紩^�������)!=eyr9������o66~L����Ϫ�)�K���2�� PY��7�z��)s�R�8P�w��]��Zpy
eֳ��0`�k����ȏK!B1����{Z-Z^���;9��ƨI����YR#��:]Żd��ل�G���[���\Cႆ$ک��5l&Տt��%}K/U����pF�Y��3J��F�T�@��[��QrzKr�2�N9�y:J�J��	�
���Ji�T���4Z.k�ߨ��SV���d���Io�����8����+$\q̃��7/bF��'�7`b���ݨ�.�(L(�����ݥ@�Kt���>rC,����+�����l&G�9��%�0P�}�� �XLQ�m�u'@�Dq������=��-�YkP�����RUK�;��1���Cp=WNx!a����c/nѾ�H+��aƾH��/f�y��ؖU/|��VCNE7H�+��ᨬ8_h�4�ߜ����T�S�=D셮�)�'�d�M���MH�-���q�ؿY¶q�$�E��f,�3�7p7��m2��<�c>����x�m�U�o��fX��p�.���8�z	v�co;z��5�N�2D�n�Y�;��]Sj�>v�.E{���r���fV�Ul[e�E��1�ń������Y׺M ܕW8\�o��v�4��@^��қ)5��T�����F2_���Ǆ2=uB}@;�m1r3���(�,E�=C�n��� v GY�Ͱ��4����;�� mk8�H�/PL�}�^�%�b��]���	l��iu�e���Ǻ]����躙_(�J�`�&k��a�������h�J$�^�����G��ۧ험D��@�{N�醮a/��@��KFD=M�b�/������_pJW5�%��ߤX\ٱ�R��o��14�?!eR��`Ԟ_��*��[=���R�[tP	���ڢ��\V+>��r�vvj⳺W��?q
f�G�N�匶.6wlO0JzE�E'y[�����@�̞�����V{��|�^*���N�9��^��v䧊��t%CZw���]�B�Ĵ��?R-��P��X�~Y����xuֆ
��ڪ5�+�c
��Ld64�ͦ_�aJ�Ip�D�P8���ZF��Sw�=Q�{8rKʫ���C��0j ����F�ea5諘��&�e���'0n$;(VC�̣���)�����B㣥p����F�<^S�7	5'��ىĹ6���5?G-�)���/h喙,b���Ç��8�K�	���
,C�R8�.�a��g��[��z�!������L�������5ڹ,X�W\��ko�{���NRb�k%ދ�Q����[�H2I9�͋��\Q����ΞP�������:���b��>o(}����)i�iv%lٜ�����V�o8�Ll(R�%���k���,1�a�9�#�Mqμ�Xtf&T,�}���w�90���\���C��_�+�G��.dh�J{.pʹQc�[�z����Q�N҅5vWQ���NA�7��K�z��5�_�Q�4u�H�����$`���.��$�9�]Md�	Ϯ��J?�/l�Q3��.�����DrI���.%�����.W�?l��M�#O��%�wG���-}��3��b�qZaD��{�w��$<�)F�����NHX����0<mO�}&�.`����&�k*��S������O��.�({�}���%�>�$n�? {5�1���-�$���<��^5��Ȍ�N�ʑE͡D&vr���ElZ��H#;��.���Ń^%��¶��6U}��1��@ʪ P����:B�gJ���<x� jħ���E��'��>����V�s^�0g-�j��'h� N����HU=��UnG��%���琝�z�