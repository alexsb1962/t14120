��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:��������uA��@��y���<����xDET>��W�����C%�=U����3v���hj��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k��u���ҽ����乊_���q�9�e�������y�^�� s�-&E�E���U�������u�z���1��vw�h��|��KѭU,���u̷�]��ƪ5�~v3�,TP򋰻w!���0��25�m���W���4yw���M{J��kc�?״�qm)�\Ɯ����ʿ:�ř�ڣ#�i��0���X���c�ѬW1?��.*(�M��F��Ι.�t-�]Rpfy��=��\� �!ru����:c�V@��F\.��"�ډ��"ݒ�[X����~ ��/'Z^r��(U8eXbݞ���'~�y�Z�����ѣ���d�_*�!#x�4S��2�Z��;���$22 ��v�p�8|q{�M��~��i4H�2�͕N9B�{�q��	T��if�t����m.��y?�K��p����>݉�/��`e=�L��i	�d�x��i�1�ᢆ��ČI����&�[f�[�{Ϟ��{�#��H�k��|e$I̺|A{������G��h]�d���[�^'׺]x���� ����x��{\��#����`�2pzgM)����"\���:��9*�@c��Q'N��a�3t����Z?���7Ѳ�i�l�c)c��cf<���zə���!ͭ���w#��#)�X�D���oD	�*m�:I�O5�3�UJ�ȕx')�(�HjYc�Y]��`SV��)���*@:�D�ɿ3�􀰮W����丗����૆]�+�iED��9��*�%^;]:�Ў��kYU��FԂ-u�6qX#���`Go�gk��SG�C�?��.�^:!��ML�1��n�|���ϳ�`���/�ScK�K�@��wCb�JJ��2��b�mVm4�� ?�F�ӎ:M���N��� ��0I������{_��8O�T���Ƈ����"D�j����Z)���7IP)1M�>�����}`Y_�^m���T���c���o�����&�����,�i�S7����(���_�s����`�M�q���7�r�7�}Y.3�����-�S��#���8A1���)^�y���>����ظ!�Ag�x/Q�E��C h��`���{7�ӎo����Z�^:���B>V�L)!kR ���U�N~�OJr�8B�2i*L纘�IR��/b��ϡ `��|I�0�*��涶�F��#�K�՞{k��8�M��Ȭ��3g�=M	�0TS%r�3��r-9��Q%���O��0ѫ��k���q�RvѱSǣ���D��Q7�S�
��d.QeͲ`�F�~Lk�,�e>O����gi���n�����k�TJ��^��?�]��]cى��v5C��!�v��e?1�����e��.��{ ߴ��l����$��ls����w����*cU�=\��v0�\���1$�ԏ1�^��ͤ��)е;��0͢|��YVΪw36jȔlҩW	�W�UW0=+ؖ�U���p�� FÊ��Z������#T��>7��N�N�bQ��3��
U�6�����v�+GW��w��r>�Ap�_^U�>Bg��;��a� �I�~G��ٮ0���T/q�0	
b2_0�$�ɒ9m��uP����(� �����Ҍ�sЀ!�NC���xySF���r��?�=�fu��9d�(:�je�y����	�!y�Ax�^����v\���X�i�4^\�&��W�u���S��%eI�>�xez
��j�H"s�w8�֍�g��A���d��+���J�gD�����B��<��0<c�1lA2r%�w�ũ���^E�
�z�75��zS_��(�[R?'V{�YX����6� ��P����v(sZ�2��֟y���,9������ i@B���e�n��Z3߄���������C��snl3�w8�=NN�%���Iu�:3T�<�{�(��y�Vcg�v�W^�܄Ǭ��XІU���{�~�!.e�fGa<O{����+��@r)��q��nr�k�lg����h����U8�.W^��\�A����ӬQZBX+��鋞,��󕚗?��̥p��E΄�>ŋ�͔���5o{H'�:B�бӴ�3���0�,�n�%�`6��z�)�b�T����_���J"��.�$7�:�N�/Q�Y�n����i/�<�t0��W��0�O�"X���6 8�s���_cפS�n+e�Nʝ����:3�N�9�6X��I�kɟ�̏L�՛h��8A)�GӶ��^Q:�AA�j<Jcg��̭��o��Ic+��쌨DI�V����nS`����lip!�)~����9~.���CN�X놷�P%���]�/��Jh�G�Q+���U�����4W1�J)]؊�_[�b���̄�kCz#i�=�cGD��US����a3Jo�)NT;��;6�����]Q�D���!��Y	ٸO��Zb��|�TD�Z��B>�Cw%�?u��?Ԫ�Tg��8]�u�}��-�^82�nM醚[Pkm��{�5���٪�ߎ�M�K�����Ъ�n��v�$�;��q5���1�xƈ�4B0��n*�ĺ@�G�ZoN��C�/�s����<�ߴiCjy7�A��I�K�O���TN&�;��:��FKu!�Ӷ�]Vq�҃��EY�9U�GA(H�[�9h��D��8>F�9$��n��/5�Wtv�9��'ɐm.QǸ����+&&F[X��}��>]-�x��ʥ�N	ci�res��eA�^�y�UA���w��
;^;k?T���X�i�����O�kM�cS�����$�2�N�6�՛lȟ���l���KB���L]������<;v��k��X\8�x�	'����F��t��(�~�V�t(C�Q��n���/�;��/v��mta��L�f֡m"ܣʋiJ�`i�zP�:�h���c	_8[�X�n��M[)V������*�OZB�������,���V�!����1̳ך��	���)�W��'��ҘlTf8��m�� �Z%��L��O_B?ż�KAX�4J�x ��r���%�ߑ:^��"G�jr�53�Ue̼L}���e.Mc�Kg�{��� *��Op��Lb��H�0��P���Ȳ�
�����|��O�AMWc}�9a
(5�^S�nd�Z��[bAG�5�Pa.���Q��ؿ$-�.�b�n\*�E�-9�[�6T�G��"���*�	w'�
���:�G�h�o��ST��	)�(֧�?��
M�fM��ؾ����