��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:��������uA��@��y���<����xDET>��W�����C%�=U����3v���hj��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^(Q�`QԤ9��<8��IϾ�} ��P�,X%��d^|�������6��X���@N�ykl[!�IҌ�x�*_Y#Fx�[����Iu���?2�F�r������[���_��ͳ��Ϭ�#G�G%$v��]]�(��$�f���;��ǘ�xgT0���S��{�.�k�q���j7����dK,�ۭgѩ��t���h!��'�3�x8��Ϡ���j��N]��1]���Rt��<��ۯ�7&?$�0���d�L�T�?�M���F���.�W�EnV��0KF��3��ᆜ͠Ϛ:a{�6��/��Kkl��,�;%C�)�L�~
 #��X�ǧ'�0��q��`��L�L M��v���b�	��#M�
u�;�^QK��'�����}�/�@��Ś1�`�)�ƌ����t��a����Ʋظy�!ϑ�>��.�W�gIu�`��N)����e��1i �VQ���?��Dn٦�F�-�Վ �u<t�7��� �PlY;��°��l�����P�&��dw�Д���L�j�{5�*��~V�C�}5�
�tAv��)]o4��_R�T��?�˟1#�>e�ҝ�So�*4g��/�Ǵ�ͻJt�@������"}8Uc��9�-�Q����j_kb/�=��G�Yǵl\y4o^D�5d���h��M��2|���ܓ ��?�8���$Ǉ�K���Y�h"2�)]o7��v�`>/�q�'�ǻ�k;HAg%E�4G#��1�Z��Habf!Y�V�yʎ`�+��sy�M|<(�+g�.�"=`�&�Cٝw0�ao6L:wo9�F�du
w9������gْ��.��z��/J��$�1������k���Z�6�H�*���=�$�����ݷ�@Ϥ�rJ��[&�&ж����cd���bU�t�䢧�aizci聯(�w<������'1\%,?�a��:w��.�#��p{�����c��a|g�N�˂�>���}���б���~�{��2���%A������S��0�2m�_� ���9o�ޠq�<�����h~(Tw��wVŐ������/'�E��N��H�RW&%�����h;&K`���>щ�d=rK�J.�ꔈnm�l�b�� ���.^��#�~�I�=쏵&$1Q¬�V���i�ǿ����x����vB<�6|��0nI?��P�Je�g;*���igz+�G������x�$���{28�?(��4�Ǒ��fJ�&������^̠CQ��J�\�/tcC?�h#>��J����
�� \!��}�V���7����~0 �:'~:���]v2�����V�R��d�n$��ͻ~�����Ɛ^w��<�?q�Gqf��(OoM�65���_�]����&�� �Vi|�73;S8��ݜ��z�#c�n�cL��+�c~�a���`���R�X��Y�K��M�ߗ���$�TMGɎFL����*�U�S��OJ1�>m�	�Ý����g��fKb+Ѝ���V�Gk �����D�"�$����'%ΘR��؆ ����c�_�#��r�x�ȵ�M���S]*	����>�C3�������d����'�T��؀ �1�:ӻ�A�B{���/�U�������]L��pf}mmӍ`�#�>��O�M �$����U�=�kf���-.O_�h���2��H�']P���(��C'z=�i�|�3��$��ŧ�f�o��BB����Z�F=W��'��~b�z��2�����0�nX4\�x����<!<�, B�� �`A��](Ǻ�VڃPO�K���k�zDW.	b�Q4ڴ�m�N�G�8ѡF�%*]�	�ۨ��pC���~�=�������+�)3XR(Y+'�w-�B���&P4�[%]�����K���c;����~sZ��n��������}Ĥ'q�!A8@������X���HsUf�VP��4&�֚a}�t����Cԍ���Be:���f	3ßh��|S��ʘwvX�f��t�;�B�4�ˋL��z���L�˯��J��c�{b��6��o��=��2%������6���!z�������H�Y}�M��`�J�o����v�aT�wm-k�G�����vWd�4�pqf�ţpy b3]�̲�̪I4�	�Xh<�	���
 ��� vP�v�'$"�S9�&.�S�ב��;w���Ȋ�oI��B�ۍ��yY3�W{�i1���Ro�/�	-�(]�t@Ow�L�D�^��~m���)��u���ږ�g��>�!d:R<�D��T�����3Ϗ��Zgr�a��H������6���Zx�g�	>E�s�Cx
�MD>!�qb;�W�{l�b2���^I��2@�c���Lh�/�H�Z���AC֬2ꖉK~\�l��0Sg���zJv�=�R��x
D�Y(J� S���nA�N(w%���	>x}$�����+]��{("5���$\b(��`��"��J��@�-m
��G糼.7pxQ�Ia�I���e�������4��U�<��tR ����)B�O>�om��}Q�R�ϰ���=�h�yv�mX]ҥ�Z��4�+9m0 ,ev�Ct���P�}-��s�\�M�	0�x5��F:����9��}��	�*��f(���0��;����{��lɉ��{��[0���>���0�Wt�'��A��ǜ^���+2�44��HVvzM��pR%�2+�;�F�-�i��*�~PX�[���p�$�f�#�j�V��z��R���U��N�	9�x�&����7�\]��af�M6Kğ��#Kl��yw����M[K����0�~w2�Q�����x�O����1�[�;�W]�4��Շ'65\.f�5����d���MA��N��E�ri%���y�q�L�qhՔ6ʵ�s�q7�S���Y�pĔ)
�V�����>U^���7ͻ�S_��\�:.p�c
�seO�D�]����3���G��ۗ���s���W�(��m��[����LD�mS̱��v����O����I�]#�9���k��F�Q�dz��ŉ�ӡy����>H�C�� g?� d�P��Pa�A�:���">���#���K�T�����fwݵt�p�^������W�Trz��҃�	�{�/�,5��������	����$t�쎲�U����f(8�*bJ<��U#��f���z6y;4]i=W����l61;�ظ�R.ֹ�5��C��/��82}���}ܠ���?8R}f5���\x��w�(�1YZ�/_��37�'�3ϋ���M��sy{����8ʿ�j^\�\ڦȡ�&������ �`֕��y��s�&ٟ�ς��h�C��.0�����U>��`�	ʣY[ɣ�Y�L�=;H�[��0����KL���{N�HD���<���)UVyX�����S3Q�`9�Y�L"������w<��stU��Y�o(r-�D'01��k:��;~��(X��fCXt����J�v��M5�N
��ن)5��Or�zbV����:��q�(�B����]�3I�����`�Z,ˆj���r*�Fن7�n{`$MK)�q'.�Kû�[͎>��5���zs�S��_�s�QBY�m{Z�.���:��6-N/�浊�r�����(���h���8��D�AG��3�~W�7&okuz�ڈIo�wwL:����j,>�Ǿ�l�Aُ�+�ױ ��A�:�9JM �3:�oL�z���;�t��t�0��*A�a���Y^�mE��I��D�*�'�ĬT�	� \�l{�������5��<�X���K�b��'ڔ�]b��4�Y/��o��\��h��N�2Jb�^�p+W�8�g��t���A)y�����A��FIG���l�K�fvn\m�W��>�G��oOI��e���0��X�}Z&T��=!�e�3,��lp�̿l�;� ����y2<k�+0���=�56������<��O� �u��"��䳟k���2p���[�����'�.k��5lK�`�!I� ���}���`-���Y�g6�?�eC|��L��������1Ô@1�1WߙXQ�45E �54o_rP���M(�VCۄ�.�GA���������Zq���C��Ĩ�=��$&��X�7�W=w��ڧX��O%].�EGw��	��x�Ca��T������� zM<e'6��nH%fu��s��U�M-��1��Ư����'T�S�۱�:�ȋ\��-�˃�O_,�1�rSŌ�T���łw!8�:����n4.�
_��ȓ�n:L� ��7{��� �GG��o���+�TSJ ^
����nh��W[��.�ϮW�o�Ц��]�̙W1㚦F��@�ʰ�;~�[��Ou�-g?�r�FΠ�?�WE�3�᭜h���/[��^��^n�׷O�bĸ2��ڍCk��'l�Z�k���z�,��	���VU���vw�3��)�� ��r��i|u�����r� gM�O�L��{��U�[×�������W���Ϗ���_L܆�w���x��T2����g��s��_������a��fv��9�ą��5���x�I/?o�id���"�nvM����Ku��Z>Y�]��G�V,Ӻ4O��C���w�����'�5,^��\��Q|����_Z�ta&8�Xa�Q�ui;�5"������F�pՁ���v�>�H�ΌX�"��ą�t�	���W��7����9M'��'(�#��
9{״/��e��@jHW�����ٳ	j)��e��~ie���cUg�|Nv�Bع�|eΜ5�I<����w�#�y���:��C5̗.�X��a�d����7�Dz�!����E��J������`C�c��@�&��؄�Q
��wUK���h�o�Ϸ�o�a�:�h��	]�s�7�Vk����V�CET��-�����e�*�K���O��<f���r�(��-��"�c��,�[���2�яq��2�*T���@� \C��L�S��2K;�nk����c��܀w^����z�bfq�Ez��vf�v3��t~9��j�|��j�j����J��ݺ#鞢yݗN�9�e��'2��~��k��V��x�k�Ǯ���������!ك0��������4���Qay���m_�\U0Z�0��~Yrci2��ݙ_�a5�ҭ�XkN�i��"���<x�����ԽN��)^^���H2���T45�;��Y+IB�Gw��0H��W+�'�� �ɮ�Q������ذ":�W��x���'c|�G9���zq$��(\��<��&�ܯ5��ew1d�]T�Xw�|���9*����f4��������F�۹!�dP�~"���ݮ[������|���`�ǥTv�T��N�H�����-���,jɞ@Lb��~�.}��B�>����
�Y��l���L~�������}�����⊥�L'�������n�Ҏ0C�H�k�!'��Yè�F�+�>,Xh�M�Cw����9��J ����eA�O�S,O�������T�L���L�e��?�+ibeqe��J��,�m�.m�@�bޓ����E�����y)r��'��� �:O�0�b���P��41q�lừ�����>�Z����dQ�S�t���@�Z�X��q��t�.�m;�/�v!,�a��7�,�\$�K;��t��#�U�M�6�Zu�t�pp��|w�w����@HF��b҃����cg@�%F�wX�S6�4�MͲ��>��9����cc��E�X�������#&r�Kr����q����Z{wD�	M�c��(=�7��l������i"a)��sg�h�c��(�l�M�䈂C��}n\
@�T��P}�Ʊ�&�J\"��M�.z �A4��&H>��u���%�a�4ļ�H�D�ǥ���L���^�S.z�P�5f�Z���������ښ��f��?��U ��S� �i��]��[��~�X��Aɿ�=@&skz9Љ��q8"$R�+߰�o��)G�w�[�)��$c����s^���M��ʻ-a������i��Y�fJ��W�f���/��`�iU|@`I��;5q��1]�<cx����ʜ��'�31�ؐl���ޟ���S���xO���d�i���0��K3/<�q����9��A�<��*���rX�t7l�Ha�ٯ{-��YJ�Ԓ29ٰ|9�M����'�N�u3�cG��:��ݷ��\s=����	g�u��k�w�-w�J����j�Wk��m�C��SZ'|�7�d�����cRy�����Ѐ3���?�����]�1b.�`��t��(��`P�G:��莟�3�,�5�L׹J�������~�!��r���¢Ō�L�c��.�Ø�U��w>d�Sy�[������ ��'_�=��D�����q*g)F_��;�VҖnS�	�)W2a�!�q �'j�_]iP �\�9S5��2Q�B)�x1��ҍ*��g��T ��� �J�W��{���D��)gEݸ5�����YKz�)�䂨�Uj�eMx$~���q���~�Ff#Mݙ��9��1�qη���2m,�q!��w�䧵���M�)����玑�s,��L����b8un�}����	��l�H�zfg����JC��ʂ[�>�Y��p;�kz�/!4�����f>|�lJq[f�?�}�Ug�1U �?1����ݾ�r�3��f��P�������uџ�W�~�N|�ѢFZ�M Q�NM�%�ʛ�&>f�y)��5�"��%T�Y3��+����!�hZ�>[R'���+���������\��+_���:������j��L�҂�d�M~#�ը���p�}.�u�v��u`P�h��۲���&��33}�t�����4]�\]}���G)髻 8[�5��������^��PABf��j;i|���j��z
𡘩>��NQX��D-H?
̱&<�Y37G-!ד0hB��������o�!5���)�%�#Հ�U���֔������$G"&d�n�t���U��c_����o&u��Zа!M� G[=~Lq�gk�c&��/��!�D	����.�BE�q�5�"7+�B�{B^��Z1���ڕ�l��Eq���M�K�~�a����/?���]}���<D�W�(}��-���P��h@�њu�\>�& �|�1��
����k�b��т��
d��e���ݳ������PL���v�L���V�o��hvz��\%�Qf�\7��z��<.nf'�.����3n>w[8����.n|�;
%P6e�Q���=���%�bi2�P���P���.`�W˱?�b��`e����C���3�P�C��XU�X���O�F�@w�6f����N��6L�1��yn�?sk���	=eZ��g��M\�#~�@�$�Iư �lf����n4B�h�K_��X*"��ۡ d&��Q�r+��=x��	%%LnL	.q|�b�s� ���!+�(����ޖ?���)L�Q.�;U�]�����F6��[��Rj���%8a�[S�Ix�K`�ܴF��e=�$��P=j�c����/*B�H���V�1�-���./�Б������RG�o� ��Ai�K�CbÖ_�����&.���4h'���"cl���P��m��V��3`���X�8|ʐ�$�@ρ˗��x�6�:��K �<iVH��!���)k�� ��%U%�6��.���a�wꀾ<���[�T�>~p�Rt�kx���υ�s�l=s�zj !H����I��,d�����;w�T%��t���A;�����I���lv��8z�a�)��a�Ej���Y8U��HZ���a��"���$��5JQJ��U���^�~g��ƃ��O�AR�F]*��� Э ��z������K���fsxΨ�2'��cK���8+q*>��(l��2vM#�p�6 �nb��	�X5����"�q������	O�a{(�S��:�鐱y��?�$��C'��}���Cc?��E���b���}�hU깆yjͱ:hUW����t!�@)�EM�����=�\0�٣
b�؎ۋh�fz�^s���a����	K�oV�u�w \�����t���!z�m̜W�ēC�_�&֛���T{>uհ8�p:��*�f8���o�z����o"Z��]w��{���$�|�Rڧ�{���H�>�sA|���19����@4gn���B����Ke0q�����`�~�i܆V��� �f
8��	�:�Ya�=���&EN�z�FB=;�͉�cim�IYvs�(�`ߛM��J�o�����q[�i�/S�Q�M���^�[�w�wK0��f�2x�O�cb�Z�0�OT�<%q۳qcaz�]�b9Lw�����BZ�z���J��$ч���@Wřf[��<�)�x� P��I�R.J���H �6z���w+1G�X��{?&cեS�xݫ�4Z��1ٞ_/����B'�͕��p�"���n&xb��	 ���>I�AY��\Y)��v��[�Q�9;���&#��?�ƞ���Թ����Ț���oj<��|����
^����d2�.u7K�]?�\��O���6䅀Q�^j+��_�G�u1��*iJ���{qOI?o��όdڍ�`1�¥o3���8��� ��0��m���� �e�z��f�z����ݚ]��J(9�5<ؾJ�.X���ѩv[�n�$"xW�m��`Ғ��g�!U�n�֠Uj�g@�8������L�F�	��Z��z�[?�1�9u���~ʒHI$V�bn��]�� �̈́6 d���R���d�g/>�Òg����*� �9=�<Ke�k��I7%�u �S���������WD��x{��̂I�0���+�k��h��:���&	�!��I.��W���U��e�2E^��38�cl�Y2R2�.Z������k��E���3T�'���2{&jn����eQ;�L�6Ok0:�هŭ@@:�W�W)�K�g�mG՜^U=Bq��8�ً���\��Է����|B�|q�8q����gh�C���N�	D�$	vž�`�#_W���Sx�_IX�P�����̠��"��/����(�qvySi?�$�����|Td���&o�6�C
d?�M�y+i��_ٰ�V�q1H�J��}��_�.���Y j�a���i!��}5��$?�xNХ}�WS��܌��e)Y���{��h��;�gM�1��a��o��$;1���!�.4���(��ξc:�J=\������m<����zK�����Ņ�Ag�PVb�ju�
�w���;���
�.�h�) !�0~��mN����� df�wz��:+��u����9Mo���@�p���:E�z��wd��Y9n}b-�����.0rRx-�8x�e�"48��!�cn�p8���95�I�\T�(z���NE�k�TRJ/��f?�V��5Ftv�����L��Q�Q3��62\Ly�<�tpM��� ��2��)��B��������9�ZR��"	�U뢔�>?��
i>��X*�2�oڻ�B�����EA��Q�c�#ғ�K��w��@-n�*�7Q�Y)p��"�N�z)�:w�d�!�=��ĉ��hE�	����AW�l��䮑5�g�ż�(�BYB�
R6z�w�*�p��fY��p�sd ��%��BJ��h6#�#s���hC��x]c�>��V��q�"�rAB,�O���[�����Wl�7�wד܊�æ@�]����ﵝ��	�>o�Z����z	��.�Vȅ��+�H�}Ns�z�"g�;����[�g5W�����3w�f�`<��Ӷ���Z�w�A1�`K��9�v���{k���RX�W2�Fzw�:=����y�s*@� \;�I�"��E�{�l���o�>;�}���܁��5��̆bz�I��yٲ���A�/��ׁ�ᰔ$�j9�UI�5*���#�G5@���D2�cUK[�u�et��~�����IL��1��V���t����~Ϸ^�N�(���	`t�-f�K���<(㽍g������}��Kvn�BQ
ԓΒ�}1�ʣz%���@L$���K<^Zug:Ԯiv�T]w35Ts�k���Ŭ}yբh�.�qalŧ�N�a���R~�f�Y[�Ej2|�9���uZs��L�&��OR��*h ��L^й�!�����k2�/���!�h��i��]�w2�._L��x@����p(�#V߁@�g���x�5���~��D�?�$6t���ϣ_ӂ"XgFxȣ?,���F�������QÝ�y �b[)����7��t%q�뢒��t+/��SqrF��Υ�P��Y���,�=��R��J�@�y���ߓxK�(֖��V�r}=:[�v�40`�NdB�t��+ o�6��e߾^��f`��Lϭ"�@���e+�h����욚 ���߿@�o�N����ζ$M�+�q
�'Hj���:Z9CvJ����և+�v�.�v)|K91���!�E
B�\S1��u���tvA��LMeÄ!G�2{��V$cG�FE���ȕ%�4���#e���v���J�����~p1��e$t�{�?˩���ü���i�1�MŜ�����(��<|ʯqi�X�Ϥ���S��>u�N�5���b%Ei�lH�)E�mH{���)��O)�IC9.P�w5��>2��HX���_�(�Z�Q�ŐC��p�fv{�j�[�c3��+���@������Ll�v��Ǳ������	IǺM�V4@T_���m�8 	�J�j ⰽ��� $���� �0�5��Ƞ=Q$�3�8_���i�n"�v!P^AJ����^���$�v��@��f0����ѳW�S:Էz.�+�t���뿶���ݬ�
(1�kMc^w���\K�b�,m�,kI¥��8����O���5h�����rm9�g�m&��@݁� Z|H��v)�ѐD"M��˜نe�.(�X4�H���q���xBاV	�j�uZ���Sę�_�հ8�$w|��$&�VH�85�o� <:�B���9�^��V2iu�W<5D|���|�T�I$�i�~"��0ȷ�2���u��NO��<5V��a&bt��g����/��|}���I��%
l��$����N+4o��i</�@��U�1��G���2�u8�ZDg�EjE��֪0Z�j/�Iji�<G�r���`��������t����&��~¾�	:2��?�iG�}B�=C����e0}��V��ہ��U�c�,6g*(2�K�"�L>�'Qa�����D^}p<�Vg=�;i\�V������;�f�3��������/�J"�X����kތ
�ܶȭ6����D"����@��(>_�J�N	֌:[6�%�y��ѽ��X(,��U�oFb]2��s�ş�,t�
�a���y[��F��c�56)�ң���&d�c`$�
C���u��{c40D= s�;C�CQ���**��c4C�Q,�@������v_)��E�:���\���gB~�(�Q���������J��1�.91_��zv+�/�ƹȺ�RTtLX/��ke��}4%�9
���N�y&-o�/z7l#R�Ҷ<��� �vN�]��ãfQ�$�B��,ˇ�<�޹4F '��iu��3�p���(H��Jl�U���Wm_#�����v%̯-���3&�7��ɳUB�c��:�lk��,Ywq�y������$���e�#���1��]Y}�N�,������e�nF+�c>K���@~JJZۈ�I�i�C�Ǩ��'W!� R�*e�O�c���� ����
X��b�,cƕM/`a��^��4bU#���O���X{�!�ʼ�!;�oX)T$g?�Rd�*Pt�۟r���y�^ϵ�Z��'_5o�h�u'zq��ԥ|u)�2��=�h�km|�V0��._��z��b���s߆F��h��FK�SF��_b�Gz�'%�"��JՌY�#�N�zOz�#��F�ɹ\����1ҡ��},��P�H5e� /�<�,9�e�R�թ����Mg�Hj!�}�Na���z��R�H���4���׺16up��VR�˵����[�KG<���kp�@y2�^m_A9E�/����V�ki��A��:��˝�*8������E�:�.FJwq �5'��S�Q1��L��H8��R�x�v����0e���|x�9R�6;���m�Jx�;�o��sN,M�r������G�N�\�4��KV/N�_P�^��d0�j�pN/}q���D.J�=-&8�m#n���)x�?��<.�L��m�]�h=��x���1=
��V�3�&��/ݲ��жCT�k/����ʒ���_6��۱݂�H/�$K;���y���osÜ�쁖t�ʅ�|��Z�z��Ԝ�vRFQ��ڹwR����I�w2q���2ʏ!�<�)�00�e2�B���N6� ��I�z�� DsAS�"t)?����ܘ�g���Yg��j�O���=	��3�6KKϸ����nw�X�)Gn)��.�9�~0-(�_��Y["4�m�*��}�Bߧ#��f<�=�V�ַ +�c^	���ci�:����PY��\�X�a���=�� X�O�w_���j+�R�zt2sӳ��hZ����D(�����Z֐��m��]���<7�\q�/���@�h�L��k�H-��9I�ګ�n��o��xsj0�mP�P�=D'�Y��u�0p�BQ
��Mc�YyGu�?�eB�j��prl�٦�?D�1�O)v��a�:ܸl�p��\����Eb�=���57V���+*��疵<���,�,�>E�3k���HK\5�8�yVU��#37����:����	w4k�������s�l�ǧn��3jT�KVWW��7��$9��H!����d��v[�Y��%:�5_yVJa(+?f9�
�K�韘��-O{{F�e>�b��~s��xܑk�9�{~8��
�@W�-��(I�A�����@HI.<�І���I*[���\b5Qa,"�9�I0>_�05ޅ�n�Su:���v�})=���Dg)��[�뀮؟�mֹ녌GNH
�4a|%~���A�ڕ�[{��R�.q)���S�C��NəSCҕ*U�O�k�������g���R��c%w�d�<�>�#B�I��rz�U��ެHp��3� ��e���G�j#Q���6�����ϡ�F�������^���}]�
G�)�@!�����0�3j���mJ���.b��l*YZ����Q�F������l�}�"@��]�<�_�!1ɋ�Ag���,�Nc�u��=��a�VJ�Э��J�Ie��b�Ē:T�)��&�)`"�<.�H����׫�&E3�a�Ϣ�Z�pe#5w�N���e��w�;�����+�#�״�ŭ��U� ���@��
gh>����ZzaGbe���j0B˻�z2&V�e����0�	����j�D8dDlh<|�m��0�l�iP���{C�5/r#����m2B;Q�{/�6�/���y �;q(e�M}�%AʤQx��$V5}m�	,T[#c��p]�yW����ʬ{��{`(���yH�r�)rφ�!�V_�>�� �9 v�hpA������FpA���ՖL�m/Q�C����k}z5�����O��2��B'g�<��I�w���cb�[)ݎF�<�9�><"	}���n����L�oӆ)�*;� �`0FE�\�$�}��ٛ�`w�QB�z��M=�������c��%meʟ9��*)S�ø��$���EoMb&F��F� ��HZpw+V�h�FSq�@S�B��t��+U�J9��ÓX��rk��(�D��>�נ��"����XL<����Gߏ�՛MR�f�΍��C�]�K��
�K1T
�.|T�1lE/�9�j� 9`��1�|�D�~B@K�x2���T�Ƒ�aO��m_�:8I"�ݜ?���T�,�)c�q�Z�08���%���Ni"�6�hO{����8xGj�m�UK�Z:��7�����7�Z�""L��N{���s)KO��=FM���J�v�1Y�qM��ב��m���0n�G���GPtb�l�ɒ|����0����H�ʟ��	�Ъ���"���OV� :c>��y>�N8B����?�u#B�%C�+�y��
4��߮�&�=CV�i��+]-9c6�@����.#���.�ui��e�{ˋ�5>�`7��<���Se�N�� �lu�����!�j-��9�:t�M����Fת�Q%YV�q���&���l0�{�"x�v;}�|pSmR	�7s.E�}�Z
풟��'D9��mT�3�D�[E+A�|w#�H�!�3(B?3�~H���TUz���"׃�k�`���C5�ٿ�O7[��[��dL�c�h;��a�O.ڜ�����`㇠gct�Ch>���?�!�W�I�_cRbv�|iODse� E�M@�yX���:�{���ư�vbu"���f�K���3P=���T�F�KT,�vO2�/�m��a�5OUll�
�*�j
"C�iP[��N��M��Z\��]=y����F���S�uH� s�RĔV�x3����/�p��z�i��4�Y[ED+��3�H�w8{���ӥ�LB���iU��Q�lX4|n��O�~�2��?�Ũ�闵�����+�R��cy^}ĩ���q�1��c}	��l��l�2X�t�[�p��D��]�l�J��g?,��qP��j+�]�2��Zh�v��W�;�����DkCLC(lJ�/��w;cX��jmD����md"�P��n_��G�'�q�q�Q��;�8���o%e�_�8��ϋ!�x'���ք#��	��:*v��M�V���B'0��t�E�d�ZS �x�>���
@��dd�YU�]EBEO����9G��M�ʵ$��KĖ��?�/��۴�� &*K�5ku�)Sz݈�.:,M�����"���0�'�C՞�+ljhӿ��g)x�bG{�^�T�n�M��5�9�.,��Ŷ�]�D�95�r����MQ����z�#R8� ��1<�N!�a<Q�{X����\![.yR7,P�~:��yj���P��|�!�e\�!N��_iSg_�c���
��V�c�qH�ʁn0z�w�x���E9'vWغ��j�#�e}T�}d�Zb�]Kdn���V�1���^*�y���F.KT�F1w�%K-�,��{I-Ba�����8ў�o?H�87�O���M��8ot���ǝ��aKlq�v���ȼkg�%���~���9��%��r�S�8Z�l3��6/��-IiJ�-p2������Go��7�r���㳿�Ё`�E��j桳L���!��s�.
�+!jм"��y�vV �R10!=lh�~���H��S ���k���v�6����;�gSC�@�j�(���~?�5��� �A/㩼�ug{�4�c�O,�Wv�SFP��W�����U���W��Q�˿��SZ$Fa,�e��$�ڴj��W��5u��I
A��0���!�V�j����[�L�W���������t��L@>���;��s;������ϔ�Pnm���y�f	0�P�h�h��v���(��g�qQ����'���^���l�cd�l�x�7|��m ��sk�{j�Z�	�����6�N�� C���I�v�T��+�A{:���LZ�l|鉋@d��T�@�������Nz~+g�ğ!���}�Q2�����;����s�]�J}�+:��ܴ��LHdW5<��M��M�%����b�;�4F�F�Č����J�]�+{���w:!� \��6��s{��u��F�����"{_�|x��?�6�B�+������w�-UE�n��O�2�$���T�{>�������O�ťG��?ٍ��|EA��<��佣h�8w���:&U`:�^^�Ks��[5�=*��b&��O;��z���_?*�)~���p�Տe�5:`��G� ��-��J�6�B�lܔ��g$���zU�Qi�S~���Z�ҘZ�`��$���f-�����%��̺�)��������^y���H�8�k`e�xڪ�z#?�ί��36M�|M錙j������t��1��@	�������e�C锛w1�!�LR'Ě�O�{SY:.�&������8��Q������5-P��bJI��:Q1��C$��!Y.e�������qݟO� 1X�
ֈ��m�%�VBCP;U˻�f$�Œ�:>s��X�=a���w�Ko`���Gľ#���fwIj ��)N���Q}��x@��yM��o^��| 7u#��
�����#c���HcOZg)��^�*�Ą��G����'Vg���m��&���+�\�}���9�k�=:P��/L���v]Q�ו��_\R����! F���3�..v�ܣ���޺�{��6$\_�hr�W6���v�� �V����ޭ��f�JD���K�e�E�� js[��g3�م�߆/Qؕi�xv|U�u,��90l����<�l�~�.X5��(g�-=iUק�q���	`wn�ɕIQ�I?�VPh�5�,92�i��üF��O��=��o��k�F����8)�rq�W|�fb)R<Z�$|Qc*џE�f�+��m'+���2q<7��Z������L[נʑ�ʣ�q�*͡�W�|�r\�sN[QebOKC-��S?#>73�²*x���~*ceІ_����N�NO[~��Ж��t�}v�γ"�.>��M�����ch�&sed����%��+��͐�Z�J@1E)I�.���vh�z螗�/X|}OA,��E��҄]SY?o��<;8_s���Fa�ɵ˜O�v�l�֡���
<���>��t�����g�z x���W1I62,i�3W�E:{62�O�YI��S�=�l�r�q�{�{t���|��M���D�p֞��MexD��Cls�����4<���U�ړ���*��O��]�_D�ٞ�>���w���ɩn%����4:�:��[����~�(���eE�i�����t������]v�x�T|��0�&�if��M�R��o���X�Ӑ����e/t�;j8�R엘����Uch���j�$&={@��M�}/�uh]�U��R<9�$�Ь����
t�d�h]�08���巄�<s�d���kn?�ܶ��a�n�3�z��̽��$�P8f�"	�*�����D4]~�14=�9s��^}�
�WIw0��_�+�N��?��M�P�`�ϑ����{Qwd�hZM|/Z(�+����Ӳ%��%/��ܓ�`�@�%v��.�7z���3W��E����0�D�x� ��<p�"XO�L5eӓJ.~�b��W&=iknm�U�v�׺�H����^x�r_.�'4���U�_OB��]7���(�hN��Z4�oc����krNĽ�i��#�;v��B]�9��?�^�r��?QF�)/c^b�W�R%`�#6���T���2
��T�Y~m�sz��Ā�[�1�G�����GA��MEvsU��4�������-����Aa:�Ef.����d�]�b� h�"�,���F��sC�[p�!��ϧE�I<j�Z.�L[�T�w~@�s��;��"������"�t�'���bP��f�3�5�f��1��ɭ�J�~����;���q�,�&ypa`���t�=���72uJ��CŒ��.�	r���PB��˃��Zyl���+����-h&:e&�|,$�H8��1l{���O؄���J򄳋5M�]�刭/��_]{�^��V���OD6?P�ɠ�\{R*�0>�@��J�l:��z-�e���~؋陰�a��3�ȵ\)j�Ej�V��[�܈�~+��ܟ~���P_8�etZ���f,jk�d߉Eɶ�$S}ŞS���X�����k$��@�f����*=ج�l�;�{k��Kt���b)ic�1�z��X&!�(�r�	V#�ʹJnR>�`���`d4�����!��`������[-%��<��N��G�;��l<�Q�Є���,#1q��Ֆ��@�,t6-�-p�!�C�a�`Mo
�GQx� U����-Q%�F�������%M�ƻq�o@�x�$��GDC޹��m
��	$ �0�Yy�zN&	�x��jU*m�Kk��c�ʹ�94!�Rlұ�dier�d���؇�O�S��ޠ:��ݭٻ$�N�`(�C/�.�OP�0Rtqo%螃Ts3-v$yj�b󺈛X�Y!as�֛�"�����(C�f�_��X��gN~!�o\F�TToJ�'[��T$Q-�1e�Dv�S罚�3��Z�'w ڣ��<����VU����:;K��pr&n�~�a�8�\�yA�|6��
���GXl�S0^����V�Q�A��:��ô9�:����<����kI��S.�έ�Y����:�/�����B��$|��'��'�jVX0�����M�)����x���а�X�N@䀤ס�9x�_��7�����7+��W�JȏzA����?'��4��a%�Urq�ځ�Ϗ��\�����&���ݎFH�����ٸ'@s`�s��UG}PX�6Ι�Q)t�nǀ��A�V���7�?����I�P�?8�~�'Dg%�!��|[s�ޯ��WbH�g�^ї��p�B�ԡ����V�tM�f�w-v<̌�]
�
1ȩոi�����b���>�(;�t��d����;4�Ѵg4�V.Ҩ"�y_:d�;0�F@.`����
�v'p�
}��Ը������s8���%�'�@ݥ:���GV�@���B6]�����ȓ�e�~׃'//&�'2�L��>��Ȝ�dGF)����s�#6��k�Sf��t��K� ��g����aiy��#�Xl��ݩ�D_Rb}m=�7j)���+?yI�7nw���-���DW�n�����B��j��/l���g�7�#9�Ǵ͋�]B�Yf��6v��/�w�ޚ�"�x=ʰ6��c�1D,��r�A�<ɔ�eU��5�$�1�+Z�ќ��cP� 9�!`A��䑞�BR���VȾq�O�-����0r��*dc�ǎ�~B�<-	��̏Z�����$��\���T&�P�ܤ-$��i/H.�{�L�w�}&&|9�W��:��Ȉ�+9��L��R�ڤ(���~ϬQ�#�cSi�����)��̜1��c:���}���_gH!�M�0���F��R��8nc�,1�^�c�{y��n�͉h�@Co��̣�&"�ݓ��_.��'��F�� �Nm����,��)8`�hqEC��I�wۀ��T���A���Td����6�îmQ�
�VM�PT��W!UK������e3Wjf�k �Tj䩎�qZ)m˄�����&7 �R�%��@-w��9���Cnһ���5w���G�� �FB��f�.�qބ7�)S_/Bd��6#-�]�(?Nu�h�K��t��i���W�ZU���d�*�-������v��:�j���lg� �n������SK~�����߲�U� �X �w�~����Ѵf�l��\nr������l:��׭��6f]�$�q�YoI�VJ����B�!1��Z�vr�R�:b,��:;�å��G�O�e��V�w:�//���ݜ��%���r���H�������������F��ؾ�JZ�#d�5�>�N����N`N�FCU�=�ђL��{24>^4�9�HD=u�]N���w�D�2,���7�~���*to���g��"�}�fV �&�9?
�߅��K(�A�3����K;����e�E����q��K��lPNc�j���ͪ�P�џ��G_�����wq���͊�;�<�x{'=��W���U2�Ku�8sX�-b�+ ��Cv��y������7��T��ȭ�zU��|�����E����a����
��Sj���<;Ѝ3!��.�g߲�R���`���?��S�nn�����p����CЃQHj-��ᡱ��)\�
���Z(�XoQ����5ٜV����-&��#����~W�o'��e�[r��bSڧ���g%���	E�00�XB��Қc$HT�aw���/:h�����չ0�俋y\�r�^�k[I8(���#��H�IE�P�'�Z�Um���X.�Q�I��,i�E�$#�,\�{�x���.Y:t���*&�<4ؚ���k�y(Zzn��5�N�J�
�G�T�#Ϝi�*��t����5��.ɋ����l�Yt�N�6�0뉅4�!��:�xJ�w�[������<?���%Y7@T���ժYZF�� �<k< �����z��mKty��G�� ă�r���>	^J��KdS�s�e `�����5�V_:l掶]���K+�F����&���yЉ�bS̈́.�<$La)@����8�E���w�c�<���O�hF���Љ�g�z�����`�;���ԃ�9�ї�.4q��@!P}�kf�Ǎ�C\KdbU���v����,=&��*W�n�w���r���� ��ЅK�� ���a/H���e������\j�YF `�n�4x�H˪�)���*A��z��)'��#k�c�p/Y�_}��ԯ'x�x_�tc)�j���K�`=���n���rD��׃"A�)&9�=&ɣ��)�����d��`��27�1�yЯq����M�~Q�@��-���L߹�P��;[䭢�1h9NB���U�%�_�)�J�DZ?O�2gõ0x�O�£Ey����:�Jot6)0D�ݸ ���W����A�N�Z¾�-g�w�Z-N��M��Ky3}