��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0]��?l
�4�!�ߦ����"�p8"	~��kB�J)��NbM�L��\jO��#y��r�3wA�y�}�S�{�����X�.m�lM(��R�g������B�*�NV�X-?����$��$�3�s�`;��y�@�u�ߗA�R�|�Ԝ�+�)]f��������҅i[^�"[��t��00��6�ĔR�*[�]�V�t���9�c%kz�Q��*N�| ea�z ��@������mU���h�$}���~�k��'C ��� Z���>J����ׯ,�'��3@akCc�U�U��?��a	6S��K󊀧uh���Z��&���9�+�)�b�В���ɀ�t�]z[��z�/`� !g�!*��P�����I�<V�� /o"�����@�g柅˳���.���5����9�i��)�!Ҏ���f8�vh�3�Z��ZC�:3Ϲ@�+��&�Ư���	��������Ϋ< �����"�����!b�'G����Z�!�R�l��Ã���3�����y���H�>����/{���?R%|��n6���gJ�2!b/ΧW�}�/FM��%����� ǜBk{�.�-�ّWz�*J`����'29�05�J�NYŪԚ��N�F2���������q��y�-Y�	����D�0���7��%��,�-.�O,P�y�w	�	�JT6'�Z�Ҟ���4��\��י����Ə��g��y��E��q�"�ӊ��N���H��`����=l�r�Ed�tP\��� �c�G�����/�('�'˷5����+��3]ʸ�:xõ|D,"���V�d�@��^Nm�D�dK�+l����E�ȟ��_��O�՟	����ȢM�6��������U�²��;偐&r�+����q���_j/�/3Ew�?'�Y���7ϓ,4���W�X�`]���eop�B����nIN�_K�����+�-�J��^��8��c�.)��+eR\_�-�/��?���}��@�|�VBp�zq�4���tsT������wPφ�(�,/��3�3~����]4�_x}����M��t,�Wv,�,�t����#���ιXz�^U��#|n���q��LlW�'_�@aQ�Ѽ��Սu�7�q��"�u$��NɌ<�}DZř��tW�	Feei�iH�_�.+9�-�����Xe"����=n0=�~9e/�B�Na�L�e�[�	�]��Z=5D����๓�^�m��=�˼�3A0ba�|&9�7]6���{Qj��M9LAT)��q��ޓ�f���t�1�S�\���8g�8wb�q ݖp�&Q��=18x�w���i��T,��"Ef}_3����u�*م�𯿁���zؑR��2ie�[{�`�hy�8!�Di���4\�q�����$�6�S�P>eR��h�lim�WBb�&,F2,mr�(P���A|%X��n�Ԭ��~���K��c'���_ױ�u5h:���d�"�aM�l���0�k��Tm����$���#!eM���`2T������ǅN),)�r������,�>S���;��&˃�[!��ăj���g�#A{�У�x7(1�2�&��ޛ����I(�0d[���:�ܡ����0Fa|���nS��q:�Wd�4��"�s��MB p^�1�WRl�W�&�\��X�g`2��[��`>{�����p�^���{�_	P��_fX��+�5ً���Ky=ɺm�E3?���8HT�pD�ml�S�5�b��/k�2@o^*�=�����b�����o�a�z��e� k#x�nkk���K����t�8��ZS�r9B�����MD�wN���b���C�ו��'�o��*�j�O�*Ǵ�3;��SE���5}i+�]�eg��:��IE|�����*�G��S���qO���N1���TKt��2����n8�ՙ�n@Rq'���+��%[⡧�g&��~�*��}ت����$���@�nЀ�d�wV"J����\���lCHVyL���7�����j:sG�v���݀,d�,&�D6Ե-��gߚ���y�l�蛴ۮ�7�`�������Μ����%y����$K���l �ӖƮ�U��8pK�y;�x11�P1�~@�;Y�A̠�+�^�M��|��7�v_�IK�0�����b*�-zY� �p�^�;�L��hU��
-yި��Q�����\���PίM�ɗ��R��~�X7yHn.!�ƚ.ǻ�Y���0~l���/��c(�98�0��:�+��8�r�cF����d,Zo�_����\Xٛ<�`b��;��Θ�g��D�._(�j߇
F�q]�����F�+/�~S�cǵ^��}<T4ޯ"!4vJi������G���^*�4Z������LV�| ���c�.t��{Y@�4p��	bGz9�F=9Ƚ�ha����<�0 M��Y>2��Ϫ���