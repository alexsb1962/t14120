��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�
y>F�Gϋ� 
��*�4QK(��7$[M3�E �N����,/mY���n~���M�ȸ��� �i�ӗ�3h�`D#����V'���F8����i(bʭgU��1�".���x�Dc��*bn��Ջʖ����h�Q��ߒ���iq^����pϋ��6>����������|uvY��:(��z���(�u�;$8��.�-�4&��{�G�����ӝ��)�v�l��'N�O��Լ� �KqT/Z�D��Y��B�tH�Ța���v.R�Ps"(9�W����@�[i�<�%f��Q�CΖ:��Ð�Q)c�p0&Ȝ`3���e&����&|����H�#��{N�S{��ڧC=��������p�>�������P��'���z�r@�=�Ҷ��-mH��EC��*8p�M��F�,�9ۀ�@��(���>�����.d��e��9����ɈIL*du��|=k�U��0{���GFEa�4֜�G�˅Z�z�YEV����1�FEa���L��:Ǭ�����%�9�ڽ��nIf%�bL��=^� �'t�VL�Ψ�Y�}���Cdר[<B>��rhw������C��8L��;ղ�n��$���4;ƨ}wӶ7�7����:��IcA��t!���ĸ��9M��z�-�L=�ϟ�M���4����tA�����̀x��u �5��k��=IP���J���������H���oq�1�{���5��׹����w7�����8� Z�2Ծ��ӳ��W�)���R��D��Fjwn�EJ��oQz�@0ܭh~�GX7Uch���n���)��:#NG�Xh&���@��W�Z�-�k|��'��5=�{`���!�-Ĩ ����:�^�J5�4���>,ab	^�H(�F��c�������4������|���Y����KAv1�_;a����pK��=���@�2�Yz�z� ���R�R���yc�HH7�����?�.����؀���8�4��q�|lgN~\��ʫ��:��θބ4@m��S~��"I	�O~i�Wv����wY��R5YU��Bzޣ:���d���3�,yQD��D ��2Ȍ,7�8xz���,����D�ލee��eS4io ��'����43�qM�G��֦:NdX�݋��&a���ݐ;�qeDZ��Vwұ|L5y<u�N��I��G���'peԀnK�s�R23��6!��n}�Uwy]�6���q��1�B�F2�_]�p��=�M�^-�xCR�r�`�/���5���zZ��>������F(�p(y$Tv�//N�8�����pd�@���M����`�v/��_��� ����b
��0&���mNԄ�5b(���]�ssP9N�:��@�z�b�(g*��!q�'����5�eO��������g�U��Lf�Z��)Z��x�<P3��(�ѭ�A��(����_����(,z^۽���@�&t�������yL��%^V�I�b�ctOZ�A(v+%�D(	9BM?���5�ݢ��|�mh�v��'jBh:�Mk�_��i�?���I\����ŉ�AB�p�֗�׶r�Ga�LpK���:k�������5�.o�u����`�Ō�Ǡ��(��GI�AѺ�Z�{*Hmv�� FT��r��ca�^Ѽsچ�*��k?�=�II2��1S7�����1F��8���%�@a��\�ųF�Q���pnㄚD���«^H�j�j�m��󲄌eR;K������������ۮ݂q؝u�i�~N�^�\G�l �痘!�������!�҆������z~I˥w���?�Q������I��+���4YKfp���)�& �X�����*+�Ĝ�� �~#�O�Jӂ'!K��o�b��{���5;�0��S�!��anP��h�Aa����	���f�!�r���tYGp,;�Ǔ�Y�%�2|�*����{�N��V�m"gp[	�(hj예���gR*�f�a݊�CLo�jLb��p���xHc-�
�u����Tt���+������>u�y�Y@�l��1qu12\�L8���Exb�~w���XO����C�L�A�~�->�<��Ie"���F��1�|�|j�I)DzƖ!��F��[gpwB����%��k�YxqXv��[64�j�Y�R��en��I9�* D4EJM��:��|�E��)GƸ)A_�i�=�B��S4�[�_* P�
۬h��@o?k��脅8�=���<�c��AH��a��.z�y���n$q�\�9��,��~/�� F�����ȳU�^�I������S��E�p����=��A���RZ/�>�[�n&��L����9)$_Q��ѳ�+8@68�w��6���b�Eŭ�>�����sCcԧ��t�G�G_85��}�6x(2CW�d#[�L�����f���X�(�jn�r��Q��^w�>��Z���1�'�'x�#����bՌ(��J��0�Z�g�/[��hJ�][3�p���?+��}�OOLZ��Q��06����m��(sW��"c4�B��X���>!K��te�q��<v�!<��A�J��#�q���=n�X�D�}�`�r�b-�%���5�7
���f�;��8� ��-�1�?�F,�ŏ��e��fƷU�}�:k�jXn��%pxvzv���Dq9�e2Wb�3�҈�"o�z�T��$��ax�Kf ��P�����( o4~ڎ��@�\/����nI\���vjӫh[H6\	B�퇵��ȝjM��]����x�y�sWM̳�P��ux绎��QY��*a��=��y��&n�=�=�+��_�l�������4O�ZZ����j;�1���S�Y�b�`��:��������"%�_�94�!�)��V��G���G=	�w����ެS>��O]�"�	Y-�)o��`���a�g�P��(��f�k�f�AW�PV��!�^�
�_���J�I��iV^�TY.r��+E�����怫�ȸ��!W^E�]�-z���b��ӌ�ئJ�z�4xm�'K�@V�H�x�G_=E��^&�ƕ��?{]M��C�(��A�V\�	'+)�n���*�F���C�i)��r�Ui܈�FvG�HR�;lC��-ɩ.wx
Z+��'d�\��<z���-9��Xq�#5q[2z(�e�-�8����Ɣ1��U�jv�%��'�kT@K����A�)�1��?����ϰ7=JLr�����]���_�����`��C'F	g�j����:D�|�%9�t��i�xd��a@�5/y���$��!��]1�O��{�z�F8�Ҳ�Y��U+@i���B
X ������� 4�s	����~�N��π/H=۲eF��,�MY�j����GC�"6Q�:-3d�t=�E�&T#;6��}�Kh�ǻ�EQ��m�R(G���{�e?��]�� ����^V��ih�A�x��2�Ds5Y�)�A$� /��NY�d������6���1��ud|bh6_���9eۓ���jՁP�v٘�r)�w��_�/ݛ5������ͭY�� m��ɒ^jQg_��Q�%Yl�N�r�,:�����#q3�oeOe�Z�o}��kkB���l"��F�NC��4�V��df:��#�[R�Q,_�^%�SR)	��v�? t���J���[��5��%N��p6>��lR�oce��x�\ؐѮ��o��ʩ�G�+3�j�<���	q=2�t���u���hwr2v���F�s�t�F�Gb���e�����<��=�
���C,�C~з���;;_5g]�o��5𒘲��4� �n�O9!I>j�|g?�����T�Vg����'�Ws�1]�Pڻ�a`��|�e4�>��<̴�m�.���X#�Rp�Z�v�Ev�>������8R�O����{[DZ�r��x�m~�{"�<��BZ��w����+v�5a+A���Z@s71����CFM�����-v�����IW��(���(aD�o}�0�do��U�a�g`��1���{��yA\���|�g2]q\R1I�B�8�G=b�T�E�f>׳������	���+��cB����s�!]N��&��27��ߦ�kQC=s�'�������[���W���o��e���M(> ��P�bt�<�	Z�Ry������>$�э���џ}ќy'qh�7���\f-r!H0���p�:�O}j2�6zk£�6<��(��0��@ Jyo�󧧔&g����?��M�\�T��������x�I���r=pZ��&7�@�1qmsI��{c����{lB#�:�1(W��G�_�F�YbS�h"�C�E� �u�@�ô�`w`��1��S4��������.��l+#�;oRB}s	63�����Q���m���"�<�߰�[�K�P��ȏ��%�&��̘(d���fL:�R��~�ϋ0s�osle���K�[?��5�Ml���p[�C�I�t�Q x������^TW� Hv����y��s��-qX��*]�YD[�y��3�od�Ł���j����Ű9�Z��r���v�P�. ��z���$������eIs�u�`��MgC빗��t~XqɸT2n���w��,Rĉ�1cﴩ[טP�Mj�*9э��_$Md��X�a:n�RA-�CMM��?Z�?�a��ω����z�+	���h�j��� mԍdy3vF����x=��_���TԪ�͎#1��.��a�#��
o6�W���>>㣂�T�e���L?�Ơ���]�/k(���֕��WѠU.H���m�s��Pz���D�	gc����,g���]� 
��T[����
�2��8��H��򶒺���wΦ��+Z��{&l���;U���M��+�yw-X�cix/3�U�)�5sf-�*a�ɺI�cZ�;�}��yF�(~�4�l��ph*�"��~-ye�K��3ԟ�hd���SQ��"Π�Z�d�~2r�#��ighz�gh�CQ4WSvLL�����j�RF��F�:�U����T�I�|ո���8�[�e�ե�d2SB�k��ŗ�9,�Y�4Z�(�f��k'�ڹ�M�Frp� c}�l��vf��h��5�C^X�H�̈�G�<��_G��b�}� ���q��(HH����YYa�ެ�Jz��V�����%|����E#��A1�&z����,/X\����T����;."�䭔�q|S���C�$�d�%��H,q��C�OQN;8���� ]�_���:�i�G�ɰ�����sSn�U�=��p�^+��zEb�ݴ�}�(�RvQ���!��.(��%�^v���N�9x��||O�R!���O�Z�yu����SĄ���k8�^������:_#����Yb�0�C]��W�m�	x_���D4�f^�z<<_���x�G�Yʗ�:��3.!�և��I�V8��umI1Qʒ�Y!�0x��k�D��<�&����(Ⱦ�V2��&�cW^��ɖ���=�&|�n'I��KĿ���#[�i0����$2��9L�*��󶣈!�}��J-uP�*!����T(V��^ϨI�fud%H��D%��?��1-���0�n9XQ����v�������YdG��m/�M���?��7�?��Ҟ�
���� M Ɛ�$(L^�����,��\X1]�3ɷ,$"D�c���v���髖����g�a)!f����l��yQ�v�>�9��(�b��v�%y
ptY����dc����H���+v�CR5e,9�����eT���F��g���'Oզ*�a*b�
�L�=K�*�b�w}o|��_E
sΒ�UU��r�n�-�:�6���π�F�y��M:h�.!t� �A��wv���1�*�D�v�P�\A�"�����1{w��v$GM�} .EƵs�����͗n����M$㻡�8����y� .T��虢9�j[�U����ǐ�* ��m�e��{�<��S4j���IK��NÚ�f�̛�M�� �ۊ�fX���M9��b˞��_��U�����^15��r�lB���,ccɦ�x�-��Ure�b�����gn�V���6����:���o_�!n�,�nS���aI�����Jp$H7�ھ��q�S�@``&�Uָ&ta"�J�_{:��I'��3�ޮ��!��4j/M�tVs�d-�ߘ��W�)�R���F�S�g��� rA(�68B���Y��UP6�yV3`a�u�+�B��4~g�O��L=6/�S̩.ZɓP�eN�?�-�`�Kp�`����\���u2�+�K)�c��&��Ãa���[�nJ�A�&�l�,��wL԰����Z7�I�^�Q=�\;;�N�L�<;����/{yd��O�^�ܧ"S퇌;���}���s�,�!8��~En��r��ɲ�iLm29����>�D�c�$볽#~����Oz�{�FQ�`�%)��i$诚wo���#T�@�0��6��|늻��\E��ѕW=Ӱ^{l_g���tجҾ_�� �̛�%�%0��F��&����iiì��Q9Wk^-%�9{����3'g0�7��w=��%N(~���>>M�!=�����5kX��u��Y$�;5,� �rU�gQ�9b�p4�r{�@l���>���!�oo��P)���e�r�I�i� K�z�"4����-L�<�Y�H�J�'�@2T�����sfG���Z��p�VDor|��r��e���➳��v�9��`��y~en}
y�Xx��B#��52&��o::I�}�����1�~�EU�"Pb�Z��y�䙵(�+��8!�)|�U�?Oz��"�x�y�u�C1?â���=[�|��K�����KR9�Ȍ���m�%T#z� �pL��?;�����L=>��ظ�Z��ߖĒS�|�Ӟ63�,�'Ø�� ���t.�-������cǍO*3�����F6W�E����)1=őY[��#`ѧ����;���{�^���:�u�����������̷#����M�i��G��rƣ���Z�>~����M�%LBH�ݠ�ц�Hі �\�2Hj^'��;��q˸�谎v��|�%N7�8�^Y1@$ܷ������o���<��$�F��ʪ��Q%C�c	�����W�*���K���I�2��W�����"�UT�Y�q������Tp��q�0O��M��Y��yȩ��G���\is�(uEN9m���ې���ilo!�& �dE`��n�s�Q�:2<��ƿE��F(����[�z������F��~�3��5X�,���*�:��S�;!BO�g�7Q�����Y͆��s��G��ý���0ʽ T�S�f����-:�fÂ>�P��@�mX�W#�c���!����{(��Q�;s�hrdC=+]FZ�rw���X��`4��K���W�v>5���a��=���/>!|17ՙݩޅD4k�g��u����\o�a�`m�%��d�ѭ�Px��>��l*͝N�����TA�����8T`
����H��6.>�.�Ќ"þɛꀯ`����
��k+�U�kMh]bf�8��_D;��CSW��Y��c��Ӣ9M��(�)fIӶÛ&���u�����w������|8��R� ��`3f��0�����X���b����{K�3�)�J\ sS�qC@����xo��c![ZG
��:(�����'��t��!g*sNj�.[�D�^1U�Ȭ}`A"�Qa����ۻi�=��o���S~�)���/ ����,��N�у�|��	�A��ms$�R����͎ʜ"Qv���Z�ޞc�	EA��n�%e`��^ƐU����m�#&�ȩ���tjܦ^ъ��.
�9nz���8�YxC���e�����.H��=��Ʀ����Gj�����}��tX���ߕmӦ��r��<�F0AB�4{0U�]��P!%�:AX�9��!����͢_���G:�t�D#�ǂ�
�o�����"�O+�e[���I�
��3v9��qܑ=Ssw����ń�AZ߀�s�ي�/��cx~�)���q�3���N��6�t��ui�����X5ZdMfȑD҉"��P�/t}	Ua����������7�:0�v�
�'5� �%���`� a`J�$�dQ���[�����]�[)5G�v?SfZ68�?�df�5�JZ�6�`;�H�#?�5���Y�*��G�-Y�I��8�4:��Ʃ�P<W�[^�7�� �иb^�ܪS`�"�����Pk:��eI����0�fҋ�*(�lNJ�I������%��$s?�0�T�=ߗ�U}T�)�Y1������<��o�{&��.
<S����2�S��@+�s���r�.��"m��Pl>˟v���j.J�����j�$H�9�I�%+�d`���u�kr��U�N��*9�+G�����Av�hk&���=�I�λ����^{L���-��C?5�a�쁃��,A��ے�X�%9*�כ&�����
�$2�߿�ff(,rÊ^�����/0��E�R �G2�9Z�0��	�l-��6�tQý����Hmڣ�ժ������r���}%�p�0�����.x�.�;2@Q����V�^6�C�<y1ʳr��%�Y� �K�*ƜWT���+��橱���>F�۰p�I(�ì&r�x�bg��3���Q��1�ZtL~Kx3E9�A<�i���������X�u��_(I�&���Z��˛j���=���ZR�y��r"�ڌ�2���`���;��W�U���4!�_��-�p&ݱ��/�E���&��S��Mt�:�gNc���b��>.]�i�n���U:T�sY��wK#��D�u�"�ȗph�1'�vI p=憿~�P�W{> ���Ahf��HS;*~�5��j�$;��6X��L�������ۥB��Y�I\�E�/`�&�`ۯ=���"��p���jeo]���x����ȇ�=<')��,&�Ҏ[|��o���!���U�Jng�(�Մۺ��H���Di�k�a?��a��*�\Ƃ3 �ᭇ9Y��MuM�"�蔶�/g�n�b��0����S(�&-�3�wp�-\�c>ڱ̬:�;���bɜ��AY�O���i�4��Z��_1�Sds,\�8[#q��Nt|2�V(��F�|�4/��89�U��B�H�^C����R�܇�s_ŎCz�է�JM�ߴ=�u�$�ς��L���<�l�p_�o\��,���ד���:w0[��g���ܕ�����>Mp�b�*�5[��޸+X���<@O:�ϵ���ʌG��B�U�6�k�/F�Ye�فsDp�{k6�\|��!og8�V�a�m,���6(�P������Ǵ�e�Ѹ��Wi6�k��A$����C`GtCk;�%#��r��4��8W��mC�+�a
`�.��� 9�*)H���*�p��t2t��L�˯"N�$�{}�Nw����hK���V��A�_ e_����4���S�K���;��ٿU;n��4�S�x�!գ�Qdb�
�׎���z���>�~NaiRbo�N����"t��JU����L�JӢJYZk�hly��V��p<R7\���;{��Ʈ��\��9�Y<�ވ���t��;���E{��)(FJ)eSwO$������Y�#���=Q�����x��,z����F� ���ㆂp�%�4v�&򧭓��Q4�[׶$�姟����d�#Z�@q	]�d�sՀOޣ�S�l��8�	�13��Xr��-��]���x0�a)Gwg�3ر�%��{<Ο-�A�b�h����������7 �@I��)��
Ń��f��H���TF,����%�wt^|�7�qc��ho�������ľt+�Å��s�I��f�E=���j؋�߁9�����;��~�.PY^�z�cm3{t�Y�n�gv#�x�����WI� ��фSs"N���Y)�=�}oea��٩άW�&F�\�2���n8�ȏ�{˝��7)c�u��Ra������*�@��G)#!G���6��fP������P!�hFm@��d��(�7�=L�A�>��[tb���|��������Qk��ĩhf��g���d�m<�0�e����-�Y��n���	s��5X����� �ڻ����8(fP����>H���V�]�ZB�Ɇn�H�!�|�ά�E�N�����޳,q��-xP7HږnQ� p&����Ϧ=�\�QDur���/���oup�>/�5������A��r�G�/ "�:�K��zh~���$��w�&¿ΙVH�a��k��ĉ�_��L�$�M����K*HE�	�{���#�Hm�∩��E�h�Kc�IIUqȂȫ�����_`"Ũ�϶9!ޝ�8 �?���J����K��>pݜ��PF쵄��矛��V�	C�|a�h�����u�����Xo����g�)u������2Ւ�C���H��T��u9�PFV��#�`�qnYE��2�a'�6�C�g�_!�oo���[P�Z����xO��9�GK��szw��f4�(ʻ����jti1{|P,y��`��!�2}o�D4�<�YS�	�V���.�P+��󮑑�|R�+ �7�b	���5l	�K�����4��_&BM���6���5E��3g�0���M��y����}�J���C����b�<"�6�i�	���h��^�	zt� �:�Y��^�'K��j�x�Jg~�����{	�ͳs���EB��������0���wA�Y���p��/�n��6���T��8y�e���ލ�t��7N���N��V8}���\�[��Ll#:�i�6��uۅt�ψ�B�o�!/Q��eȖy喦�+�p�.��(�.ϫ�=��$�PJ9D�B�T�JP����)���m�s���T�j��]F��QQ"f��;=��Ox"�"�3�ң�D�i�k��U�M�:�)'�\�2����^��K���H�OXZ�G���|*]�]��E��b�/?^J{0�QRV�V6n����#�v��	�MR����!���t���t�Ժ�+���i�OJj'u+˳
&��؉&�O��	�ϳ��F^-������aI኶��2�	�k���e
�d<��?��5�$�L���\{X=���i>!���wLM5��R
�#�y�\��ɧU��a-Z:H?ð�rD�I�P������坕NZ���"�h��\�~W�9%�@4��{(<|T��	w�.II���n�s_�	�f�%��k�ݒW@�)A���]%��~���MWU�ρ ���wf%�,��fB�д`�BwN���&}H��S|�*ϩ���wt���Bq�t�� �
�?��C