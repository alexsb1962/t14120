��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�յ�'�)���ҶtЅ�(�R4�K.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I+ĂiW,���D�+y[ف���rn��mo�����(����5���&<˴m�d
����]��;�I�����)O��Ξ4�"�\�� ���K�O�{��
2�D��7ީ��_c\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<2�q�U��k�8u[\E���@N1�w�0XL����[fe�Hs��9lSUQ�S��)���2Ee�Y�R2
�I.��	���
����k�������0�?�}4��ѕ�������U��=>bMab�	;4��G����a�����(�I�?g�f �H�Z��1]���%N
x��]Qu ���������	x]̍��;��V��
:/,-���	���Hߵg�4C$#;W���]w t��������SۣF߱�y�Zk���GT�U�{�OJ%
������7%OU�z�z.��e���L�Y&Q�\7�	��,�;���<)䟓�~������ЎG2`j��Um�!=�y����h�}�BK9�H��^$E_������b,�}�o?�M��;]�=��)�I��)܅���Sւ�~�T�2�bT]�܊KMb�w0�k�8���҆�|n�����|Hj`�~^T�ɴ��b��9J�Й�m�z\H�� 0��~����p�:�C��JS�Ȕ*Ĥf���J�D{g�P�r�|Aښt�  ",��9���1� c��(�U����	x]�<���e��8�t�~��,�O�W��s�!5�S��H���)��������ҥ{E�?HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ��Ny5�s�JFAa��Bzb;ym��+r��JʅqNA��d��1�:�Ω��
�/�r��]���P��`�.�D���J7"z��cX��ѬL�1m��+5z�P�_X�I�?g�f�L#����2=�l�����4�c��ҁO�����ߖ�g��o�4��?��d��q�G�+��T�����h�6ؖ� onc�����rYd�ea�;y� ����t����M���������b9����4�6�t�����\{F˯�+)��n̈́�zL͊�q���Vǃ���߼��� .�����ݞ��D	��U����	�I	"k�+��v��z�N������i��b9����:ߐ�؍��R��j�.(Wx*��|��p��h�d �'���Xw�f�VHF��>BH<M�z�]�!����M[��Ǣ����K? T�ҋX����>��l%i�-"K��^��Hm��S�)37J*u�������ݹ�0����['����?���F��ʙ@E>*;�¬pX��g��U-�e�,���6+��\�!wn�Ŕ"�����/Z鎬����
C��8q��f�kN�ı��XK��(�W�~:n=�ct�:��RE��W��_�ړ8���/��4��}�<��/�^�Ӭ����
L'���Xw s4S�'�i��`�z��4�+|'Tԕ���ߋI7��-5|>����n�xY�J��ev�mS��0�-����#u��Yk"1/���]���lh &�=p-iu�`���`�+N��?���&���#�{�0;�}����\Ҥ�Yk"1/���]���lR;�{m�B�5��k�:A�	S�r��AR1<�N�؆�B��W+`�x�o���{��&�e�5
��Ib����rs�i�jf� l�Ǜ������CyW�f�tR�wX�Հ��0@ȹWpH7���
I@1���t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s��.|Z���I7��-5|>����n����Øf}�
�?�Gs_�G�k�:A�	S�r��AR1<]Q�I����踫g(�r��!9nV�[}�@��L}�
�?� ��h�Ơ�k�:A�	S�r��AR1<]Q�I����踫g(�r��!9nV�[}�@��L}�
�?��`��׊��D�of�7���A3�(N��㎏qló��@d��שt�v��I�`2ڻ�ΪZ��| �Ɛ����n9�ycP��$m6��i�0�OgA�I�y�?ܔp�l
d�R�.��On��M��������4����/����DP֞ RS)$�i��Vh���*ܑe�W����n�4�{lGD�V�B�['����?���F��L� s�j8l������_ρ�OpD�of�7���A3�(N��㎏qló��@d��שt�v��I�`2ڻ�Ϊ�>�����!T��a���s��0�(�|2;$�JأͽgF"?�['����?���F����H�V�����,ycP��$m6����)�Y�{'%s=y镇 �H`|vXvs͋���P���L$y[)/�C?wm����ҳj �{��!���c�A�L'FC�v���]v1�_ُ�=�P{\� o~֊&w�R���yv4�����=b{ϡ,����x�-�)�$�Wdl��n��w�⽒���M��������qb	��G��W+��W�� �}�@.�:0�#}���{�sv}'W1�����Z�טy��j��k@��5��:7.SiB׀���!���c�A�L'0#P�O�D��QI2�*�ڃgڹ�E����W�6?���� c)�K�Q��ǺΕ�����-PE�9/�)����I��I��)���W�w��fDa>�Y��֕�*>*����8H��O%��<�*�AG�
�������?�d���&�(�6k�4d?��n��Y�10y��&7̷_��yC��S8�����ZK��Pq]��Z��~w�!:s��B� ��a�x�(�H�`��{�Q���l�,��3�L��B� ���vx!�읽��HN��R��?�d���&��A�bJ8��t����M~V��	��yO����w��fu��y�8{���@^�4���zȌ��t�h��W+��W���JĖ�Y�h�nџ�e��|�Y��ξ����LUG���E�����+T5�O�%E#P:�����φ��<�6�@a� ���N���Q'݀�=�յ[+8��H����Qw�c4~Nr_�mS8<�n�ݚ�Н�{k�h�+s3����b_X�XV�b�z'hۉ)��d�7�q�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�s�Yls��8��GM��-����!�`�(i3���_����]�C3����/�i4?$|�Ĉ��(a;��H7�: !�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rG߸��S�Ȍd�p�e�5�.�g3ZE��g�Hb��c�H�mݜ���,�ǰ;փ���wE�=p���Z�����p~z�r,:"�G�}��d���!i{k�h�+�/�i4?$|MF���y�|V��	��y�f�HYs����$ll���6�6����D5�|أͽgF"?�Q��ǺΕ������^�̷ؠJ��:�����@���Ձ�=�n�4��Ǳ߁R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#Pq�\E��0�}CE�>���L9��=>*J�X�$��,ZH��pC?wm��`q���9�z��,{v¿_.��45�I�{�P�՜���,�ǰ�������ݮ��&V��	��y�2B��$X|,�E_�CR��L(q_҂T�q�w���t�v��I�`2ڻ�Ϊ_��s�֙]�m4p`�Xp�T82g��	��#X�1���������s����Ac<�p{�5�O�%E#Pq�\E��0�`j3���Fm�b�vA`v@񴱝�P���Q�w�R���ykb>���pP�|x����.�g3Zdj�t��C���j��~��v;N��-2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hDj9�J?�H*�^ݙ����2������[he���Aɤ?ʺ~Qy��؄�����@rLj}^��6!:R�$l1T�n|s�)>���@}[Ǣ˩���.|�vA�VG��++��5�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc쩲
 se��rm���N�0`��:'����ֈ[�z�Ծ��!�`�(i3��0�C�D�Eyz?]4��jyP�����膗z��!�`�(i3�5,O�39�"<��5�{ �_�t�'�J�:}9e����8���y���q�9�}P�ux]Ѥi��}4�4/�q�Q�n����Sy8���W~��,���Q{�~D�T9w�[h�\��t�3Ah	)ޟ�I.��^�