��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�������*p�8������)���	Y�pI;&D�c��Ĥ��tc�)E�����0���X�Q���J0�wR���Q��E��!U�F�w�跤�/�⇰;5:�i��bZ�j�֠_��]�v��O���y�>�Yq�O��RC�ک�V�t|&qu���ݩ8�ug4b��hm�/�i�D����}�`�{���)�t:�/?@.�h:��*�R:
�y�NI{;[X����.�o[��HY�ї��{e[�2�~A�cW�PI�wC�LCݯ�k��n^�zti}INx��hA�W.�gIM�?~��{��47���}M�Z"��L�I� 3t�MBsZ�Ӹ��]���a�2�)�q"�P��� _m� �C�h�D��O�5�ʴ�r5O�~���5_mN�P�,�)Ɨ���e����~9���b���O�\�Z O�R���B���3j�A1W5����\�I>L��Z������D�j���Fu���0bQ�WR�@�(�f�N���y��W�5�mݾ}���0�%h)Z5B�DQ�E`L���Aq�Up?�q��h��VNk������,�?��q_�Ҽ%�3�S���i	pZCgS�4�`؀՞�@J���,8V��r�e�|��Y�Oj����Mo	�,��z�؇:6�(��{v6��
�=6��»m����
�Ǉ�B��D�#r'Yl
l~v��Yj�!�a��4?.g6�Y�>W��jG[n��P���8U��d���=VĊ����Hy-P�ʰ&�4�gv��q�%l���:��􂮜�	P���023��-��$5c}1���!��h͇��Jb�}G��kS�Y1K� �𼹪K��,
��:a&�kK�·����Q$"�:�z�V �θ�U{vݵ�ь{Y�C	{�g�����_�i�� U��n+����'&���bJ8)�9j���Hm�)�*^�����:{t�Ыx���3O�w�6���I��` ͷ�u+�[.}q5����j�� �I!A�ڗ�!�_L�Gim���ІI�!{��4T��|��A �r����tqO:䘻^D-�p���s���D<j����H���hf�	]�4�,��E��0�w?ܱ����	�Z���\M��	�ͺ�b7�S�!�Yꪡ����;��v����h�f��R�O԰���f3En�`Vk"!�:G}Qm��Sl�X$�9@���~�(66�u���O u}���ӱN�.�y딭��:�qP.K�v��栛�74���I�#������茊�C����Ö�8�@�`W�ɶ����ݩ\�_�����	s�����J[!�>��ҥsߣN���K�*4�G���5�����y���P�
������R��q;)$JA����ğУ�'�Q(�k+�2#�����5f���Ԃ�Z�o�;����J#Ճ�J0�$���JV*5����׊_��#K����Ni�c�	3�]`�V��XA�o�婁ôi�������'&��l�X�r��Ɣ�J-c������,���/�8�
o�^�4��C����o�����_��c��	y��2)�WiP.�u"��wY���,LAW=Ȱe��R�K�O��6�g�{貓�E�C�"-���� �Q���l�$��+Ef�H�#���{��s��3�������Y9�7�e���i���FGyd�nr���w��c<�sl�4��y
�&�;LQF�s�%@0�T�����K���hH<�O��C��ߎR���!�����L�����,�,Vk�7-2%�f�S�Hs��uOĕ�U�#�涻������e�ip,׻n����_O'R�> �+waK��ɻ������e<a�XD>)�F����K§!�Q{~C9�^D�	��+��T
��<� �(��q@a�}�A��\Z��Q�}����	i��f�^-]�"<�a�v�ea��}���y�+zV����5R=4Z��	N�q'�灝^�K4_3�$u�2q�k>�r�}�B/������+oՕ�i�{��_n��e�J�֠c�5�&nW���r᪪A�n	�%���{4��������!#�g/PԐt~���-�{7$)<�-�Ǳ}����U�QK�@�j��T�Ju-�YC 
��J�/D^�ͼ�%�3�bz3�Jh��!���G1i>�.T�*��U)�$��ڋ�Z_�k_����)�>Om�;V|k��Z9Q˒uM+tʴ�YO�ȅ�ULۓ&�.uC������d��yo�g8r~�W:���/ȳ�2�!�E�`�0Xﮄm�4�W�S����bo�1xg�y�SY=|t���q��8�����`p�P��$)���FF��w��
�����Uw����#�=2����r�فec���:'��.(�c�Jַ��Qi�R� Ei�x(��R,��6�74(�������/
7�Lu�B���q�������ȩ��\g�_屽EhYQ� ��U[䁃�������4e�Y��.��|F�����y0ۗBIO���>Db�@=3$���	*3���-�,
�c��4����#V�S�?(����7�UNR=�����T�J���m`V�+������<@���	a�{�Vm�Rhh�vj����Mݔ?�Հ$`�V�Ȇ��=��>�HO�Dw�I��ύ��T��i����U�VȡCe�n���C,�h���e!z���{�W��-�M�Q���C�$�u�_k�A[��ۦ�J�;����GVe���Q�V���:[3]w5�`y"h��S����ŗaqԗLL"Y	* �h;�|ά�^<9�TCG{�#O�Y��t7��y��g�uP`������7�s��L̈C�gs_$�hE�<����+�C�~��%Y���%OR��t8���SÖ5�}��K~��\��3K�����_6�ɡ�^IdD����)��^;Q��Y��X�fs�DF��p���,dFW�/+��@��VF�&�n�T���
�:����������&]�k�T��J��r0���*;I�X�tp�+n;��Aϑ6f1�t����`p}����i�*�Góp�^'�z�[:r��H�ϱ�^-�9=@O/D>�B	g��ְ��>�i=�#uaq�C�Q߭W|��6D`25����6+��x��g4�u�Xl��1���8)h��糢��TpB��۰!�&������^�a�ka��k��8��->n��}�^*�N9��s�b�)B�/�q�V�f�?Qr��ߟ/ii�8a��t잏\����`��\��ci!�	��l���~J%:b���NI�)�1r�n�ф�<�.����l֘��U��@!�1�Lgf��Z���'˛s�@�T���7�P��x�PiN��Ɇ��])>�U�v$������Y���8�b#� ����~W�4JKnj2$��X7eX�#�4���8"�FZXe*��w���Y6���cE������� D�=cl��q�IFgh��(&vOj�ů��<�5��M *j2n�,�0ס�F���w�ǳ`����lE4�f��U��*�h�U+�n���J�bT���������#�;��u(����_p�N������	w���_�1q���-�"h�W���^0��S��O���*2�����$Ã���ױ�n�j���S���I�Q@� �Xjڝ�J{?��d�64�:�2�3��cOL�����~e��~����ci�s�5�.С���MS-���tѬ��BʈF��4�͔^-����>m�\���ps��B�=^�U�$�UP�|_�m���ɰ �/r`	a��zxm�#����n:���F$kѤ�ېogF�x��)��U9��>8�$��)?,j?��~��IFo�.,�!'��W��]�(�E$��Z��:��`")��t���rM�zL6��SSdV��ڷ�Pk�%(�:f/�.˺{����s���8̩V�R��5������A��l��!z0s��L����,L��&�{�=Pn2^����!��6 yc�Q�����6��i� S��[�����C}��T�:�z	�h�e萐#�ھ����N~���ʼX�,־CXմ�)�����$��N�D)rN����/�O���]&�9��*�_N����W͈H��Ѧ��!�5�a�a��?Y�T)o�tǊd�͐��]�kh��J������+=����0������jW��6��H�:��.�P�.4ܬ#On�L�P�7�����3h���k+T7�gK��]bߨ<�-�!�.�ن�'2ߡ��l5��6�KL���?<�Zb�/pՉ{c�[JOr�U����٢��O��Fek����b��Ȟ�9��U.`�mm.�������9��nȤc
�@FA,�P���ߝ��f�N�-�\���܄L#fQ���vc !���U��I�!����ʏ,Y�)75��ݎ��nQ���Տ1ǺD���F�:/��CT�!�F>�o� �丄&v���������( T���T��;~%�;*�fb=b3~���F@�E�e	WR�.���\'Hɗ�M��Es����B�����
��V�FM@�rvZ��c�����������tb��İ!�y�h�^���˷�* s �eķn.�F�*Do\�=g��-ŖEW�督 �r��ge~x�̖ħ�	��4��3ۋ3Ey���Z+��7��4�ڗ��؆=I{l�����KΦ���zQ00	���=Q�������;�$ �5x�����k�*��6��a �y��0�@h/	4nrk�����x,'ey����������x&�AU]���n���a��������!��e�$�V�'�+)t<[�����}#�f�vw�X��+�h/���>��	��8o�	7kL�9ip�`�ѻ�m߶�q�
c�!@��W�*�:���5L�Z�%,Ź��҆�]�x�C�0ElVZ���(Q�����a�ė��p�3�c�pQ3�Ȥ�̆y��ȦH���M5'@����*1|3R5���UN�GUKbH�U�&+�>q��8�6$��[L���
BS�\��Op���S�C�S�b��QG\=�#�0(�<�����N'�zEv1k��=���#�7��^�F����(�-�T����\s�5��;[ �)��[WE{a
#ㅢg:�yKk��k{N1��v(�?��hf�1��{mcdw�΀Y�s��O$�� +���J/.�Ä�1J?װ�:w�M7�IBB]��d9���
َ����Kը�B��]^�$Z2�"��d���D29�bb[��Sj�8�5��u��3BDU��B�Կ��g-������[ ��-�(4�;�8f�E�+�d�Z�9X�;���~��/o�L<�V/�l�Ԋ�=/y#����P�L�_�01TkR�����Gf�pM�6���_�M�<wt�N���D*�~1vx�hK�M��kS�h7�k
�RΏ����;�4>��Lr�c%&�@��i@�Rv� 
�kl�?!���#��z�'��Zp�y@w����	nڝ4UfY������Y�����K2g�I5�v���=r�V�Jk�Q���Q�x!��C�
��ZXG^(�r�iڭ���f��0i��@��[	�o�
�i[���W�fc�!��7��P �mU�N�R� M�ܓ��ŊyP�?�rOw�t��&wkZ@;k�Wq�6�U*�E��s����\+a��ʰQƜ���#v�ӎ�b�@o�.z+�[�����_o�
�"�9{� �P�#��q ���!D�A�χG��R�<�Gi�[`�G�{e���~a�G�*g
{�n]cz"ci��sp*ze���E�:*����s��-�&�B������I�1zD����{�|�tT���7ۂ����G��U���1�X�]lo=����/�2=��y�GqA0r�-??%�T���i��R���P$n����lA$zq��833���|}9�Т*�j!�$2x�(0�`6~W���A]z�WL�����!����f\����Vj4�*��#�Q��sQ�`H�S�(�Z��T���4���/��[����{R��j��W<N/��|�+��C>�����������}��n툙��*;��:�8����҃o~X�	$`��G�S���Y¨�ۯ\10��%���������Z$�ls����/vCr�� ��~E��FC�Ⱥ!"{���,L�����,��vʎm��
�|�}�� ˘�$�0�~���?�`�X��C���A���# !��
\H�}EP>��z�*̸��{z�fg\��׷�E��`�c����J����V�<ox͆�G�y�oOf^:����uܖ�� ��OL�4V>J��t�i�j��5Ʃ��;vt5�C���K�����[����S��_����N��k�ZiiQ粕M1;·��N�Ic|O�,Qb���SQ�I�\�ٷ%@r!L�ԯ�gZz��|eOP�dw�<�$�մ�{1�/�������V���?��>����Ɇ�T�j�;��e+�-������~�C�z$��Rz�k�UR��2mNzI�
g�a�����'QI9��8�q�\ݽ����d��"[��X�2��kN������#�ٶ���@�0�+M;�2J����l����Ut���G��
��^����x��)�������R}�,~o��h��,d��KC�%���S
'�/�����8�}/����g�V-��-L`��)a�߸n�N3rȧ~ҽ��<!��(>>S�	��������L�`[�i�"Zo��˛���eO�dFe�V��t���
d��I�ئp�u�`�������`N������@ߔ�d]s̳C�2�����$L�|q����m�!jz��w�A�Of�N�j��u� :� ��
)S/��~��џv���}��OZo+ɇ�M8 ul��*+��c	<j'����\�Oͦσ�4Ti7�/�a�E����:7yq0�(��#��$�" 0Mo�����-�ҕX����Ϊ,9ZO援<Q�-sX���h#�����t_r�/�z��6ڸ��:��g�"�yx.lĚU@F�j>����?�92���`��N���˜�h�G���ަ��m�<X����>�C�I1�D�(�������DY��C��c�ᢍ=�315�q�ˁ��(��>�A;���"��?�߮���8	���J5k�VN�k�؏(���!��� p��4�3kF;������e�X�{)é��]�)���W�b&�J�9�Z������������6sj�P���m�a����ϯh�ꕈ�,ȶ�o-P�g���xS��zF���?s�.w	v�BD��hw��5�U�|4԰�#��b����
c8�SOp��a�_ N�Dܕ�5c!�O�mi�JQry��5�Ӈ+J|� �J����
	��NI.�ݼ���l��ֈ�<�;l��G�T����6X8�"���"j��ۭ��R�v�Q�Q�@]�*ⅻw�t�P	������4�2���8PKs�M�)Z�V�=��Q��ޏ��]����H���|���5/z�0���/	�S)�f�HzQRnF�����Y�C���Ho�䗥�$��f�������M�������M��h�x2����Ƹ*�,i�M-�E�I-��b�(�ۻ"$��\Й�?�AVQ̐�X�g�"5u���'��'����d�,|^u�Ly렋�PM���j���ʲ3��~�h#T��E������q�F:��=����|�,5��Z�ݘ���G������*-��qy)�N��j�t���,��[,�����AC�P�-�����V�sZ���#!N]6�]�1
�����$�؁�2��y\��z%��e
�Ǝ�dƹ1���J#io��d�ȹ`��d������?���,:1��(�]�ǣ��i�v?⨒ �ZX��&��>�[�icR��	���P���j
��Op�/�C��FP��
%����F�c!|DtڻkPw7�{�ȯ����R�}Io�Q���2��]�����yz޺��a<�7>��Q�h�d����?gQݝ"�@��ĉ[T��YjS��7�{���\�*�|������l)�����T�σ��6�vL�kglL�<'����SLY�h�'�[{�6��X��S��(r}*��p�,�?�^���Ր.+�{Ҹ�>�7>C�I������o
gO4���7��w�zV�KM�N�E<�� �Um=Yk�v��pɜ�D��뺈u��zrD�p���h�v�_�+�Y�X;����fz�(��O��[=ƨwi~P��x�mn�V��M.�q�_��ӳZ�CYLJbD�"P�|���­��VԧY��M���o�&m_�?
q�[�[$jt�e�V� �L�7��G��1~t5Z�f�ō�.�24��kN��$��������~�|7�$To��t��S��wL���T�ٸ�ŶD-I"��ه9��R�������t�8����M!�k�7@��5V�B/'�]1��1��`;�s�7;L1���"d!��T�a>��Q�)�r���%�$�`m����pk��'!Pk���iOv*+P�H�w�[3|���ܼ�I���OZ;dj2{K������9�ș��*��^��L��CL�x{"��3�VwȂS�vD�S��d��q�i��	C�f��F�h E,к�n�8�_�b;����cx�.y��-e-��h��w�y�����U�,e�q�<���-��G˴��ۍ+�Ȗ/�)��XQ��:B� �\���QUv�Zz4&2�<HKR�~��b�Jռ�,�*�g��6�8�t�pMY}%����C����<4��Z�ͷ�X�qԣ���$ѿ"�"b���	d�%�䍲�Ӈ*"L�����f2�-z]!�&��5�P�:�sN��ݚ/�c�p���j��>��&�Q�6��8���5�5�=����K���!G�0*�]����^�
��b�Q�a+����d�J��ߺ���uE�P�Bl�+�T$��){�ip[x��@�e�$SI���\�6�����b�Y��bC�Z�G�% 0ӌB�[9�:X�/ȂJN6ܪR~��a��Hc<�qP�x��'�F�+�~�	��Mw��G���C�Kn!ň�ϸ0�Ɏ��+���n��j��T�'Pvq�b�.��$�l�;D�6�r�d����ȡs]��1���\l�O'I�!Xij��������ߨu�쯲:��mb/����	�֕|g��q�X��%�$3n��x��Π�g�T�9��PI���=Aj}x��,�<^�:���U�X৩xZ] ����ܳ�������*���g�gf��TK�ax��oP
<�Ӗ�CoBK���p�j��O�����l����@��lK�J�����{V4~j�E���_�.��͊�����"�fv�m�u�`,���3�.r4��~�x����PdbHt/K�Y.KB�)�p�'k��W�E3D��f�C�x{��֓�6q�:,�KAܑ9�h���嬚���YP�E�Zݦ�|y=r�Bnw���߱����H΢[ѵ�S�w��,&5�����{��-|do�E&�6()*�F�EٸP��>/T�����(�V�8WB�e���!>*%�Fƍk�K<5�q��;�.��!I���o���������\sӉ�u]&�RzvO���1>�;:&�����4��|�uRe~�rI��VQ�݉Q(c�s�fV��������wl*d���sV[�L52{ʍS��_	�n#�}�P.F�g?�Y'�L�u 쀱��DV�
0�?A�Ɔ5�"R�p��?6#S��	^p���N=����"� ����<x���biES�~
��᝺�,s^-�)��dYf2e����*�"~y5�����\�˛v�1�ґr!6�jwn��E���b�[Fb%%�JM�s�M:���Us�����]�f� ;�����_�C��\C,��4<��p�mM��(�͓sr=��~�[}�/���gh�r��r�8�R<>wCź���[��]$����2����;x��l�]��4�r��`I%tn9 �Y��0�]/��)��@���_d]~��\#�[<=rA��j��v��Z-c�ڥK�Eu>N-*�C��װ7��-��D)���ɚ���&�Z�&aͅ7<϶4�Ȼp�X�.2l{�7�	�r�PT����E�1�������+l[������W�r<aŵ^�&
�ܫU"��eL�",���O�還%�$~b,e�Ĝw?5��t�l�!��T9o��(-���'��75]�)���T��6
I�F�w�QF��[��9^u�&����X�C�J���O�SRuՅ*�d�xF� �C%���iO�����Χ
~	H6�@�uS�؇�>��!��7QW1zv����	��$��J�̬�/ɉ�rB������iK�d��@_��whR��#��|�����k�m��CFm�k��Q{oKnb[�h�3����,�P#�����[��2k�1I;ּBַr��nZ���iup��ԵIKԷ��HP_rK�᩵ng�ŉs�	��[�pT��U��0���gj�ɻ��:T����Q��U	"���V��N}/'��u�/L�lI�x�)�g�
�LeeZ��Vo�)«^�q���H�����)�}������{�Y�|�Y#��sl���([B��&���F�}���3�:�.��z�_� <��QZ���hG��>���T�Fٕ�٦�9��F[�}�Y��4.�r��:���b�=Q-x�{�篆T�]��p�5�l�`��)ѕ��loNM|W�a��~T_��K�o��KC�ZP8��:�N��ĥ�y���=���\��aϾ��!�b��q�D��6r�_�����Eâ���i�:�tt���]Xs�����R�E�+��w��e�%ˑ�b�/��Ȁ�j��3�d@��#�Qss�$�M�����q4_������qS�0�D'��#��
;N����dS����pV���x�@Q^��m~�k�a��;�D���#`6&���I�!���h�d菞r��O<2��<�_���ݘS��j�\�`yL:�x��#y��
D��S�'�����4V�u�����P�"ydB��*k�>��i���-V�V�O��ųv���I��
4�o�\���ug�䤤�M�$,�S�K2݋]}�>�3��߱����&r.���Cnm�}5n�(������ i-;V,j����T�.c7�32�؄35J�A�4�"_�*8����V��!��[��Y��a��sx9�;_�F�6)��NǼTɄ��f�~R\�{��H��q3�I!���"گ*�gߑ�'|�l�+���o$�'�c�Yߩ��`*d�~uƀ�U�d~�t���F+A���<�C��V{���ޕU��-:����T�G�z4���gM$}S��, ��NV,��u�����0���_H�nh�t��f��[_��m�oP�`��(^�|��&E��X�]y�.Q���� "A��J��[�Qگȴ�\|4���]��<M��9̶�.7x;DoTn�B�c�uefh�~6�|HS�z.�Z�V���<߉G��gJ"�-R�|0� 5��$�(���S)���&������~,�j���	cE\����UG���>��&R.��\%��D~��)����d�V?�����VF\��
�d��z?�DboGo�+�	N�_(���􇅑�҆V)l������"�Jg��,^wT�$y��`K'7����s�,� �L��:#9���fP� W�%�
�e4��|Z��,@�T$�����\b�`(�Ϛ܏�])�~��i����@��Ns�M�̿K>ѧ���n�41����q^Wh��MgV��#P�����Gt��#o;0��J��MVpJHF���<����N�
���ʩ,��E|�3��j:��Q����mL�6�^��^Ǉ��1[����1�)�X#4�#�q��M�P�O���'�����^ܷg�g��s.P>����P;��d{<W�?=���#���"�P]���ԫ��0��ǉ)śr�T>�y\GH�?���2�5e�y�&�����Ax�a�#�8�e���=�{�]l#C���#�=����Ȑ�"ܱT3����i��X�X�xjڶ�T��a&^���������P�KÊ��I%MY�g_:���UЂ�J���I�t����1�J,�ژy�ckn�3)df�����W\�]�'���kw�¡�Vǆ�h�1&�*};+�M!X��2Z�('S���,�;��y�\���K��@�u�P�:�]fJ���MD
w��e�@�"�������A���S�-L�����`�{N��	&f���|r�c?�]?l�\h�Ԏ8nr�e�i�G`�ҋף��1��ڶyL)�Pz���#���?�=�̭�R��b T'��ǿϝ��'��J����T�6P��S�����]*����?����|W%�iI��[�t���Ƙ�����#��HR����������v>g�P�,3��h����[/ ��db�8�#u
�6!�[�K��+>���.���a�D�bS�:�:�ry��"��[]��3��6)`�W0�h#�����Pm����X��o��l���c�`Ks�ӹܨ�l��	!�Is�p��sM1!�I/3�`q�v�T��E�ӳ��P|ʮ�dBM�r����`���?��R��Y�:�����a@�~\�
mn��=�"c��e4w/-Q�M��|�+l�I~�<cA&��=\(:TzR޳nf򗫹��ς�֌e�5����;�敳st��
Z"����
3=�0J;x+�'�s `(:�I�K�z7F<[d�YӜ���nɖq�ak	��.6~���C��g;>�V��ɩ�p3���MV�ҽX��È������p)뢊br�>QDH��F뒀@"�]GC�wa������������#���^�� a��Gbl�+�4�]�Pi�=�1�m�@$��I�i^�'dMq�@,~Z��d��� �Oԁ�?p����!�SY%E��Xgp�:ϴ� Me
	yK���=��M���T/�{I���c�R�kW��t���#� �^&*����>e�0ɋ���m�b^��H$��Z��(n��D聇|'�W�}L>(:����!�Rkb�,i�X�������"�K��w�m̶�����?���}^�\^�=����Zۭ���b�����VD�I�+�:[����%RU��h�A�dm�d�̙5�ʞ=��U�_�)�n��k�l�#ol���V���XB{;� �_�� �Ճ:�yRD�ȗ`�z�b+8�ɪs����t�����C����G���9~�_��t01³�$Ȟ�%]� �5K�e�l62J��9hYUiHt���9�Ğ67�Q�>�>����Hd/�aa?w����m���<|��m8��������$�1�EQEX"p�!�g�j��my��t���Z����5�9���h��3\��uR��.��zj'�/����o�aZ��f*z��;�P�%����R��9��Y���]�cp�/��#��h�)��v`T�?l���W�!,mP�1s!�s~��!��iȮ�����,�߼v�'"N}�m퇔Ŵ����b���I���t`�@�v�Q)���$Sbn���j-W��z�~-/hӄ�I�<Y�|��Y���z'�E��(�<飼6l�9�>�Y;�A]A��!�2��6�
��͂}f@9����(b��p����O�'-�J+oR��>T�����E�Y�
jnTɚ����Y��Tc�`O�3�	YR���tE^[C�$���Uh��8�A�A/~�o�P��g��G{�x���n��IG�9؜疼���駱���ڻ�|��o���45[�5�G*�k�K��x-���isfH �P��4"f
#���5�~��{�`f�}c�i�m^��Sw�����a'"IAOc4�D-G��bpi�^�c�ٰ}#e�J՘Ұ~��P�w�0���'�������`�z�0M��
�aH�>F��:�ۑ�i}���D갾�
�Em���4k=2���T����^�����<�����k����c#�Ew��F�f�0e��⓷p1D��9ꢑX�Ճ�1�wŢ��y�� ��LO5M���C82��C;c��`��`J�<��s2�=�{��5�T]��~0H�����������y���4��.����;L~�����H�&W��6�+��@��=\�l��L}?�/�;.�82)��.n6D|��ڞ�h
��<��w,4^��N t'G��K�d{9fD}�Sl;�c�����b+�� �J�Y`�
u�ZC�,�����d9;)��J["��<�uX�Ȭl�+�k�/&Qds&;!��#+�n������z���:KU��/m$ω���[�ݥ,鶭��"�`��H�5�v��(\�/�����4$*K�/l�����w<YҔB
������[�:�s����L4��j����q^ke��o�qW˫C6���C���g׈2�fY��%�ͼӼ3{�<��a���nײ�C��H����[7ʥ^<�Z����J8��ժ�O�ҁ���sbe:������x��������T�OP�hͿ����z�'ѨU#�mKh05��Y����H�]�4����[�=�M�_�L�ٙ]q݉�Mg�r�4<I�����*2	V2e��ƥ�u"��RI���E��	�16�o�Q���i���i�4ҥ)'g���D���q!�G�]&Ҥ_+v��<�W��ޥ�`e7m-��P��kI�>CQӊ剳ޣ�CR����i�<��J��8�࠯�g�2��T�ѱXx�j�ȅVSzI+�D���]�5�h�3�ּ��l-gZ��Gb9C�A�{A�m�$D��62�T^�pg�}�^Q;M��#'vx�.�I���K����'_�`�67���b�M�>�^��+�����@Ч�r�� �A'`�ְ/�BYma:d���Y��ۓ�A*�v�0���P��<4�w�ܥ�"�D�$N����߷�$�X��H�]�xgˎ��Ab���nMF�d{��3�K��5����{�+��"x��Z��7�\5'�#y����~��ӛ�G+�O��(w���`}������)�����_LU�a& h���[1�J8�º���k��0	��|��� ��0g	�^y��]f��	����}}C'�]�F)�P�����E�$��=m㓔������A(R�ҋ�O�R`�7�<#�j�MeQ(����\Y�a��*s�ȑs�l�>2���V���Xsw_�QMy����Uu`U��q��cQ��[��( � �]�J~�
BWL�R.��}q�\0a�}����mc7�����
,����pu��	v��r&0����A������5f�q��55�<��!U9cƟ�t	4�?z����4ŧ�qѽ�f�K\�)�PmûĽD�)0r^jc�<��R ������%�ePhܒX�a~���c:y&���r��[����% ��U��We��XS���Ɉ��5*wyvU��
��_g�A��9w�`F��;�vŕC�Vk2���p����!���j�F��1Tdς��":�o��4�G��#��`z;n}�LSq�l�M�td���c��A��p���h��1,e��z{�ou�Ɩ�-�����14&��V�ĔJ+��W��'̸珶����!�6Q\)�) ������=�j�!�UP$��¦�& ��������q�������o�)ˑR��G��֛���B�2V�C���G�k��!C'm���0o��Yh|?wtm�h˵����Q���u��xB��x�W�/��H2<�<V̍�oQ�Ӄ��D]g��ʕ���8��y��o�p�l`R	@B������ħx�7ԇ�gc����f�p�Q��@�lQ�T#��"��&�T^����;>������R#�JKς��3b^V]��8SUԉg�i�x�K.kJu5��DV��%�����vkb���e���`F����uXc�XBf����[�Fj����si�ث�^�j'���ªaŞ� �l�t���%�Ϫ����h�9�f�{�w��n�*&��ӗ��D�~L�K&b�a��K��e�l,,��κ�����|�NJ5X"K_��k&��SZC�n�>n"�X/�eEH�X7�P�M`rmH�[z 0Y���ι>�����v��72��Yx�N�~���t	��:�'W5��~Vc�%Cep �e��ƞM�Y�w����0�6b��$�Ѩ MǂT�,��&9ԅ�_����k;�Q��Ԣse��Z[V@m��m�^� |�y#(�q\`fX�+�u�.�����r��8�ܧvĘ�rr�su�ZujlTϣP�� w�+�}���kP	/�`�vy��W�&�)��������bg+m�'��/jӠ��X�]�ǰ�G�},(���lG���V"9��UM�Qn�m?9�|�C��Ħ�b���O(�[i&Gb�+�?]���P�vcN�t�-!>����Y����+&)E�D1;==�+�ba�U�q��Øm�/�M
>���<��^퀖>Y2��7�,d0���v�v��Tv����(%G)= � Y�^�/T����@/��-3��U�o�j���]��7����+T� K��L�יY����������KNKǂ��eؔ@� �E�-��O�z�6ʪN�8V��K<?�nIT��4��`���7�O��f�v�zY�;�����K��ܙ��i�y�I� �l`��'�z�?�<hy�˔zƋ�6����a�)apEr����f��W9��W��#��o\x�5�VQ�����C�a:�]~��,�O��Ou��V�4s�0ĴS�;ǬTZ�2bs�	�m��撎i9h�d�]n��_qg��q�p$-�.{%������n�0��y��+[�y��v��8��c�0��ivދ-��j��A#ud�aa���<w�%���s��L�+�BFAg�̯=�
4@q&�s|�n��'�ZÚx\�Knb���d�1;Zf7�is�ϩ
<��{�ig�^L��9�_gtY�"�ϡ��ϓ������ؕ{�oV�By4��D/��se~�}:-��c�p�sN�<�£�x��PI���� ���g
BHe�HZ��F�"Z3%wA��9�P �J-B~p"����.��'�x���mk�ӛ
�IͿ�\��C��"���@mE����6� � �{�m�Gg��j���1%Yf��УϜ�kYf�ժ��'z�Я�����^c�4�Ek[�0� ��dQ
�v[����>��E<�G����!�Z�����M���ַ{�x������WR��1M�Z��~,t�Γ�{�LŠ���WJ�E�c��[ɪ��C�S�qq�]��B�P%��v�_�PCN��ܦ��%3��o�G̜��7=�gS�;"�+����OgQH�s�\�`S�j��>M��+I�i��t�͒^�=�Ẹ����ߝ�c��Q��N��tW���	"��I���3���w r��3���Y�(��y�z
��7+��;RM��N�S�U������fBe�HV�s��7��� oݩMf�_lI���� w���y%Zd���������j�:/�1�Qx
�a3NPF���X`�Kh C��n�G׿"��}ϵ���D$�l��3���ٍ��LC\����ŭç�u��G:?�(�x<f��TF�o��$�<��i݆Z�=���cǝ|���@� .�wa��>�:,�d9Rq{Fi������GU��:��O,|܆c*2��ٸ`)���@nX�]7�r1�`��5H��7&T6H'{��2�J{�R �rB'<1���x���oHj`�A����G��OM�� ,�FI�1�А-�$�>KܠѺ�3&��|r���s"��~�p�Y��qde_V}=�fcÊ��Me�O��fZ{�6|�ڐ� �zJ��*�SeT���g؝a|�ه�]WË���QF?jRӣ��!�2�W�r�7�Tԥk9���4�T��!����ƈ>2g��sb��qR~&>CP1�A��CK��R	}r�f�{R�w��Ur�T��uOTH�1�Sy;���#Ì�h|��-*ӝ����I���d5�g���B�\�]�>�~�t&gaTiگ�j��Ry
������pE��U{� %]�U[H7�a��(��=�Ģ Q���C,+b]�~�n/�bD�����d0�x��#~�Ṋ+����3T�\�~�����R�4�õ�졛�z_y&!��e�}�j �1c��/���{b�X~�����Q�!��o@5�j�^f�*�
�VQa��������Y�C�JRt��A,9��3��4b���!���_����������5I<nB��<G��>y����hgV넢�v���,[V9(���ꀋe�'XvT	IN�s���N��w�}r��c�=w�k�/��e���}Ua�\�=���"F��B�A+�U��\�C�\����Ӏ��f��R@c6�f(]-��H��A-s�u�������-�@Vk�Bp��,������p1+q��R�s�L�q���w�w�*�n�[}8�X<�ECq��L�uyϮ�:��$��	���G��l��Œ��.k��27Z�eʚg���B�('e�\.�����`)J~��_���b_��<���4C|A�Ի��[���Â^�9������J���(��pM�a��:��8��)���	�Dv��Nu�O����F��l�] �c��1K�#%��q��I�^�P��y��y��ɶ��h:8���G�V��r��p���Q�0 <���6�[�׺L�`u8��-��ͣ���&p�DE�hnDvY6��Wj��,F�����+��ŏ�H7�@�Ś��Z�&-�p�/��:yX��C���N���S|�B��2e @���QE=�{��<���h�H���kª)��aF�s����^D\�C�>������
5[C�<��'��t��5P�����!%B����ߪ�&��>��"6!�ܯ?T�`�g������U��V5�xW����7�(>��:`2���~��H�1�:�[-���t3װS)Y1�l��%���S.�s<����d2��f�|I��D�)���h<`�������yu���Y����U���Ss��&j�O����c�ъ�x� e��m�+(�{ ���^��7 M�0nMM(�"�)�&�L7�o��B�#ql������t,��F�U!����i�Iv���x����ɚX[�h��'=� �PDSD�җ�WC��s�X��O*5��
~#p�ۂSb�ҽ�h{�u�GB��@*Bw��ؗY�b�Яln-���Ezk�c�|x3 [ I ���B��b��k���ֻ�%b��jx2�$�eY��Tf:}���������0�j$RWQZyȇ�ӁC ��Um��d3D,.��	�.Þ��4�B3�dO��UA��(ck��SՈ1�Ȗ�ͩ��ʰ��BL�y�ù!�/W�j)c
C9��ِW���;uF#s��s��&Fʗ�0k����v=7=��LŢ�5���;φ���@E��ל��w�I�.z�6�ް����8���^;�kS�m������:_��;W_�%�ع�<^��x�\��F�� "�-u�C�b������`z(�������#��t\p�(Z§]���Z���\&��痲�"���lv9C�t#a��QX���G�"R~�<);d�p��M�ң?#P�q�*uA������[T�n��}�ewh0�I�J(�B�n��2q����Gv�@Ï�e0�*�«��C��M*�m�_X�k�VPi,�Dd����>��>�Cr@�������L�x}� �o����Xbyb��:c�)���;0�~��'t@�����Q�y��E5�4��rѾ��C
��b.�H�8���,���y˙F>:�O��2�� ����ڪ_i&�����.ѯ�I9��_7p0�1S�C"C�M��u����ǵݨaݗ��`6g� ��v�i,�"&�Î��rn8�B���p�Ӹ�QX�|q��$qvR,��I% ��;�+�} +�Ȏ,z�,J&���C%�_]�l���+� |��:�T
�A��r��/l�W��zDN��5cЏ�Qx�����~�>����.% @Ky���Ýv��[�T>M|�Uwm�lUruDQ8OJ�NT���=x�a����@	�պ�Jy>������/�u�sm/M�J$�y
�'J^��*�1|����m䊃UD.�Yuo���ɪ��B
:D�v'����he����t~�����I,�PJC�[�~���1d�j��e�<q�n�d�r
�g_Ѩb@<��ƽ:k<y?�����#��0���*P���f��6���� ��2�,���0s�v�� �w�SjP 2I��� ��%��k��?�_# �]w�29���b���u�#��BB,:�H��x����\ j
H����񍋦��OrDW~	}ϺT��?�8�4�S�D��(��<�w�PWⲶ́�<��z���V���L%ukp����G���\��Ch(�� �n������E� hhP!����������#���d�w�A���G6�
+�U�b����2�>��Y�s�P$ƢW.Z[4�����+C��숣n�(pz�F����*rh���w���#F�왲\ތ������ߥ�Q#\�5�Bf]�_�V_����h`@s��"!�2��$�%C�o��ޜN�#ukn<�*�6,U���H�w��o���c�`[��9�>�Ф��}�2
�FA;����P�R�G�� �U�*��s&`,Ʊ[v��6W(r����{�;?Í:�B����
���b�M�T�d�|]u.���F�XUf�����5�:�n<2}D��/Tz�(3��X3�=)��c��gK�y���S��yG�ּ�س�K��#������%�<@��0�Q�⋊��(Od�l�+����1�殉����)>��KD;�@
�u����D(>�+N3��!�&2�#Ly� �V׆X��2�~��A+��Kf���[tZ6�h���/�	�N��~�=ltJb�Z�*N���BC�(�#�^b	�]������ ^ ���¯��n�x zr�)���;�ipĐ�=���B��b��8%Gj��(���s�L���`���
!�v��ީ&dbUE��+����y�����@���V���6"�#����i�/\�e`7k��`SO܊vXueloC�-G;�;�����ژ8����߾�^�;P�yv�e�-gl��������':����=���~�-D���57��i���U���	����BGA��@QG�V:ʨ<�uh�ξfcJa;.�-w,��[ԻpN5_:���]>�"fh�S~��HR�����L!ff���"�O5�6�ms#����Ll�r�i��Dk�x�x^^y�-!<���%�&$L0A��Z�嬷�zL�S|�T�
�w!�e*8�ĸ��ɲ�xbq/Q�}��i:�X��$.��`�֍`�±f�J:*3��L�QtmoV�(���U�{+@���E.�u6FY�6�Z��rZ���WI�@�1�@6y���Q"Jt��m�������m�3� �� cϢ��_#g�_��mش�(�߇���1�;�1Q�
L�43��3z������Ԁ�ms�G��K�NH�h �d�o�'R�F���>L�� Y�M1�:঺��i��b���͂\�p�5d7�:U�7���bї�z��H���	O�@=j*k�/
�Ɓ4\|7��刡�(NQI�"�j{�-���K�KY��L�����v�V�U�o-e* �۝Ð�Hb�P�VJ�3���İLV�m��&C��ZB��N�+/���P���/��e�g��O�o��j����e6m~�C�= P��  ��%�kEG�i��D�T�[?�:��ԣ�'���S#�2����X=�H�No�˦xuM��s���cn�Z��
�!i�kR:ϳtÈƁXꋖ�o,~::�ˬ_a���2>��f0n5WX\�����"����_��mP	A��E��kE�D!�	���HM���� cӋSp��)���u���>_�P��j2}��RzP�H�Uh%��|e�q ���Y,�A@'�ѿ�m�`g��^�pZ�ˏ�_�K�f��8D�j3�Z��\�!m� ��u�g�G��*�1�{�U��q[IHMK�\�m��NQ�2��6��_b�m��mƑ٠c�� ��fyWB���Ԯ�<Jߣ� ���H�y$]|_C�SP��A�-dhiSˮ`��F7��ʔ`"��Д�O��c��� ����k�k>�D=��J$`�<�q��w'+X�/�w��v}�O~�c�
>�$�W��Y�~���ɊK=�o��!*{��=6'��<�|�J�}A��3��M����������}0,��"y��n�/`P"u*Q�b�ni�����@��8�S�Z6iq-��#�{�	��F��D�#	i���<|d�t��ECp���y����M1�Ѝh�p��Omc���y!}m��O�C�š�]�D� G�O���Gy���;��%ze7�Y���l�(���(\��s�y�i����S��,=���44Ez쳋�Ѹ'.�b�V��y��z&�����u[~:P�ʸ�7�C�9ı�t���v�noB�NP�G� Gb��$9�#xIZrCP�z�9����p�"ȅ6m�~�J*P���?����<�X�`;�u���gEz%@��*Ҩ.�l�TՇO1�R�6�,��o�c�^��/� ��Dz4������!j/�0��tZ�7jߔ��e|󭂻�ї�Ԫ��Pɲ���Ey��B�b�G��D��:/7���j���m���W�LC��Eqۈ'?����SH�/��mi�(��}���u�����*�F��rK�%�i���e���3yq>T�@����\.FWn#E8�9rUnU��q���p�ֿ�쳓Q6�f�L%�s�N�R��=��\Ǧ7aА"���q>W�1Ϛ{!��kY#�����)�I��e~kU�8��
�_�A�V�P}�_w��FN�E��Z�M�+��]@��6b�Y�3(e���4h�L�1.et�6���/��[����È� �}t�W�p��Q���Q���5
�L9��q\��SY�Y�ʧ������5�,�7�l�l,~V6)�N�E����}l�J#ӷ 3R�\)��U�����x�?(��Հ�7�w����0c
��~�Ӱ΍����4I�����q����b�2r�X���S��|��5�r�dդ�]��#G��fE� �\�ֲ/_��"hUD�����I�Lk��K�f��S)h� ���.�t9���uT;52�
c|��y�
��-���;�J�*#����M��D{1I���I�TѮ����J��6K��fH���|D���0#��̹&�-H��_=]`�h_�l.&�T����*y��5��l�Ra�V� �g�r,Т%��g@�)BB!Խ�uXB�ՈX��]��"�SgAf���%m�W6�2�5���vB�6�B�vh_I�U`4c;��_��\���� ,zރy�7}<lq�k�!Q�G@���������[ۊ�s��q�p�(Bw)׉T�}��_ڐ���H��;Ȍ��,� ,�x�����P>��5��R<�k���D?��c���L�q3������Q�0?\��� ]Z��A%�:Z@��>3�.��:ݽ{�L{H�gexT�rV�O	�Sm4D������>�oո'����(������g��B֡�n����Dw�2l����(_�A��ϰ�(Z�e�&XX���G.n�=���j���;�=w�cI���E�E��x�v���YX���q�kx�$�f�ŸxK�Z�����1҂��+m=F��@/M�&H�������C/ |���LP:�u�Sx����D0�<�G��_��HyU�6o�f��C"��ۍI���ClL�2�����o�2�7&?@x8�y7��oG����h�y*��l��m����=!�G�gX�ʄcJ�
>�t��>s�zz� t��LR �`����FI_d|��Bu�L�?���
�#Nǵΰf̥S�#�utk$ .�	o�9�+�P���q�R�m�Z�{��H��C~�Q�����.G�n|��Q����ݓ�\�K?K��Q�ݓ��u��x�=�}�"6��QG��hݷ1���<U��r�Iʱ�3$��P��Ob���+�n��D`�Y�%�zm�.��T0�(���L �r5��u��	el4
�
,y1+M���<V��� ��ɛfL��=��$�4��ËoeE��Y���'Y���R���P2����=���x0��/�Ȃw^\����ְ��B�T>� X�<�42�#1����ȏ�����>���c|��4暯�}�I[�Jo� �~�����@��!wr�8��v�I�~�c���%�i���_68\� 5�ߐ���M�Ѳ/(�[�	�����&�A�	'/�w魝; ���d]��7?���QK�T��d*+A�$S��M_�K�=�Dwd��I�Ā�&W��2�5���<��˷�����9w�,L�-��N��*�1 �ÄE;��ڸ���fe y�9}x��[�BӇ� �|��7ckg�Zb��!l97�7�-7�i,LT��������k0����U��1�(j(=�f�X@��z��&���qV�gDbׂ�H�����NЫ�*}〪ת�I�l��~�� C�z@��'< &���A(#+˼����	�����a3�{��[��DخI�)�],#��N�lԈJ%`�9p�:f�Vͳ ���e�������n �8����c�Ԋ7�W����\Y����
�l*�vԞ]���Qb�*�D��t���mi3`(�ȯ���۶�r��mp��� >l��6�ސ�^�Yè�>���˚&�V8���kuf���g�Fs	0!g��TPZOA���ݥ�V4���V� Bن=��T����x����5iݛu{ ���D���`&s���y��(`�]��*�ߗ[��W�>��E���3���u�*�b1`bht��Y-��~*{��?�M�΂�9.:���E}1�XE��v�o?r��v_vВ|�l5o���)3'\]	�3�X��Q��	�{1�� ��N"Aij�x|�hƌY<�B�C���2 ��0�HP-Әk��1w���|��:c��C|$vJ|�n6���kZ��x)"R�Z�#u�
�HֽT4�7)n.�*5J�Y�4B^gB�O���\������(vL�:  d�e��q�	�Y��`���!ȝ|O#D����S���E�;��VY�F0�-�=Ò����q	B^(Ŕ�?��*����,	���oc���z��q��nm�pr��$��)�c��J�'`���(�e,ЪM�=��U�1���C!��NC�GB_�B��n�(��ީ��];��H�cH�\��;�+���wq����r��L]�0o�"�Z�2̶��j�QO AH���ZaL�&�78�DV��&��Z��]�2�����TץZa�A%�բ���S�O>��	�m�5{�����*��E�3�����z�F�n	�5�o���<�8�Pd�~o�_6������8ҧ$P�O$v�kU����-|�#�Y�n�:h�;�mrՁ��e���-�a�n@N���b�s3)&6lr�WdmK>[Tȏ����V��2��&��&�V�N�f׶��55I�NQO|����U!���!��9��t`�Rg�u�O�Q����U+
Yh#���u���z��$�3%�ɚ�IP��I�����	S�?����ў�ю1����k�
b�=[}�I�sp��ov��2SZ��l���	[M���2�����I�5�(ru�C�a_ϓ-��{�����"���s�C�ķ0�JA����.ha�h�f7�Ω��nXs.��!��O���t�V0�o�9��8�9�]O <y��[G7o��Ԍ�r�!e�qRe���#�l�>���T�0�bd�v�7������{�D���Z�k;�GC)m��X��"��+}:M��o���#7J
�¬�KD�f��s��������'l6`��
��=t��������2��
�k#�?����$���m���Q5Ȉ�A������G��r�M2s�z�_���)[��;�M����X6��X��7��8?��@�����
T�h�_pm�@>�^N8�?�Bv|j�2N��.c]M�rKU�{S�n'����*����,����QgVqaʓ',&��;.�]!լ�����8�)*{7�Χ�F�uL�),�sW��X���/����c����u�2;��V���DFyÓG}[�-^v
Ο>:}�T0�#�y�e�l�onF�,AO���BC�<Y������{�֨Q�E���� onPr���`�?I����k�'d��v*S��N���U�nB�$@�M"�`7�դ���IٲS�?���N����%b�J�W�ź�r�Un{59q� ��lq��֠x�f��xD��|T`�ɶ 
���mՁU]�Tj;t���2qC �[�Um�IP$�ވ?�1d��c�';|�+uo��ءp2]N�V?����9�DsE��"�FTV?pJ�x:�w��Ś�+ɇx*輕 ��7��_:=�3'��ה|���Z��Qr6[�)�h�jP�t���5����E
��4L"V:z�󴠱a�
j�C$�4��[�c��=<t��a�=�Ȗ�N)�au~gT�ߋQ�~��ug��p �R#(A�W���>+��S�zHe�)B7y��pW�t�a�UCe@F�<ۯ�c
��U!�5�e:�L^� �W&A������n�=���[Q��3��	��X��>/V�I�ڳ��Q'Ts{������} � A���`�@�LU��N�O;�;=�z@��j�'��*q������~��t� Z���ˁ�ң�p����	2�������DX�����٫��4�1�戥����XK�?Y=$ۓ�!�"������N�_��%�g��M%���K�K9ο�G!�K�d�4x���k"�b���p6&5D=u����9
!F�zI~�({闒Փ����{V�ս��-� �G�W�4��$�%�$�R� 3��W{�I��X`�"�YDğo�(��5U���qٍ��u�[�����@�Nۉ�����U4�q��^Q��~��:��l쮯�Hx;djT�R�QR7����i��۲@}��B�ح�+�>�~y`��-�h����;�b��N}F�(���*��� +"|��{����[���������7w-c
H��W���
�.�&�hk�����o����OO�:�e��NK&)k�����	����{���UdN��-��H �G�Ã��̔�Q�m����ɺ�\ �M��Gn����j�d=�,h�5�xRtL�����
vXgo�FUj����m�k����cdN�v@���OY��T˗�Aj�ϳ��2�:��!��y��T�Q�	S�@�yb��w��hۛ�|RO�9ͥ`as���L�S�w�#��<��?�P=>]{�&�HlL�$a�(�JJ��A��Yk��~���\2�Z$	#r��?�̫Xu,9��B�??C4_lIhk��"�?�@9�\�[ ��z��w��!�{���<�Q�V����t�H-�aAT2��
���C�gK����Safjo4!�?KΣ vb���vR5����;�����/BcHP�. ��f�n�f�� p�%Q�cz��̛z�u<;��y��n��Foǳ?�͘WQ�ǝ�F�� Jz!>�a�:�AdC|��i���|�#��Oa;�Ђ	����?�3���3]�m�x�u���ld�EQk�=  Q�D�Ku3z-�0��T�����I9>W�x1r
����e-V'qYP��ݞ��RnaK٪�C^jk(;����UxYdU����6f���YL8�[ �͑�����0�&�Þ���f�� č��N]h���{E�оY�:�%� ���yXv��kңv�*
�$�,>���2�3Ź렡�$���U���� /�=ܤ�jk�S��iBlj��7@Cy䝋%3J����T/\��M.��S���+�4""ʩO8����բ璗�j��[tkEI44�`�r 7������A�kwXL5g�y-�Μ;9.dA�����hE�x0���0����A���\ڢ������bm,M%���pX�j�y��g�"�d���T5S�n��q��E@<�ݛy��-S@����)�h4��Õcb�wJt!6M�|!��J�\��,B��'���a�A��L5��k{@ú.�p��/�1��◣ړ	�l��(��T�-�e+x1yO�b�=����������[iO����ƪ0v3��9������������D��|���D���7�gu��X��Ў�F:�X.�E�Fw��Γ헣`R�����Da��nIm��ÂfoI���Qr�΂���^*���T3�<�Qoe�}�ø�Yt��ɜ��/�Mw� s�*�E~,�ޖ�#2!c.*I]��bH�j��Ŕe�+:�Y���zG-Mwe�{)�_�A����8d��L�n�$4��͡�G8-�8����}���z�g<TQ�3a�qd�����B'W��Tr,�J�3w����ya�k��Zᔣ#%��g����Y���~��/�"_�!�:Ͻ�o��"���v�b醡�.2��
��	��U\�ba�������W���9�v����3<��D���q���}BV.��C0D/0�7����rvVsV�ԮCf��/�lF1����{mV�Gm���8,! 2<"O����\=�m2V�J�рz� E�"M��[`�1��Ф2��UУ����I�!��q�f�ϑj��bbh����M��g��D�>̀^80�A�-��z��/�����*i���!�^���3e]��}��ο`\܆�z|�S������`:�Ő� e����T�|�Yy�i�}��A{��ݔ�K��zTFt�<�r-�Y(�{+oLk&{�V�0.��Ż,e��Pk;�w&	�U�b1�P"��ʕ����&�`�f�@�/�k���M���VG�m�|$2���6.#ɓ�`SE���{�utn�jտ��˪hD&���^�����h}�8�筚�zȽ��v�V!�+�Ʒ[߄ߋ��zW~���ݮ�<.��ֺ1�~��[�ZR�&��O�g�~F�+�NNWb�,'y����x���d�����hT���4�O��o�26�2q��TQtԩj	��}G� P�;䙻r/t�5z�J:�)�r7��ٞG�S�3g���f|����~s�yYX1�w��e����:���h׶c�m��y��w
���5�sSj]��3@G��\��%"o\�b��(�|�z6_H�9R�!4�����j|�L���߰v�1��1 � 5��4�m�!
S��A3g���~�cKw�yO��u&2���>8S��zv�_�ך��O��a��}�y��J
�����tt��r\`���v����h��2"R1�o"��'�nگ���s5B�\���x���D�����\�e�=��ϏDކ���R��*��"�;Z-9���R�Q�ρ�#�nV�;,^ I�-	 �Ԡ_��F�֜���3g��2<,QU��c��`���g�rY�ꑷ�͋WR���Yy�տZ��(3I�1@��/�Ȁr ֍wv&Gt�c��~wD��p}�em�񀕈F/�"N�c��z8�G{�f��^�HZ���qf�~�{?����7V� ��b6QĤ�N3oj4�Al��k��V�X�P�۟�΄>63�CT������	R�Ρ|����"Z�:� �%����B-p��l��Q�]���| ��ƕ��촡��'_mQ,(�W�w_�su*��T�S�E�J�;�7���ۖ�3Q�t}a&���t�]���#ư 6��2�%���J���७ɸa�I ����v&�$�������1���F��;�F�����������G�~G\W�i����T���>���8�C���(J&��������u�ċ��J�A�tbP�nJ|�#q��Se��Вc���<�U���;be���n�.[�K@�?�_d����Eѳ�Y���'�	A�x��![uq{���,�>F�� Ɛ���ť���'�t�'j�vHTBCS��1O�xzO�@�}��^�H��_���a ��J�3��BËo��:�Hh��2�SnL!���ʪ�v�KnA�\�ю���I|K��,�����^l�'�K C��ͯʑw�˨?�am͔��6�,�?4��mQ�^�" �����Wġo6�$���;�m��4�	��C[/-"h����lUB�6rIaŧk����?d��Џ8ME����E��S�E����H&ƤsV��8�-�A|v�_ǘ�/)�8fEv�ܠ�N:s1�<��,�3v��(�S^��~p�ɭ�q-������F���pл1p_�V=��p�D�A�hD����<���M�<_gq-i�m(І�}Fv�:9G�j.�9~[q�~��C:b�>��s	<�^!�v��� ��&`Z/�����t�.��Qˏ��]�j�S� ����kܕ�]����JvUĀ�b��cͭ�B~E�37�2��PH�(�9�`��io�
l�&���������������$N�7�6�yI��mw�\����������3Crjk�B`�|���\sv�oO�Z�@S@�cs��9�ѫ�d��UF�@ht\�a��Ap?���,�ؙ��4�L|���f~Dt��4[�j�-Ԭ�M�
�F)n�� �zӚ�rr8��#�e�ϰ2>�m�|�h�p���B9��^�v�����.���헉{��0��i�Q}C�۸��~�~d7�'�.�%6G4-A�+C�I��O���ZvJ�CA��<��?�е�Pr3���t���Θ�����g�C}�{ԈI8�:r/�����ݶ����Z�0Jq'HVg����/�������[W��2��[�����֧ �f0��m����U�.�~ly�s�V)��u�� ed�-��T�^k<��Ħ���v;G/V����S\k��>�֥PB�W����B�^�[d&X��ʓ�-%D�0@j�sf���
�21��
�܋{y�W�p��ee� ����t�|��A"��D�涻�Ez!U�<���܀d��k�P�u� �L����Mz�^&r����#�i�U��ƕ(���mL�݉�M��%��Ǘ�H�T�y�c�rS�J�Q�OX q�ǡ`s�&�A����֫6bo��<L�'`c�X�Gk�F������n'f��6�	�jш �d��g�F�k�a��h$�j��?��&s�Ō�˽H8�Q�־��aϮ>�T�l:��o��fI7�nk�����f(W�/;�,�L��d�&��3�kRu��;k��n����'�/<H�������;&����j�.D&M�K�y�Ks�בp�ֈ���K�7=[�эH�)�Ō�Ҏ���j�j�=�0zB��9����/���T%]vp �,��y�t��Sݜ��KD�����&��M�eI���?v�����\����Q��ӥI�+�i�y@|�`����g�I�w\�g�қf�IS��SR��+���s�a�nΗ.�7�u,��|=�k�"���Hc�非=1������6�-y/n�h�\�y��x(&|.6�u_k�+l�%.��}�����q����1-x�:}t�b��g(��J�S4W�,}'�'�y�˙gSm��]�R�v�*��s\��$$
�X�H��AbL�UKƔzj�A���<�����@Z|��6)�At߼�X��h�ɝFMW�H��y>AO�p��\f����*}P�=����K�jUBA(E�P�uNt�6��^#%�*�<pG
''����������+P�u����1�&'����Kl�l���@$�hb����;��l��,����`���K�'���9[ٜ�mX���8�H.\�\���W����<�f<��+n�|~m�����M����Q؇W�l�������^v�.H�2��:^M�7���>�()Y)O]�3?��x�]�r5�������JV�Kl_������<e�vm�R
8Ĩ���l���	$č�塲�^�v�+��k1��༽�&߀�P��!�&���(?�XWޢ��j�9����z��z_��Q��D�u�<w�&�$&���z�Z�p��4� �o|�W�,.���?&+z�����W��cy�ww����H�-C`(���XǏ�ޥ��hV���7���<�����`�Uʬ�%
�w��xTK%ڧ>��AA<��T���ix�ܩ�h��ǥ�&��V�a]��ώ�A�aH?�x�Ƅ|wY^�h2�t�n]\���}���U�;Q�(�t�� �+�p�?��)����&