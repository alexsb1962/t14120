��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����rC'�[�7e���5%	��Ά�ZY`X���D���#�I�^��қ��
���4�e�4igȩM�O�´�3�]=pr8{��7�׺�ĵ/n��pϺ��/����?�}�����{�ܝ'a�|��F�c%1��_�U�"����e�ehxs�f��76���|�ˍ�,�.�pz�����J�m�B��(2��ko5"�e@%�
/������1���x�E��bqB��rW�����9o���s�"�3��<���-	��ϵ��d�,K�_����rz9�)��}]���V��bxtO%��@K��_
�kgIsw��@#7�+9�YY>���V�D���*��%I��B�s���3�[3���=U��=4�\�Zo��	+/�yQb+%�����n�v�J�;@�������DXfr���L��@�0眹�m�]�0��vʍjG*�t�jY�LV?h�=L�:�4���Np��=����υ���j�m� �@4SH!T���u�o�?�h�d��>�@�-�t�Cv�͈!h|M*RDg=��ցh8������c^����v�ߜ�v?�s�˭$H2.|�P�|7��!�j�;m� -Wb���
@�Y2��@YB�_��k/9͘��_"j�+5�N&���RV�>�l*����5�S�+'\�o���d9�G/���,;5�������a�.SY�A�:4I�����{�[șk� ��(-7
3S���<����YѵI7���u}��ox:TĊ���!�W�A�qZ(��t �%�`��V��K[+k�*��:�N�N��������t��m�p��ˬ�Ř�N� 0o������>��+��_j�l���U$>��6qm�&�H2OK�D��4�h���/�]*/����mf/sW+��[[�k�Z��G�$%��i.�5"ӶT��gx*�ܵ�	�Ͷ���@�.�.�S�OG�>��7L\���^�8��ی[
��=9r; gز∨߄8<����Jn��P>���~�M(�m�Fs7����ٛ0�;��[<TkJg�e���5����[��E��S��f����N {a���ȡ�{�_��g8�uᅯ�$lk���jp�8/�&�s|����M*�1��0&�X�'E�nsm��b���̮Xq7�=�+�p��Zjr_���"Jԗ\6B����|�M��J7�#��Ȃ5�+<�sk�31�9�7��)~�廄}�O�	)/ԧ��Q1�;VB��-1u�0S�q��@V{�o�Gz��Md�����C�Z���i9�*�t���b��N�ςK�t7��jE�I�U�B��f����v�ã�D���E���+������(ܐN��4��6�&YZ/�L"թ��)�&nO/��}Ztmx����L�F~]�V�G��ԓ������ZJ �Т[� ��ҏp�2R��r���|#!%��� ����C����²�a��z��.%k!��<�/%?�=����MNW?r� �8�+��#d�t1BO�/����ݽ��2U���g����ߔ�@3Њ�-^4=�@K��1,�R'K�M�:�nj�Z߱�k��~R��ʆ���P�:�o1i��C���.��k*�f��ʘu�1�QK���i���	xH4�.�Ib�p����X�C�F)����!p(w �0�j߁߁6$15���~�zj2h�'-5l��%;Km"D�-��Z�X
�{��2��G��LvK���7��ٺ�h�#02q������I����Y��g(7��<���"w �)��lPH8�`�2>f�f�ޡK�<���PYi��3��	[�S�6�}��F��A�U¹?y������e���φ:'����,���/�M#�Lh-݁��W)��ʉ�w2�ϫ]1���ʘ��P�E'��U�2���e�-6��,j��c1�mˉk\�cA�Ci"����O��~;t��3	��jF3gV��9;��N&W���9���WTEۜ�'֨s�F�e	�����w�%*{��Z�B/�`n�C�V�.��k��O>R���H-%��Ꮔ��
]��1g������y0 ���.��C�M���L]�uT� �J�ol���|����9���� b-љh�>���h��`�8~�q4�u��\����5?>�ٱ(,Wc�L+"$b��V�N��]���SȹH�I��x��J��]{��(U��Ǩ��Р�������`;J��Rvo�f!M&�J�R�O���{0L�y��"��T�&L���2U��s :C��j��p)_�aг%9Pcb�)JT���F�p�u�CM]��M�Uy�e5�:+U��KO��o�uB�����{5�8�m��@�LS*�㑃=&#纐�����/�'l��ñ��KOZ$��7��f� jji��]��Z����|UhS<þ=��`w����hЗs_��`:�Ɯ�7�Y��Y��*Vr�ŤWC�|���6Z��@�`C�Ҹn���q��a�W�qܱ�t�3��E���#�6W�*��>a�`�����
ݢ3g}sc+r�k����~�>"�2m'- ��o݃:�r��c,+ܕ0w���y���@X���p%_�k]��Ic寿)9��y��_5��Y���2�+�F�ۂF�$c��[?���(d5�;� �tp�;g+��,1#�6��l.�*�5�{L�8�ڱ#����ۅ���н��*���2K,���Qr�C��Pƶ�c���G�t�!2BE�0�qܣ�J�Q$�L}|�9��_z8�b�Y"Zn�e E������ێ�5y���t0=~C�3B�ݲ�$��l����ZA_��mM�j>��a�k���Y�4M��6�͞/uS��v?�&a�������(�)Ջ�ۥ�X]~���󄹞8���N�����|��e��)@���MJ�Gx��5�����+Ǚ�&��E=�&k
�I��%��|.Q��2�v���ed�p%m²NUS���l|��6�U� ݕ�d1U��=6Ϯj�k��u�?��
�[���'�$�E?��n�%�������s�4:�H,D�-A(܆<��͞f�]��� |4׺TLL���G���/C?�+9l��j�n���ظ����<iv�U=�1H��u���Ɣ�طp~H��W�Zɶ����p���Qcb�S/v����9Jt�w ����:	��erw�#�Pг�m�i��ˠ!~�V��8jrM�^�hS�([R�K���B�N�@�x
}���άem�CPz *����mʮ��Z0ץDN+$z����Gʏ�3�*J�dA򼫾�ro�Dk�Z�[kj�V��	�w/�X#2b�|�î�\ A���{������ّ��&@+/F��?ظS4V��)��P���!zXr���XB>�`�Ը(-���I���Wg幷����,7_�z�Fs�<�<k�=6�⨆��"vR����Ĳ��U�#x��~�o���ef8R�e��]ӪH�3q�Z��8m>�z�5#�q%���;��Z�`���~Z����0Vҧj�a	�9�bS��Q����:"��=��ǚ�2c/��і+ٰ`��U�`̎�Q*��7���LzK�m�'k��9��t�a�6��u�j�\�����@�	��3�@ry�>%�����p$.�y�U��V�[_�U�>��}|��y�ٙ(��؅���i����ϳ"�q�_��\��2�˺U)PJc��h�1���D#���	Tf2���z�]�����CJ-��7�u���ƴ��?{1P��z���cd<�൳�Y4�0�p��Q9 W5$� 'I�������\)G��7+U��t��~�t�b��'��p��X���w8�o[��g��:��6w�w�����q��"��T��iw�5�x�VqtS�<����������vu,���� p��%�ʥ(�_�T��M��0�R�a	��v%�nPWD
NJ�������$+:mN�'����IX��s�[�$
[�Kw?� �@�x�	��k��N������(��U�j��In���=�������Ӻb"����7�� �^�h�L�9��?���ڦ���QnΝmٓ;M��3	�b݀W�x�yk��0*���y��}Bf8�U�������>y����q�I��n��i+	b+�����!���5g��:��4:� �t�Ρ�k��JyHf�]�2�d��i�*"oGW�Q~$��`0r��	�k�t�--���Q��G���@as^O*�f�W��s"ĉ�u���7��>~�oF�}�^ERz�0H mu�� �}f�>��;6�_��K�q3��0XD!�[�.�S��p�
r	��� ���&s�l>�KAf�J�b�r��R�(���
3O�OA�t�|Z�lw�\�C<�}#3��Av>c�)ϯ�޽�8�֟\u(S��ڃ �8�v�A3��ߣ���C�J�����ۊ����E�N�h�8;F��)�k�SVɪ��W�v(�����T|�[�=�<��䘓���������P(,�0V�+/"5��Yr\LIF��[�&@$�R�[����j�Bw�̈́�?\c߅hN*걆���s�W�ϟ�k�P���8R�r����SN�5U��e�UQ�' �������~u
s����+y8����A p�+{wþ)�g !*2�ս�P�t���30㡬`��5��Μ<���EUB���\��O=$O��EK�Y�$*�"!�m��o̘�������_��%��Vŀj����N�j|Rݹ$�%�+����-����2�e&���$�KID!�Ѯ)��cqRr�A��tWp��ƠR_�D��o52�F	W�`��gXf� '�S\�|ꂂ���R�W
��w���5?��B󌶗+_}�N<�%i55�tf��$���{g�$O*.o5\�����0T-�]�ڪ�<��B���]^-c(U�-�tS��I	��;�c�\e@���&O�=�1$ilq��<��!}�P��7&�+u���A�;���!(`44���<�2��)�U^s�6��7�;�a��wZx�h�YkҲ�N�-��d�`'w�#�������xA�Cjpi4
R�]�S0�`�ab| Y��./!�h	��X�{I�=|����������D�U�����1���H���"[=Ș�B恾����� �5%Y�^�чg�I1l�OhRΥc��A�Y�����	�R�Ty# �&;�z�A����Ol��������q��θ�Ӈ���c��q����7�O%&��eCf�ۿ���kM��k��HsǄ�sߏE��u��+v>��I0M�����܂��B�ٗ���d^T5�%��!����t~�:�NcŽ��T@��;}�v����k�y���qo�F|�Lɺ�l��5��J�&�`�O�[��XzorP6������h]�h䅀��r��خ�f�ˣ�~�j���p�^H ő�0cl,�]"�Oda$z������&�� �(�.��%��z���{k+��[���3ڦ�����MB�G���8��Ln�xDt�+;z[��av���P�W�z�=��꿒�rwkD�$MQ�@��xG'��э��$��6]W<�̩B]��ި�3��J 4)��S��(B��;k��5�W�_�<z���5���:u٧�>~}dө-u0l��;���Ln��t����������� 1F��go�ް�K\��"����pJû9Js��͡�]<L\D�O���#7<��v�2�GEV�������ϜX=P���[��	aG���X����H��V���+@d��4��2�l���dC�����n�gۭ٫�I�edBؠ�|�;_�i�-9��� @w��/-:���<	��G��"��[l?+�:�{�N|�r0{�a9C������>f;�ؠ���ZO4��h2��+����)�@ƚ��ӆ00D�4D�zgX���v2���e�4�e�\6u�(�E��z;��%%���=�eD�a�]ļH���?>,kNTI�c���\� >V�zPh	�F��w�Hl����-6&��+���a?��p����x-3{,����_z�Lv���Qĺ_,�-.���R��H/�9\�Dr�a��"-QcjQEC:}`Ti2=f���q�*�(3m�Z��姐�1;ٗ��-v{T��ݼ��{�"�b��xBG���)��?H^*�2�hT~���Ԇ��-3];ٻ�y��h�2�D(q�d�2�MK+�J�L[�|���=p=.3��7��q�sy�^��|�4E:b��u}
%A�:��ƕ����.�ri.����7��<^i-�]1��6s����DO�_-��w��j���@u��;?o8�q���C
2n�8�<��5�U<���Ku���~��];�A�K(+jj�U��54��� R���p�^�e9���_��a���h��
�ŤI~E��ȗ%
��B���z@k6�+�<���Nc���!֓�G��cµߺ��n����x.{�����5u�f���>��U�aU.��j�)�7Z_�N��[�T.a���M\���ƟO� �Y�$z��������q`4�i�.�Q���o��zW��2�����)9�ߵpi����֢�:���D���q�2�Vӓ��(��x�t�V��o;|�&�|��-L��̾/C5�!O^��M������X*U��Z��cn옭.y���0g��2���M���2s��M�VO}o�ʢ-r�"�oy��mW-���G�5��ː3���CE�����W���քLp��I�"���#�x��ar�M�s�X��y���ӿ�7���?�	Ir�c�]I�6`>G7=��!b����Y8�x��ǡ��*�8�ߥ�\�!�!���qHu?_�;���HZ��I��P�=_�E��K}�y���ՠV�,�N�1=/9����w� �P��t�?D��
����v߾0�؄����}&P�R��{�$(�S *톣Agܵ�E�)-�w|���Y���=%�<@���U�̀�Ӭ|�H�F�ND\"A�]�$ �{9<��z���-�8�@M�� ���u��B���u�����BS�ʂ]'Ѵ��;�e�Q��l��V�@�?l9�I���
 +qf�P��"T��^C���YZ����\������pt�|V��=�z٣��R�~��_ |�x��a�R��x���@$�صL"��9�3��a�T���Ƃ��Fk�L	�pJE�Y����G�+��`+�(�a�y���>F_ac�Q���`g��ި�9��#6-���U0m�ո<]�DX�N���!Kq���GV	txz@�7���z���m;=^�/�X�nnr��d %év�ٿ�ݴ�5� �  �j�!	�s]u��:+8!�q9�T h��u+���;ȶ#���(r��8��ӱpr#���'����z0m��Z���8늋�NY�'�q�u|��]NO��nA�5p�V>�z�s`�s������B��	1=JC�2� ���򸤧O ة�@��Ą�i9\),�u��3��߁�e�w�@Я�9��%���H۰允Ӝ)qb,%��5� ����Q�j��C;�іmV���VG1�-��-��އW��l�����+'C�α��j�)�Z� ��xD~O�Ȓ���ߓ�|Y�ۖ�{w��С�u-o�oP��5l���γ�܉n;IHz��x�� ;[T*jt"�a���"_&�(�Ǩ'c}!t#RF�-6\ެN����h���l�{�ɸ+W2U��>������F_	��H~von��þ����޴#Q�P)Z����p����+e��� �T�]@�V�3n��$�*2����Gy	��>��?��~�R�Ě
�O�
��� ؋�n����կ�=�{�㋥ "n}�XG��\ma1�S�F�s�� ����y@���~|�zj�㲾����WFI�HѦ���38�tI!�6�ԙ���M�Lm,HT�C�@[ T�1Ȭ�JU��Cv���j?�X�z��Kf�`�$\�=����
���&���_㥈+]%�X=��ӳ�75S������s�6�>�J4tWU2���0�����5��vn��O����^��g�f_*�~y���"�:P�"|�ɹ%3B�xz{�O?��6}Lt�e�&!�޹%� �v�l���C�1��>ZN8L]p �w���ទ�_T���T#cNKC2y�J��op��}2UO4TJv+1����;�������mW��F
�t��ɘ�cp8�J��BN����l/0���0Ch��:)G�n�E� ��z��c	߆:% Cv��H��DG|�c�H?f�,;0 �(�\i�)]*�<q���:f	gϫ+R�F���Y���DP���w��DA����y,�� �y���?sXӮV<O_���}I��>Z�ѻGZHq	�G��)WG#w@u	e��X|!��/���Ɖ�
%SH���GH}E2(���S�������Q��؍c"%���`��Z���Ⱦ��f`��PW���@�])9ֈ&��H��:Y�MT�(}Ge�$o{�E=��p�L��N�ܭjX'�i�������k8Qc_(}e`����w-$!q h�բ�� T�~v�o�`R�Ēnt�ҚSͷ�s�_��}�d;�fr@QGR�K;�0gWS��cd,�B�Z5=�TuY�`NP�1w��g�Pݑ$Q�7�z$���I���#��5Jtxg���uz[�5�OI=��t�V�\Y����|żn�����|%܌;6^��r�[^MG�H���� �����X�7�k�"H^��{!x%��v@j�ާe��j%ߴ���.�x�ޞ�ҧ㍍��~u��1|��
H.@4��G*f�>mDb�d.��X'�B�e��y��?"�!�Z�R��1v�bQ�9U��&��"f��:2ȡBU"�� u��� ��=Wxd�F2�&Xh�#(�@�����/=@�h۫ʕXz��阞�[�r}ϛ�Gs3H�-Rm�ai�%W��	�)�B��msU쬳���ɄO<�Je�ZE]����y��Oݒ̷�z|m�I���K��&�S�N�MW��s�i,�3�p}��kIy��L�Z�l����{���[V7:b�i�� �12�b�k]�xx���_rý��R�E����ߒ�.#Ύ���96,-6f��n@���V
��A�hBS`�W��Ŏu����zt��t�'wQ������}_����w}���RW��v+/�����`u��ޏ�B��3��᫷7�����m�1���܏�@nD�XK i���0@�]�iP�xY�qk7T��@���p�^��H|�(��?&����>S%���w��(�5�S�O8Ѥr�-����dUA�&��6��u>��%�[2�9L Cq� ��^�WE�:˙�=�+@`r<�&k��q���йh%S�}6�̀���_�R�b7�G���k#�v"�[�*e���P�.wڍav�e�{vS��QJ_��^�P,�1.����GЄ��L1�-U��Г-��(4�����F^��Et�}���|$�@j�H�8h^=�"DwJ!�F�me����s�ݰ��N� �Iˌ�CȢ��hd�;���)x�ePow�X�f�����J���#nk�=������ .���Th��Z�(0q�]g�i=��zj�T%�_*uˠ��BJ���O��^��S�b�`u�!�yp^�*���7���&��=���>��k�e��H�����˺����x���4���~x�9���:��!�W�|4>���0e-��) Wl\50\���ߋ�?�˓ n*-G`L���l^]�������<�/�k�4�]2;�ʡg���w��+k]ń�҈l��WƄ�Q�F�\�6�Ƽji&:����&��o��-� F�AF�Jn��8J�7 w>0�-h�.�!������	�!CL�������_�li�9�s�W,[�oV����le�[��WJ�)��,Wl�:y
��1&�}�&ſfɿG�G�RE~�ET��_��^�n#�� ^�l�Y���]��A{�9��.K�:�T�y�vߐ�������SB!AJJ�EԔ2�;����Zkq�i���]򞫝9l�J#6���:w�@ ]��<��zA]�z��U��7VN���~����MD�sL�O��
R&G#�r�h�3�XY�u�H�L���ե�>���Ȭ�G�-�t���K �i�E�{��t��tt{\I&Pw���z9y��B�Wi�@�;���^�ZA�fa�:����o}y4_G����kz�W).��}�#�������PP*��Zn.&Vv��Ԉ4uZ���)�CYn�x���=e��0�*`� �L�t���eT�Tk��	�ue��`��l���X��?�0�3����R��e:�t-^OI�"�QO��V�B�����ØP��+u�'����7���!�3%��>��_:8�;���;��|��L���� �}6��ۏw�ƂB/�(������L(��$[���J3.Bg�����>���z���*�*��9q���s;w�r��_�q4�
��7m4C����V�f4��_�L}�?�����~����|`94�v��α����8�.�"#��%�`��&�����:7C����r4���r��K a\F?,�{�h������l�c��*�O"#���}v�[q_��Z��	+t��?f��ë�'z������=�tk@b�x��>���ǡcW��.��Tzcf�'�[!6b@p0�r���V�[�V]1ٶf��p"9�H�M�e�`$��x����]ўr�mȾ�RKe���o���p+����O�';�)�R����Ί���\��;����(�2.g	��ۍx�o�i@�6#_��`[�U\�	`�=��� ��X%�W���,�^wZ0�/�?�:�0mtp�N�5��>���d��Z	M�ւ@�7"/;�=��*+	��"��A�M4�nv?�Ւ��
��ȩ�k1r��̒m����K&6/��Dב��lL�YZ���0k��6~��#q��:f�j��z�k�'{�I�8��#��ZH?��Q��J*,.K��n�/��
��x����ծY�;l5�P�S�pl��Eo���d��-��M��f:Z��q2��Qq����h�b��q~t��a*�Ӿ�(���9C0�.M�� \cq	ߤ>�����@�<���ݥ�*����sr�3nb������Md��YD�V��EՄ�&F���:e�����B��GG��/����,�GX����/w-3�;d�$���>V��Q��=���~��>{Sof���,k6�6�V�1���-���e;錍�hX!�?f���_��,k��2f/�"z�x�%�)��
��	c����h�y��/�(&�"ذV�q+��a�s;�%��3���d3�bJ�1�:K���竲MZ�d���9JȾe��d��5x�a�!�f��q�K�U6�_o��|ȡ�|��u�8����:��uX�\_:��g!@	���Aji'a�=�jw�du��\���dg�O������|s���'��γsn�os��f�"�X߬����N��יؐc�J�rl�8��KQ�r��j��bї�L��K�0Uo}�J~Z�l���<��2����ȩ��h���դ���3����3�3{SW���#o�a[V�c��a&������L�}�i�语�[*x^�[����6VD�I����a�ƀ�a�Rd��F��8B8b�G���PQ�K}�����,U���6<i����l`y �T�\�S��lA���tC�����܀��h��԰/L�j�i)6��FN�>V�ʰ��RN���-C$��������!�2�ϱ�G�~��*	'X��{ȗ8���Մ�h=�D��K
��T�0�����o�o�)q���v
Ǝ�_��Ԑ���?�Uƣ
��k�!�=�g�`(��O�t.�n犢�DM�
2�����u�i��(���c��%A@��sI(6k�]��ݫ�C�2��$YNo���U�w�8l�e��;�m6[��!"�/���C�P�(�G�9�Q��^jN�BB�-h��8�Q���T
O��0�;	2L�q_5�n�d<O�P����>��AXf�9̀+δ��`.��f�N���Tj
~�Z�Q��7Y��!�����rw��ۇǬ(�T^���|V�fXưt\u��{�P��p�y׈�NQo���]1��� eR�UL)�2i��@o�Z���mݐ����Q�]M41���(�UK�g㐹��u�y28����ts��c�0��y]�
40z�./mU�Xe�Wy���K/�@�Ӊ��	K;���;�̭���-6�N��'�qƕ�~W��^��"���8�{�y`�4�+)-��B>\�h�ƿ����O��MDWw���W�i`��~A��ݮ&�m���hR�� ���~���gq__�.25���EJ޷R6h�P�ű�~�˫�5[�>�Ҩ��W�P7�\��_u�͂k�2��E�p��Z ��\�fr#�^�q�m�n�Izl~�q]i����|��pb+x"�K^��f[e�Dٰ�=�:�����~}�V�8�3^tn�� kW�|ϡ�N�U@1:I�d��GO!��jc>��{�ǲO��1�y�"�ߊ�,�6u�v�o��������Ŵ$��<��!���P
�HT��/In��k����L��_WME��*A�ڡv�3N&D�ٓޭ���a}i3f�_�J�3��
��żlF�
v��L�<�#_NEn�_[(/GI
]���6K�E�@)�5@�%t�E�����,F~�+:~�^��	�p���&��@���7={��8���K��}5J�*#�C(n�&��A���,gF�7ޒ���ʧ�A��g㴅[YHNK��KYs.�,�ݳ]%�d��K5��[;���m�'_n��H�2J��r�4�q� �X=iCC�ɗ�~���d�~Qly���9���#NWJ���R�D��o�a�s,�'��k�1�Z�E���Qgc��&?:c$��H"�a��3��gx�Ј�w�3�ݤ���d@����=,^Qz�_�@�F�s9�)��D�<�V���{�ް�[$9�*z������� I���|PƲA�Bxk�����Q��x:z���M�S�� �,���c��j�1!�/gK������8r䃁Ow��lΥp�<�8�`)�K:���i�*S��R���ۍ-��mѭ�IAB@$�a��;�9]�\����D{E��n