��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����]�V����9����D	Yp�,&�ƹ>i����r�O�z�J��X�������^�ꃺA���&k�S9����zѬPr��˶�d]��;�h��7�mںZ8!�ꡎ�u�6�-Z������. �w�+/��hB$���\d�?~j�����؇�O=�,���V��O�7#	l_rǪ�xL�zQ8�f�rB�*'��L��v�*�׵n(S�W*�k�_#�X��2b�CXRd�sF�*�zY�� �{�,�xs#���
s�Fз2L�_�'�y<1l��X�_��T6�u4����+>$kvi��j"�A��
�%�/���{s,5�w�B�/~9�n̲=iKE&�b*ysу��&(�40ȵ\��,d�0����%==bX؜���1�J����º�Ű�J��%�������\$U���霈�9�G٥��U�r#��La�}��r�m	�h@)B��.�l�o�H�[y��w���<�d�K-ړ�V�2m���1.�Hj˄�jʋ��9�8����T�U?) �i�!�57�/q@����uCK����O� ���6A��1���<�A�ӳ��y�_�:Ơ�m���o��Ǫ��wt�F�����j��t��b@҇�!=���`QpTg��+A'��*9��B]�/�|��K����V�i��mv@n�'Lk\Ӈ*�s�4-r_��vil�-��
�8B��,	X�^�Ky��ih��sr'^��7-��8�C}�{g��_\0�Թ�1� �^���H�Tc�������|�s�Q�G;ꆍ�s��#�w�0�*��f��bT��3/Un�p,���/K���G���6&��e3Z������v�3��t4�E�~[�����' ��e�en�']ѥ��G�"���'0O�F�P�;;zD+�-k9F'��\�j��\�t$ʗq��qj={�@�@�R	vj����h�.������8F<�X3h2ĉ"Js>��W�b������8������P��h�����E��Z�[?�=�~�`�EB���cvm�,�p$y�>��tR��}��5T�g �Qi��~Lق�
Zz#Ab3q��xx)�������5�uQ���df"���ݓ���o	��k-z�2O:���;*q�G�y�<�?����N�t�,�3B��s5W�I�����8a}����?��j�W�,
W�f��\}�0\�����!. �$�]���\��g�I���]�\w��ŽA�Y��{�p J-��Ҩ��[>${�#�Ar�6�.J�	��E�������P��:�>:Ƒ��G&)9D1Q�}��'Y|��2���;���=*!ۓ;�M�ŕߟ77޲�����;�3�^,�Z�0����Gqo=C���?Y�<��aw���Ӗ+l԰��>Y��n>���(�FP�w�1"�8�d�~�
}��q�..B�*V�f�Z|T9����4�Lŝ�<� �f���@��ڜm�k�;�������L��*�0ܩ�Z�j�l�Ա�a��Ȁs����߈Ђ�7
��:'#�:=X�ܲyf� �Xҧ"
?mɏ��o��_$�%�tY�f�=l�G�!ª�� n���·��Vy��! L��-����À�g�4ѽ1�3�iR��w��I�q��4&<��� �G Y�#�ɟo�1�Nc�H�[^�GQv:1���������b=�?JvE��W�|�q%��z�Ss�<IB��Q���)�/3/f[�r�*��D砏˝��	�9���a�q��d+�CZ�֣�c&��ڕ͞I�6���:$�~�α>�,ݴAcb���+�#ī�֮��h/�����Q	ӻF��+g��@=�Ρ�5��r�8:a��>V����b�3�C"���T��2=I�Ա�t��Ṃۮ�d�����Z%�C	5v�f�@,���oI'��d#_M�y5z��}����x >��NQ��W2A��b2�1�_��̧��jM{�s�֯:���T�Z�� o'%�R,�Y���^Q+>xа�zڡ:2FMo�6����St��W3 ����`YO���+O�������l���	g" �,���8%2���i����2 �o���:t��#=AI�q�l�m���Xa��@�t�nV��މT�����[G8��B[����B�]�m�W0���F�%d9Ț2�����c�t�uC]�fSd�4�'����ӽ�"P�2H��)��X�Jaņ�Sgt����v�c��{r۸��7����2�W��y`\���ɴ�xrY�t�I����u�'L��3ꚥK���i����D��G{H�7>�4C�;���Q7׶�s��w7���:e9��^K�����H�����Ì���n�E��8��#S���V�<��j����GG��Ў������KQN�䨆tp]�����*�\
@��N��@�f��!k(�}������������G�?�wګ͊�ʮܮ�Y�ȱz_���Ҡ�C�>�1�!�}	���'�C����W ���c�
���G��7��X ~?�7(-��.��p Z��W%|�EG'��L%��u�OB�L��1gl1èT́F�>��D��(��ѕ��s�~��O����/���V|�v�n��=A�}Ơ�����=�g��b���N�	�3�e��3 W����V����_#/Y�l�8���V���D�7���`��AKE�h��oi���ph��іTo
D�#�����2��O;1u4��#č�:���*�.���?"/���޹�6+[�Y'J"�����,�ӽ��P'��ۡߓ%Dԛ�?�:�ٴ��^?؅����.5��!������waI;S����VӞ����1�Y\ ��+S/�G';�Bb�5w��Zo4VB�PfX�9��N�!�K�S/>�.�;����_�-B�"|��Wµ;�҄|������E���:��[�5+ދ�xc���8���t[�����p��F�F�'�d�ɖ2�L׫�!�qw
l`�߅I;���������%�2p׌�ך,�f3�>)�hHIyơ!�у:|���@�j���!���<[�Hn`��Vd$"'���d^I#�˸����dė8�]ru�&�� ~��*^M��,	�j_uo���㡗��d�B:�l&J�[���P6���c2uW���[D%@q���s���bp�wͯ+�<�L�ԛJ�H��JI�|�N�����u9o�U �ǿ�n=a��pXN~�߽�M
���w�����6�3R�B��"�)���F̘�2�|��z~�7�ߪ����� I�K�S�4^
j,+_jR���BP����i��������-^u���p'���yA��e��$�	t���.�;�g,%�-����顣�=}��ܿ��:{��2�]���k�4�+m�1@D�S�T�r�Kb�I��]#&�Ҕ�ܿW2K��K�'3~���~��ާ튈"�>w�x���*�p'Ic_��^+gӢ ֽG�
��<�ggL�����zB���=rh��俨�(^�_����⏠�s:���f���<1��g�,��U��s�/>T<T����MѺ�uI@h�Ͽ?�N4��r]�Bs�]�]�B��������G�7��O:�D*��6UbkeE���y��Ir^��q�& x��L���f�T(9.ڦ�]D�Ѵ}jGI}��Lݺ�
�ݘgܯB�s1���^�m����OZ����x�~M��*�����rr=��~�F��N1��4���׿��NǾ�lX S�	%YA��Q���v�'��j��
���_�,��IV��~�Ǐ��b��d���P�O�I�XM$sl�'�
�k��(G���/�c���B�g��f$�m���=�Y$p�^G�P^�(C��u���}c�iU^N%yE����b�Z7�V�G_T���Ƒ����A��R�Kg�σ8"GQ[_3z�+Or;�H/c��h�c�ﳛi�ׄ�<���	�z��Ău�;n`<�� �{%�	�����u�m|f��ޟ|��)��,�^��m��plt}}�/�\]� �ӹ��:��pڝQs
��c����=hn"v�yz�Z7�l��6$�S���kZ���Sr�wӺمH��P$�gCQ|^�<y���Z�tWK����"?��e0Vi6vc%�q���O{C0�m`��m�o&��KÃ�
L���:��o�A$-����݈�fHP�w�R�T�=g��T��5o�^d5�2:I�1�����i����_�8n���C}:�oe2�)��Apfꝟ���Eg��6w`�����4(�w�<f;qE`@u�D �cI��C���2pR�u[H>�I�N�R���^_{9�Һ���h���3�C�|�-�d��4���i��A��HAz��P�b R���i>̏˱��8y�P��S��7��w��P$�쒥w����^��d�Q���T2 [���m#]�p(�aI�GB�6�i�(��'�A5 �,�YBy`<f�k���z9�駘[���AS�"���;�qF$0]�E�mB�<S,ooհǅ˃q"��⦢S��:&w�Mǚj$m�NKk�-!�N5?h�+�rX��j����D��6�IL�5��ٲ>ƴ�����&5T����8=R�f����`?v:A�IQ�1:V�����7J/�Yqs���H�=�AHOBJ[�ߜ�K���vF_Q�&�Q:ac y}�����������O B-#!��5ѳDiH���H�) �O$�� �X~ۦ}�e�m���>�a�çx5�/݉#�����ܼ��cq����P=�=�j�a2\�n�����zۦ>U5֛*g���K='d=; 6�g�Q
��u��WW���Ô+���P��'*κ���4}�n+��,.�������&��M ����R�8�J(�ņ��Q_�;S��$�r����m��.���I6��|@1�]{���_�D�V�u�?�%�¤ ��S�q�`��^�MDqM���k�UZS�=�U�7oC�I�m�[����g����cy)a�"��r��O�G9 �p�K%@?�ʎ�I�t�ީ.ѷ$^�-��;#�U}`#nu8��u�8�	�I"��{]=��`�'�>h*�]�;�F�[(L;|�I��Ô�����3��ǰ���h�i-֫�W�fF�Z��=i�^c̓C��a���m�,�B�}����jw	������'�f�)�n݈Az\�VL��ɒA'Q9^�����Z�}jJ�Nci��T�X�����	t]2a��~S�4&KL<�M/�;&�>�
U�º�E��@y�s#ؚ��Ęl�5!���U ��d�Cy2�!�q�� 0Aɉ�,��i9xx
�>V�>Ҡ*\��	��aD*�/[��a-��^�G��n�)'�@��e*�K+'��RƳ  ��G��������γ�3q�Aϟ��
�>�
`��A*w!ǺR:l�Q�����E6TG���(xB��.R���{�x���5MAt�Y��Q���us����,�	��ŊJ�BK��x_p�NgK`� v:�=0��5�~�^�&}��~���@O�1�I���Kp4o��T����슰�����9�������UW�����P7��>�{3�����~������hEW�S�C��$�b@J�ѷ��fH�\��ox6ſ��c��.�b\nE}%�γ�\�5�}����kK�3]�V%��X�2|��Iu�@����w� �C)�{C�Q.���k{T��>�t>/�.�Mzd���-�t�R�d���b8!QF��/LD�+6P ��n2̧�����7�^^7�K��m���R�K\��w%N�dF�~�
%�Ǒ��(km�k����O�n`��G�n��5���{�ȯ�W��փ�2g+N;V��8W�Е|Eu�n7FN�ƍh=�9�h�oVI	������R��X�ц̮]��H��^��b.��m�㍡��aU�r��D��o����r��/���~�
xA-�.v�����}Ɍ�I����Q���;����Gҭ`��'���9I�
��lP�AR�lp�x�pks�X4����gU֪��MѻT3�<�R����FQA
r�>�D�a���F�i��D���Z����_t���b&�rP�{��ip;�]���L��|��GHU6A��i��Z� �r�CMW��W]R�N��a�|������w���;��1��aSfh�� k�5��uc����9�;\���ҚYB���hs	
��=�7�,�:��� �7�Ao��y��!�5��>hR��V�����#�#]j�M(q�vp1�M����Ŕ�fP�F����<�H�P(�9 ��|���9�U�'C�+�.oW=|��FsY�_��է� :o.���D��UK���9�BҴ�ڮ����Kx|Lj��d(7�����:]*Z�B�T�,�&S�e`�4v]������ي�Cb��O|6?�z�쉕��9���)��D��Ч�p9�l�ؐ��Z�`��5k�{Ew���vzA{uz�f���)�_��l��X������Kz�5:X?cW��#$����`�(���˶[�;_�2<BFr$c�l]W�Й�Q6'���k�x���T~�/���0	Co°�4���[pM�Y��M��Ѡ�q�(�xhm��))��V@�lVQ�:q�v�z�bi̓T�,�oز��9��[�����C?|�3s�3�C��>_�`����c����:��t���o๖��R���@�����U������j�h��
�� &�S��&��.���^r~`�Wͮv;�{���iċ-c|8r�ü�,��
�oF���,�[���6�Mg�j�-�%�aFuVJO��s�zy�����\6�Vn�����:��5Ý,�w6���������<�(�m�,�ԩ�I��"Ν;��.�m^y������0��і�\w�����pK��|�S��/ouȒ4�=
�2q�yt�p�} :����my-UЬ� ��P�Q:+?O+z��"��������K�wS�Km����ּ_֣ͦ�#��8�q�~�����=�
f$����}lр)ꁨ�����5�i���ҋ��#���!G<��Jݕj��
ވ��5�(�O�Mb�Lvp÷c<����G��^��+k��� �ƪ� ȩ.f�ȡ�4�8ɝ��� 3�?��lSm��: 9^%�Xn8,"L�ܯ�%E��z�ߕ�5&@�x�]�Ut�����U��Bɽ�����������~�h�\i�l��/_0���V��l1D�;��r<��yG�4�F��Ĵ�cn+%�٦��\�sku�.�$�������])����j�a@*y�1F�[M)�&A�gL�O���w%n��[���1���oaJ@��H�D_�6EI��߄�4�-_@�"Ba�R4~ɼ��d���Vٕ�<㉉A����f��|Z8*�x�ƈb��!�J�鰅����ğ�I[�8
���s��K����^��ʪ���<���C����Դ�s,�6�T��Y����~3p�,A�ym��9����Y�l�8��z�<��e�j(_������,��H&��!�'�{6�i�ofH)Ѷ���
\��Hp����#ɵ��B�����bv�]��
՞�xj���@Y�#�"�����W]��4H_�&��� 'D��Ў_����l������9Fj�Dn�Տ��Fje�7�Ik��Nj�Ѭ�E�l��B����j��ݦ�o���t�cJ����:�I��OW}'�`ҞAΎ��T>����������U��F�,������墅�;6�z2'��o �19d��G��̒\�]���Fض���c����J��Y����B"�C�n�]T�uG�"���Uh���U��:��ݍ�k�[S�RpB�@w�
50�,	m�t���8��*o3��Yd�;��JT�+������.QG� ^�c�S*���U͓X��`^���� Se�y ��*=��	ns ����1i_�CՍCҍ�0�[���E�VcQ�>�F��}���	E�a{ޥe��n�l��mP/Ѩ,��y�}����noh�W�Uj��|#���<5���$��m�<AF��|�9�Mn	1�_�"_��Pz0wa��N���a�2P�O�/+�i�^�d+��0gݘG�t�%���D��U�$^�l����E��
YC����S{|g�}ğm��`*�]��d{^E�[�%=#.tr�4�
������ϲ˔� �/E��'r)���R@P�׆�(h�U��z�\��>k�Ow/��m|e���$\K��UKԄч˶�TF*QXd�I��p+�&���C(��A�v�̏Ú�i?����%����-�5g⬦����dT�y=���kލ�#J��}�E�6�&��#�9�=t�����VU��hǉ4"q���>�h��A*w( ��j�eM+;��Q~�겛Q���ԝ ����^14��A����R��8-�L����{|��_*h/SM�nÔ��,0�rG��vUE34�d���_c�Z�������5S7@a�6-����cВƈg���r��ΛHޓ��n�Pl��Z����'*��S[mub������~�	M`Z��j}z/�g�C8�~V�7c�YW�cD�r������KϪ�T1����ƫ;t��Eb'�X%�>��g�e�H�b���r:c��)Ϧ��h�H�8�2��	�h~��=Kq��Ikm��!z�Ə��;�ɬ?���'�g���w���,ej�Bge�Ww��p��ߡ��S�A��V��s͑��e�����uOK��0"�Kwz��4�.�S�ģ�A&'��-3G��Q����b��%��d^bh�o eN~���{`}\ـ�ϑ��2,Y�rK8n�a�}9���