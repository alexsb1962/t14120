��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����߿�C^���
�|0@��V�.'��I��>���	ړ*D�R����a�bt����b�Iق�e�}���X��n�� �/��C�yq�89�a��<�Ѕ*J��C��u�_�P�5��*�/9��B� 3q��ɼ��*�S���8�ȬbZ��B���jU���
��J��
+D�.i����4�΋I�\��� �ir�Լ^:��2c�1.�B��FD��~����T�]F!�1���Kk2���<�<��i��"�M����L�V��+g���j'������X��֭��+�}@�= ��B�����\&�JM��q3}�V�_n��9J�"n���.��6��%��@�Dwy�����5�+(d�ǾAG��]�P�Ig�������i&���Rof���;S5�����)��d~6Y�~�N3Ӳ#�O"�<�Ɵ��E�2~��lP\��J~sa2�J�7�})��q��E@D��!8��r��m0m�����+.)�=�vV�Ѣ�R[AjR@�B�t�� 9O�R(�]����:rh܇Mʇ8��:l��)N�@�Ư���2���I�Se.��HW0�^f�o����,���L�q�B�L��"v��3ӛ�ǡ�b���+��Ob�7��j<������m].��P�MQR*B�4z���)�a�p�DdL���"kx��{��Е�볯�����7��#Q����Og<;t�^���K#;=����=��4C.��4���<
8������B��(!�!O�?D�T
#���?�(��%"�� �B(K�0���B��9O
ͼ�PbP0-��0T�<����9�懣�G�D�
�jV#W���g+�1�I�CR�����q����O�e�.����*S��%ei�����K�B̸�Ke���ss�g��P`�SI�I�$�yY`�#�&~&�F�Ӿ:����߈�]Ú4&2R9#oԟ@�������2i�o�(F˒p�>��܂�RQ2�$��!�ny*�/!�V�G���ګ/X���c�zY �'�t�"�=,�|,'Գl�U�R���D'�L)�Q�}1T�Jh�%�B+TV3�g�_uG�;�d&"|X�`�
Nǯݘ	�^���&�}�J�s���z��PFF	�3;b@�lEy���
�ufm��y��i�G�8�6a�O���7P\r�?=�c֏E��t���߉�:�+�i��,���w+h�bȋQn��A������H�=���c��?dؿ�܇[�� X�M�ڜZ�B0 ������zĿZR��m�U7�!����M\8$� �P(]. ��)��f��R9��U¥#�0< ����H'mJ8�� �T�mY3����_u1E�+��]zGw��l'���KXS����᳇Q2�PؾX!��pf�-!y���3m+�l-Zz�Z }X���Ұ)�>��O�ڮ�C�3ڋ,Nw$��]OrX4����|��G#��h��}�K5Xo�;��ՠ�lmk:2���d	D0���Z�+���@��<r��ɫ�� �̴�՟#���՛�t�I 0��c-<�F��3m`��*I�p�P��^��)���:�N�#�UE�Һ8¨��W0[���f|Dh�)��3�`lW�"�A?�l�i	����/^�	'q���s&4��E����&��
P���o�EW!rx�W�ia�4����߶M�n���i�ֶ�8Cؐ{"5X��yƘ2�]p5
�qX.��8Lو��j�.��t�1T����l#��tM9��o�ʓ 8�C����ؾ�<PP�[i)��ק{�5gǲ/v#�{��Yk�o׶R�����Շ+JO�$+��R����^�d���(l���d�����j\�T+�JHJ�.:^�,��22�oӫ��yqS��s���n��.3��V���6.U˺�6~�I�hE��\��o�	h�/�҂�/��ˊ�1�_���r-�G��
���ҟ��)�ԾL���ْ?&$O��m�
��v��o#��5���VS	�f����Ƞ��Sc�N�&��zf�9�4����I���A=`��>�����H�>�	�3�2bٞ@�d� w��W��u�yI������RЭ�'q��TDX=�o���-��U�z� +��h�ӏ�c-�`�����mߟ����o�Ć��s���Q\"�"�
�W�����v����ߍz�am]�`ŚU� �[� �]!Ŭ*P��E�>�ܷ�K��r����]�Ӱ��F:�4.�.�.q�xj$D���T�V�E)e?_֢���Mq{Pa�y�7U�^���Z�氇���Oȋu��I�uF��ǣ�쉩��Y�A�~f ��0{|lXΒ_��Au��>��i����8r�f�p�݉MFnM����kZ���l�Evٍ�(<厲�Fp�$':-�7����j�0!_ �2>�*��@�����k��t��G���� ^4�;<�<U� � � 9�SR:V�w�sBy�lɐ�J� 
T�y�h�,���xs�n儩F�T3X��'�H��,,�V�E��V�K��؎N"BJt��xm+�ސ>
���l4��|w������ր`դ����x&m�Ĺ�$��F���W��vD�&OI���_�9E�@���=���i̴9_pKU����
e��1�9{��f�s<��A�H$��Z�F��z��搦JA��8��D��j����A���ۚ�,�x���;�Y d�:KS�1�[;�����k����&/O�R�:X~a:5� 9�.��Y�%~��C�!�
Dq��W�/�٘�ܲ�y|[?E�����/�+7�0XX�R�0� B
@G�lϼ>���gt~q�{�C�� �ǔpJ�����p3�Wsn1���,�So҇AMOY!TzVu֨1�EѬ�l<i�" � ���E�n�\j^����;x&�ߐ.ק�l;�S����y� A��̽*�Y� �[ۼ^�W�r;u�8��j��5�w� �ߴj�G8w��<(Q���*^Yi��5�Շ�R�l��\R�Ob���>�Y�:�1U�-A��a��I������b:f{^�l�+C��_��e24w�}������R��
��
������@Z��"��f~�J٦]N�"���ՍlUb����d�_Gf��s�FTܰ۬�<�� 
E��5%��D�	@�Y�w$b~��ՙ �	����F&����P̊�*�H�>e��'M^�����a�-�!��7Em��#��<�Q��t��4���
w��Ϻq�?@r�$.��]�p�H����+`��HA&�0�@V�\bye�Ǳ|/CU5E���OM)k��u�f4�7UH�]�ODѕ�D�C6/D�*A�A2R6×�4��M�3;�^	�"n�PG�.)ls��pNg!K��7B��&��I/UL�OH�iM�I��I�߷����䆸����k!5���G, l��ݚ����_@�Q�.�!���H���Lw7��\X]�n��{�0՚g��*���*�X�\�edw��{z������ܱ�!�]̘Ps�.��'X����O�u�����;"S:����{bW�!WpҡKn��	Ԓȗ^m�7Ͻn�f3�&�]�czM�wH@'9
ښ!ml�+&��e��0�e(��J���1�`CR4o��5�I����K�܄�O3����v��}����ʀ�a�^аb^|�ra1���=�}	�.e��Y�M*͛�E1`X:sEG�1E��������W��[-���Y��Բ���Ĝ_+lG	���]�;	�Կ�����Z߱��.�3:�M}��V���t�������&GC5l$�Y� ��А�u����>�[���Ž��D����4��r�VN,�O�hN�B��.c�힦��ye�T鵼��<>T�';��)���cK~<�QÃ�U1�����"�����}݇���'�?mjzM^�	�L�����݋��%""R�6���ʝ����n�lU���H8�A�'le.��0� M�8�BVn���f���xX�%��?� ����WV�WF� Ӣ�C��}��.�!���bi��*���~���zaB��ג���Kӻ$fF��4-=
�ۨnW^S���u�����K8�w���6��G�Sȓ@GU�*6��Ϋ�axʠ�_��mPT\����J��`�5�����$�E��yT��Ch�9LUj��3����;���/'��`�����K�F}Y���M�5_�G����/z���C�
�{*�ֵH���{�ݸ��B}�ׂ�4%Ö�y꧓��8k$l�6����~���c��3�X�W����v��=�r��!N,:�% ��s�N���o.7��I��$4WJ��@f�B^=���Bt����# k�m�޼�4��} ����pj98d��J����Q�n�ʳuu T��hn��B̐H��ڹ�S�D�*4"A�!�$[띆�?j���?��	���P��nP 3���] �㬡q�R���.hU�Rf#;'H���w�z=���3�6D�nǖu��P8�P	��� �Qp�a<�0�� /�n.j�:*��k(����yʂ�Q��hfn�� g1��*�7��c9Pb^`�b�@�J�U��K���0�/?��m8�K��l����<��J�ژ����O�~4R1�o��v�����UH-(��\��ϤBZ	�\�M����s��"J�	pTT.��ҙ�HZ�
ѕƢ�N��)ꅆ�p�u%���}�xRs��ǒ>}�ݬq�D�>�?b�8��X�v��n�&U�Ӣ���� nѹc���n��uG�Z��)&�Ne1�F��'4�,�h�a�Z̘�K�44v�S2W�WQ��A�L@��3-f۫p�`���e� i��<�p��;�^m����z%���၅6QN�B����p��ߵ�nB���+���O	���U��?X>H�:w闾��&��C����Ow�������IaF��f�LD���/�B��j�&�C��R����.h�Y���M��d��K�%:r����A2{�:,Mi����DQ�`�A�tx*��aM����XZ}4��|�74�Gn�*oz�K�XZp�մ����9~�b�8/�.�X��J7<��L]�
@@�=q���D�/�D�[��~f���d'�k�J�����1�il��"-�sb�Pk���q��\8s��F��O�k8{e\�ANU�c�Ȁ���ŵ�J3b��&S�R�;"k�A�!wR�<#�1{l]�]�a��HFa@e�����)s�]d�;f�).H��ǘJ(���";ۮ�ꉼћ~|�Łֲh;���x%�g)#7(���k�!���Bpl��](�/U?����a�����O�qs�!��ѡ�f	�{U����r��p53���@MM��(Z?4��.�X]���<6j���g6��e��韜LX��Y�/���esV�JC �R>�t�ۋN��&�W5c^�;c�X���~p��hũ�Ө�YW �Y]�6U��M$���s7z�pL�No�'k���"<N�閫��s9���/���0��&�yp�W���P�(��h���N�������`�բ�Vom`d�yfx�q�m!��q��B�J����8���4�.�*�tj�b�9��X� 'qE`����u����}�Z��?g g��{gkWV/똠�wu����2~߫�U-/��7�nc���&&͈}�[���7��V�ݻ��1��6�"áWO��/�6g	Մ�Ut�&��4���1`$��/{��������ܖ���Dm�p��7H �]��Dé]S)
G�=E� ц�x'$��Чv=HZ<m|��W�� ;$.$)�
���BKR1����=�!�\l}�"����;���#�6�� 0ncŀ	�Ε�^x7��|>[@�E@������"���F���?]i��B`6�XM:$'�1I�y�b别Ju�j[��s�\Ż:�$�F�&*���ʔ�Q�V��ʹP<�5O�oxX~>fc��ۢ_xv���_Nx�U-��'�F��,-tc:k�#�)��3���;��K ��2z�ن�`�*8��#n�k�v-�/%��� K�|k@�Tb����dn78�����rZ�'�����VW�_��Ye�=�0+��ɀ���w�x;�A�I��BzC�j-(����5p�ZV����Q�K��﩯���$�K�
]�"�J��p�:E�3�!����2�{k���V�&I�d��x8��΃kv�cK�)��+.'�/?�]�oj;��氟d5ڑ6���&@�G��T�}bU�U�x/�1�&p�� Ψ|�����6L	�mtur= ���v�(	� �y���J���-4�6�)�$rQ��¤n����_�o�)���'X2�b�?����s��G#G<��������}�?RF��i�uQ���_�AmR� ���j�����vI�7HHm�5���9�{4�@��ˠ����úy([�\CJ�4E}��y�H	�a��Y�<�C	��p��l�YE�Q�7+=U�&D��L�˒գ���X��Bf��eN�kRS�ҥ��}��Nl/F<�	�#�W�*�&~��%�c�J�_
/G$���7�E"��~8=�EJ�}�a�/H �nU��31=#��~� ��E�'9�@+�2�*d�T[����=<�����8�"��ta�*X�#�8�S�|�s�CR6?��8�Ԙ����9�x֋��=ӳ_�@A��!F���5�in%c�di_{���?������禞$����q#�d��]���!�zPK�g*��	Tg��u���� =Fd�⸫������)A^M��J��!Al:qL4�jxE-,����!������V+FZ㶫�.IO$%b��"��ĸ��ɀ�4����L00U{ H��e�N.*w+���1P!��&�o/|�ΜxǱ��$�ߧ��O��IH`P B�\�Ȉ��J<i����1s֚�i�9R����ߨ��
������	�L)(vΩG�Kj���n}C� �/��U�mGE���bQ�c�w+�ju�]�˩� �xW~mŜ�	A���ǒ�E�CR��)ٿ�9�=����%�w������{0��:ǣ�ꞝ����C�Gn�X�iGK������N6yC֩=CM�/f�N�M$�F�{xpyDn$�b[1�y����y����T�YwCC�	E� �����*�Q��7�T�D�Em�i��!�U�V��<QK�"y��� ºr�9Rޖ~�wL����x"��^,��hm��~�&Ʈ�����Θ��)��2��K��v�0�D�.��+�RbS�	�'��1k�Xx��lI�͢�;f��vx����~蓖g��.�+ل<����#���]�|�٭q��f�&{���?�Z�K]�ݮ�4dy��[G�ހ�AW�-Jj)�}�@� 2P��M���S���΋HIY�-����5Z�ߵ��B��c"�A.Fd*-5��"LӒ��I��v?�hV�୞y0�pH)�<#L�=f���:Ӆ$p=�%��^TO��{��g%��̞�ծ�WH{�F!��J�M$�!?|�����0���� /ܫ�$���~Q�ؕ�5��?k�%�d���+��C�e	�@�X9H����-��sN���\�w�㇝�婐r���%���6"�^���kbr?2V����$���? @��`�6i����4yl�|��D����J�0'�°#�Yg�G�aM���ʛ���V䒄�a�7��,�j*��P\.Ft�(�:j�����,���(+�-ب���7BGc��#h�b�2��,���	ջ4��9@h����U:xFGܤ�$W%@׿<��"��V�.bk��*�P]J�:����S
V�X��<�K*�~A>�^SL�zE
L�4��i�t];(��]�T_֬�q��t3E5�ǧĢ2���M�F��+4����4�k)�cF�؝`���+~�o�кt�F�(��p*O���O��(o.w�r���)�w�C��d�.C�����W&�"&�5��TO���<_c4'�7'�z& �N��T�v�*B�և�~'�N�Ќ���^�{j��5��FP2P�Q�0w�n�iv��i_����h]�""Zz8�0�
�*��E���l�c
T;�`>�վH��[n	�n��Q���!<脡��_�)Ey(a�Ɇ�:qp+G���Dƃ?��_9�
��xE~5^��L���͌i��x����|)��o&�z��@$r:�S�c��ʛ��l.�{ibŃp��o���m'�	{}p�`��@�5��>�I��6�f4/�g��F|ɼ��e�㘱��:e�6ǡ4�4hװs�ܾ�xK�5��_^�rWV��g�(	�]�� zh���q�c�:*&H�^�%����Rbg�g%��̣����H	ZNZ)
�_�=�l7m�-e�0��D��O�%B>�%{T���.�OnDX�����4��J�r�c6ƴoMW�q(�y`�%S�Kj#������] UZ)-��pNZI|��b�9��7���t��	�Cⵓ-�V��j):��G�SY �iKfQ�4+���س���i���ϊ�Z�)�v-&�4��IQ ʪ�ņ�D-��lz���ܦ ���[�o݆ܣoS}�(���,��|��C#�ϱ�E>ߌ�������U/��5��hP�0]*z�m2C��*�9�q��纭�9�f���,٘=P�e
��,_-J�($^~`��b¬�D��޷Ġ����G�Y��Y�X��RT^�8 ��5����)/�`z_�� �Z�m�_�#�1\������]tX����F�2Dt����[H����k�Y�:�ip�����*�:EDr�*,�f��k�F����U�k(\%�)[�:~YL^mj#)»�}��['b�#�h�1(��J��:T��-��Z�n ����q�Ҍ�WL�2���vMuЕ��!��!W�������#.���%��\4m���O;�Я�Z�j����J�h[-b�g�K"�� i`�V�:R
'�cF�NN�Qk\	a`��e.ޟ�O99t��䶑:+,�BH����}�� �f�[��)�g!�w����ٮ��P�ka��,M���\�����#�?��D�|�!�A�:�G�7�������aCJ����~�xZC�Q�֔�|�����hvL1<�鏽�Ϫx���H]Ѧ��S�fvr|�A�i������������a��VD)ؼ�h�:�-�m���M�mQ�C�����$*o��~����������d��>�=�y�y�| ?�H���ϲfˮ`}�89��4;�N��$�h�Z��<$K&G�k?��2Y��PU��{��$:[<�Q�͆�Y�*�IH�z�FE��_E/�3��iv����U(�����@��Z�k��+�2�� �@�J����F��´�=_V.�#�+�o���`J���SW��KN�5u�1QO���j��p	��Ez��A6Û&Y�$o"_m�gL_�)�Ӵ�'���š뛔?,�E(%�/<�?��"�' =9*""3{Ƶ2,�g�7�ŧ���!d�¦:�?��MxK������/�d���ѣ�g.��h����n��F�;dS�<���"�(XfU���֓��R�?Zt�W�Un��{�Vbī���'-@�o��}u�)=��w6�G,�Ր� xE���M�y@��_"�A�pI�x�({��y��:1�]-�� ���}���4ҽq-��+�(p"����{%�A՗��o����_D��>��Nլ������MZ�R�=�d_#�Ԟ5#b�Y��P���E:ས��ѝ�y�jz*��ĥ@��x��~��ٖ~ z)5a2�II�j�}
'v�3��5��#Va2�	�D�)�p��!�}n�)j; UW����������,p%r��;��G���a�v	�}�!�h�Db#�/t;\|�[��������N:��1�΄�b�_��&E�E!L]=C�aʓ�m����zc/�h�$�2��~)��\p"L�N!t��q�(O��,V
d'+�((k�G J��K��HX���"�h3-�|��kL����1~��t�[ea궩cB3h���Om��RM���^��ͼ�I��/���P�0����.�$�Ր���c�H�<®��By�rP{IB��K4�*N��N���.N� ݓuEE<�ƌvpL���ˇR6���v�V]:��h���W1�w�I���O�^�K�;Z]�(�_�������=�$,1ެҘk�Z�C����Zx
�ȳ����V�O�9!bk�H"X��6���k�&������ާ >����y����?��ķ#�h#���J.+{�N�#��B|q�<����/���ɳ��w�U�{!bz�os,����zĸ�OyREI6�h��1v5�Qri%CB�I,o��o
xy��">Z����DU��-L���C�6g���?�����v5Ƣ���_v���N�� �,��2>�N���T*zͶ6M��B�Ul�$���cga��a$TdB�;��n�w�pu_3tRӫ�����x�L��#1HOm�0D1V��rD��j�{qЦ&Dj�h�T��3��ČY�[�����*�,�vy�*��̫�/���r�@�ߕ0�;⿥���{w�,ܽ��U�XBָ�B�?f+gWݐm=�\�Jr��
o�e���i�Έ�Ne٥{h n ����A^�r����؇��Y�>�c͗S���3���i����,�f\fsj�u�jJ�|�� ~MnWb7\ɼ�I�׽�lpr�l�f��3��^�H	; ��l9<ݷ���:��X�a�L�U��l��	xP�q�ba���eRL�:��T��4ک\������4����+Ѭy�*���a���� ;�ɽ�0�\S�	�#���j��F�:S��U��h��*˘ D,��j�K�C��Ŋ�-��J�_�4[%~=��I���]�=�(�Sp��KbϾ�2L�xU�X��秪�۴���{f+T�*���չ�ː��\��S�pI
}d��fiu��y�Yry�e���.��$�ԃ ;2bhl���2O>��ݳ�~��e����6��>�R%	��o��M���PӸb�E[����$=VE�|����Mj=#����)n��,s�v�3&�Ţ���8�mol��O}��Tv�wS���)"�sg�N��I./o:#�l����$�BM��L��*-�vͿX�V��Hھ-���h=���@�q�z1r/�L�� ���Kz��~� �f��m�ۇ�8ݪ������Kl��s\lB���J�C/��\�"�-�ؑ���P�(߅�ŤLN9L��lll"�X����I�tf9�I)ld��cn�Q�u����*�ǋF�W��e�H�8���!�ȋ����$ؑӆ�pd�S���T �����$Ӈ�6��:
Un�(gz�8/�%�^�ôQ��l[Ju�d
���Z) �� ��=���0������R�"��F�#ٙ�M���?�cE��噒3Dhh<+i����\���3�=�t*{b�־��C�����8�n��7h�8 fQ�J���h��fcR�}!b9���j)(���-�C-�J�k��l���w��$�g���T~@����X�Ѧ�2���{$�^X�� A
DD(4P$��h�W�B;W�"�±�����h�+ؒ��Fv�������0�6S�,�GP���'�8fuW�*8��ݘ�g-�`��b�狚k�?r0��T`�o�#�a&B�(�'=b!��$�'�t񿞰/�س@R�JvH������nv�$� �8v�q�Ylt���Â1.e�g�3;d�8A7-Ω�J���$��2��Xr�2�ʩ��<�:�?&�����\9s�|�K����W�]��e4Q@^��W���f�ù@�by�a�Ф�y�G[a\�p��A!�3�N_�h�\$��F��{V��/h{�B7r��e�"H�}�� :ڲ�Mܑ��0Z��~p���b�W󧕆+"4Qڏ��<-��WϻNG�Vv��F�2�N���J�����䄜(?��G��ȵh޻?���|��
���xBxrN9c�N2���?��O �D�o���PpR|h�lT��Y��+�E��;v���'�o�8^��"���հl���� ]������ ��1Kt�������f�[\��w+<[m�&�Q��:N�f�B����&�4�o�����#�R� 99k�$�E��� ,����h���@��)�(5$Za0����~so��� D��>�fJwm厴�|V$[�v�0a͞'\A!��V��w�j�Ơ;�j`�]��U�>�3�St��&�af3,R|Y�y9�׻*1
��O:`A�$}g�p;ug=�ZR+��q0��{��Y��/�r������&�ME�/'�?���7ۤ�s���1���?r�)6e�E}, VT�
-��(v�=������%�Rݴ��3~�K�+�Jk-����mv/��y���'������\�y"ӻ	E
��E�W��cˤ��Ò�'I�1a��bٍ�����*;,aM'�]�/���W��9������#�uNyiJb��s*�-4�h+߽ߖ���l�Ӎ��I(Šq��F����I*�[���e�r��^!;���	�@�a��E��;_���D�����!�qQʡe�X>���s�M\������%=�k̩21��!#��6S��B0`!]�䁽�@	����w����^M����-i�� \�d�W��J�>Б"(�k�[�� �+N+�B�X���:X�'6s�}���iע9t$�fgϖ:X �"-ω�L��*��mr�#$�zO�X=<4`'(A{�U�ZR���m�U�#l&9S�e����J�4K�3��l7���f�L�j���Ru��c�E,����a@���o�sF=l�s�(�`J�Ј�k�
q��Z�=�
�:q���~6ko3���Z�
��ӂЀ���E����ۏ�7jxw���ّ����� `�i���%��揠yOӜ%�fz*;I s�W�m�/d�����U��T��H^Z���=`q�H�\�������-mr4�(�Kg�E�+vA�b���l�ӛD+�V�e����`�(*-\�����Vp��3<kF ִ���!)�s��w#x5C4�&��������7�:���m�u�B�5H�i�[s�X�^Bq�n��/{��LB�&dIO)�j��.�s�Ư'*t3s��+����=_�#`�KAC��i�"F�� �An�ڌ�u�'�e:� �_�W��.G3�����a/���W���t�
q>p�o`WH��� q�S� ����hR�l��N ��������A`��݈*��q"uV+����P�h"��jKn�3��m�T�Wsk����N7� 󩼌��2�5�@��%��p~a�2QU	D���%�F�� ������)zK�¤y����\+�[Z�W���L���ꞩ��,"�x{�6��)Q���]EV��.��\�K5����w�bc����̐.@#�C�f"�H�77�3�ͪ{�R���b{�W5��� �8-�Z��dL=7,B��;�xk����'P%��TuA�����RP�*�c�(3I��!�4�wϚh\aVwR�%Ǵ�Ѡqk��N��=����y^���_�/J�����<N@+��p���	kN5�3� �	~�%�A���Ia�{��_DI���o|60D8M�R���f�x�0D������n��:Q=�Y�c�j�����ٮ�y����3�k��~�ׇ�x�aij�$%ɒ�Qɲ	��(uΎ�V�|��4*�Y���O��A�и�)Ň��*TV�?��ܻt@0B�Z���.]�~KE�����+P�@dΙJ���]���;���E�k�J�n�M>��{5�w)4̐�4Mʽ�����K9�8jp��ڝ[$"�����������o�tdŨ��2m昆^��%)�=}�=tOlk����@�Ӛ��7FuA�&\T2wW6sC��-��j��7Z�?EA6D���W� �3A�������[:�~q0!֓w�Ud��UC)K��3[��x;�u��Jp���� �9�ȟ�����8�ڰ�\�]���%���q��"��N8�8�H5߽�)U ܴ8����q-)��B��CO��|�vE�Er��_x����J�|FPN�����A,
�XG����`6��素��@4�[9�~7�J��Y���IP�.�E{9A����m��tJ�K���uo!�V��d���X�kŸ���:ow+n~���b�m�-��JwTONa���Dj�OqpF��?
�Vߟu���Ri��t������!��A�$P;ߝw����Jb���md��]�b�BMK�ML�l��>8f�)8�N��|��?|�����sN�����K�;$�b���Q�j�9cRŨ�#�D�U/�d���h�����x��tE[9����2����_�m�]�� 1��x�r��A�T��s>�
$��ɕn�h6!��������:b�4C�����d�b?���<��k��70cz��T� i��>�kU�C�Վ��Yڦ���S�H�326�*=f[L��5��Ő�-���q�~�_&c����#ZR�n�|�0�Bc��;x(��Uj��03`�"1��p:u�I�'������7���U���VXWѠ��Hp�XQ:;���v�\�Ȗ�)�)�´���bK�G{2��Ԓ�@��E��E3���^v�[O>z��?�^� ��ڣ}��0�+~1�L�s-�y;bi�o�����o�K��B����)�h�:�NI��E���/Y��2���DL��u;6�Gk~Gg
�Tw��u���(mu7k8Mb{��^\��.�25�e!�B�������sG-Y̺=n���]��z,��%|�Ͻ����eZ��}H���W�8�k�(�LM�@i�����$	���.�
����!��;*e��)�pYz����鼓�h^�Ƭ]e���]*� ẕ���E���V�[�q��=�W*S�U�`Y��=!_�ԅx4���B�y;9�:�V�����Miul�d��MuZ@ .��nG7G["V�J����@��9�!9��6�4�����(&�X�T��B�	]>Y��(�f��s��c��N �kp��~c�5���%Y.樕��ϗ����
	�Iqĸ����v����Ur�؁�3ޤ���( v��I� �M�ެ�����,��@�i�I b�1�s��>9,��^0�F�<{�I�O���en~\�FV���i;�b�폹%%�X
te��K��)���%�����^���$I�
 �r`�n4�<\�}:r�Co;���¢�(;&�w�8Z	�� j�ݘ�`֙ؠj7^�ٹ�����L��?�=afkg�	��t>rO�S�aբFf��{A��XQ� ����׎<1�R����Q�ّ�ܞ�ëB�7R�@�q	�G��rѤZi���\�&��q���K�[�IY=�#�]m�����P�����\֭����@ٕ c�A� ���`ߵ��]_� �������}5���^D��NV����C��ZX�����32�2_�pU�AȦ셼���n��l�?h�1z�L�GA�<Hm���	�II����Ip�~.�J{�c"���{J�r���K�x-�02gZY�Q��! y�}����7�0e8Q��\��}�Ա聪]K嚮]2�k�KF�n6l���G�zmor�8W�����
�x�N���:�q�U�gPs�&{��R|\���R�t~��w����Ys(1�~j4A|N�^^
�+t�DJ� �o��mf@IA��#0Agu���_�"��>�&ٲ ��rl̂$.G��p
���C�=u3�1{�"@P=y�����[0??���l�ʻ� �E�����1 �3ՙ����;8p������Q�[=�U=%��%d��P�_���I7�"A!�El�I�4+,Aw��cH�1�a���&��Y�Ya��Rjl��g�g�kɞ�rĶ����u�ML.��1e�	̢\�a���V� kh��JO�5#S���}SMq܄�A�2J�΍h�k�/[����gɶI����˩���8��pS���p��:������o��s�
��g�E_h���%nS����'�su��o"�8�n�B���w��rc���~\DR����M�i���Z[���xe��	ì��gE��7���C]�%�ߌ�����e�#�Ds�.@V#�1b�ߚ�;����,<��$�_�: ��
�ۃO������������wׂL�	5,yi?�.☒xo�'�%��r͂&����o&�oQ�1�1#�'*��]#�����յe��J��g'f:T��k���g.�VA��Q�C���]�ߝ�D�@��,g̮yx�L�JX6><��יK�6:�I����,�lb�����.���r��ÑԔ�|lj�m���&��t=%Ҹ��s��g;���K��@2\��N[ծ�F�
���ԭ�'���H�z_�a�da�Qje�?����M5Xx�Ҹ�jN�RJ���F���#�?�Ǯ�	v�a/�r5��C\NF	�/q��o�9�Чk��Y�9˒���S���>3�K�}��Ӊ��pQ֍�t�1�?y�,��l��>0�%�:��IP�-��48I�2��pa���;�L��v~s2��G�usnY ��G��&�3�ǹ�,윊]��FO&�&	��/y�t@�|D;�X��j3�g�[�\��E12A��R�\M�#�SR��w�Z��O���Ih�B��%���� M�&
�f�6�����/�r9�8Z�u�֘��$�O�۲�:<UdXyZ���bw�2���*���9�~�帕F��y���֬��/�';��m�O�r��R
�X(i^�c:--N7
�-x�a���o+&NP�����0zC��#(�(�:{`1Ҩ��8�߾H�&��bفJ�ۋ�̨<[�e�ɧ��1�l31�PØ��a�����1����o���_,hm��d2�b6Q�$���A:A��F�+)�N׋x%�o��]�!D�Ι[�:����Kd���c��߉�r�WQ���JX(k7r�8=��7��SF���/(�`:�STZ��m⌰&Ҭ�CrGw��t�\=($S�D��e)�#�7��3F���v~���qi��ϒ�t h���7'�/�����.�(���ͯ0{�	�o����6�||,/���YbC���S�Ѻ��Z3�`�P��=g������1O�"1�)�����#v��U}�.�vV��8bv�=�Q.9��c�Hc����F�t
����J�wR�]��ϼO-��aT.�gg�(��z�}��i,>������4kC�\��T��FnbF���\����Y�C�S�?���1:Ôn���]�7����n�7C��k~�7�-����7@�hzU{���R�ɽ'�F�Xjl�[�����:d����l���-�PWK���2�#����+�p�Q]�`z�:���@��4!�<m7�x8��f��L�wz<Ԗ�su3]�[�O��Lo�w��|���uϫJ�]#�K�)�*�'�%���
��A��`V0�h����!���]��{6��`h�A�*��\�A���5:���L�yl�"�2*����b��+�p}�*]�꒫ ���+$?V�U���Y��]��>�� �ыg�X���>��=q�6I�2�@���w�)��L��߳�����nc��M^��C�Xԇ�^���o����w�K�[�z�~�P�c�^�I&N�h�'�����K�^�W��<'����l�x"S}�(m�R�v?�V(�K^�"?��
tK`,Q���l�"�1�<�_Kƥ�X:Zh�].�]9?3���d�
d6ɁG�y9���O% bj��ʌ�R_��R^ ڶ"�]n1�Z�n��W^~�~I�m���O��Y�p�so��`�ҝ�;�Ƣ%-A&8�i8�����9���D��h�J����7�#�U�<��N����{�WԻ���$ ƥ�ZC��U��A ��e�?�vԇ�M��_*�u�lFE:�g�q�+�D&Lo±�OG�V�P��)�g�~l��ew�ݔ�B�;��v�P�{T�l�Lv�����H�@�q�v^9Q�n�k����B�h*=��{r]�3,���\�W����������<�:�N�9}3��Ze}��
��������0�"�煩xv(�b� �ٮ2����H�Z���~,w�����@A=+M��Ҡ��-!�=���*�r]�_.W�\����xa�K�Z����&Ai>�R�R��n��MO@֛Sx�j�Pe�hv�X'���1i��g�@�}�\���4)q$���k���c]��H��no�t�m�t&��\�V��<cw,�{4U�C��h������S=��
7�Y[#N�x6�]:
���9��?��2x�K]G�������Kӏ���ck� ���fnUH����=�ʠW��+�<Nk�05�/J3���D��n� 	�CE��Uw�԰4%f��O4h�ѧaGY5��"d��f�����@�1�u@P��D>���x��?�>���Gq����1�<����nsE�w�]�n�Z�dm�4�*d���>�\��^F͆�*	ʑ@��eU)�q�3��PS�m�Ƭ8� �$ɚ�t���ZI
d�a��k����J��mJ�I�|<�;��Y�%k?�ﲺu�c�!D�(�Ivϐ5�*�Њ�fg�KBu�ͮ6��m���}�k�9�}�#5b75YO���U��(+�sp(XU ��
5Ǧ5Y����A<w���7��mL>2F1����+��z!�y%J��|�i�DR���hl溰(�ǚ����PY���`�d��~Q@%��bk�K����x�,
����H^��eݍtJ��S�<��rxLL\Gj^�$����e��(¥�R�8Mx1D���KĿp���!ԥH��]��bUKZ�EPĚS~���]MY�O� O
���x^k�fqُ����^̶�Q�׸���:v��	����������T�υl�G�[Y�#�"�N�k���J�0l��I�Fi{t��@L�� l��{ϴ����?��h�[�a�ǚ!&����g�e^\tP�H3�^�2�I-�P��[l��������m�3U^ݵ���5�W�7�M�N��!�S�� ��%��.#1]딬��s&���)� �ɒ��\�Y1A��2�T�X����{��j~�N�4S�YCDô�o��4>���������7v�/�U,+o��
]����H&��� �	
�#�-��jI��S)����$��g	��µ.�Od����a�,�E0u5��63��d^��q�[b��XNY�b��Ԩ�G�2(���n$��b`��H=T�4`I���}���S��ZM
�y�Ze�T6S�녷����W��'S��Ɔ�닃6	⫰�ɁZ��cX��B~a����J�f}5�)����]3z�$^7\*�?���&ZW�see��wo�����K��\C��Uz��sbL�	և1�ϫ�;`J=i3�u]��@�-2%�vp�8�6������ZoD��:�lנ�[$g�C-�p�Zy���{�8��on�\�NӪRϪ�`�rF�2� Wqc �_i�^8�3wG�	�$�{u�Dh��w;�#`sA%��}y��H,%���H�c����qC����m����$����E��"Ҙ���L" ��2<����`A��O��DB���,�
�[�d%R�Ѫ$�ј	��"����iΟ�orN�GS�m��Ǭ�ӎ��DZ֎�����	�2\C�Gd��b��uI�y�ߟ5�@V���v<0G����lX�LD-��[PXx�ƼO���ѩ0�B�>׾=i_�
�����*x��r}xXSu:�5޸��'�Q��Y�H���}P�.�.	��r"D��%��L��Ċ�VI��mM�bB<��"r������u��VC:N��5^�?�]?h�{�i1��.N6/�S��Ї�Җ�k�׉{_=��}E�1p�y�y�L#g �xː"b��A��F�c�a�nM���?�x�5�̋���[��d�P?rv�fBHS_�۲�v$���%�a"O���!���)Z�_���:<��;pߊ
���z�sW�"�j�o=4(
�\a����]z������C(�'�c���MK�5�*�M��o���=s���]�����q��頇AU]�qA��8�Q9�m�nI�NkrÞI�F�Q
���Qʈ�n^<%b�c��b9Z�>黡!��~O,�#P�� Ǆa���Gp�&�UH��`y�G�O|���y������?YM=��b5�:=�	����jT�,�>��6y/�sU��%�s��#�|�X���[b�6�����~W4�Ͼ���Ng�HK\���: c`@�F�Vr|N^��CF�j;Vƺݓ�B����s�������չ�X�R��H'�e�ld�z�>;E�;K%���u�{"���)�E�G�D� _��LPE��i�0h��29	���v��
�Rs�#����O��
q-��'��>d�JE?� LU(Z�*�����[z)ь�OZևL��BsQ���N��م!t��1sM�FΑ��PӇ�$����'K�ncx##�r���a;��H+OC]Aw`I������]q�H�j���e	<.ʤe�Z��ҭ�U>�#�kM�&;��@睷�ҸX�%~���cc^x��G���V�F@15�g�Q�w�\5J�if���_,�K����y���9B����F�Ģ�7�n[�(o�Թ<l6���Oo��K�*]���`-�r��s�u�k��9scaC������v��}*�Y��d�{�gˉi�y���������Kc�G_�e�Z����B޿�Y^�F��r���{���eo�}H���ѽ�B�%����˵O`\Y-��,Xi�LK4���'4��-�X9�Ό�Ǌ����(�p��<�AM����t!�h�(�aq'����껁��E7�h��4��_ 1S2��`sD��vٴQ��Y@+d7��'�H��]�VB^�ވ�G��S� �ۋ5$�I�u�rt_}���#��~K�f���DN*���,�^Z��?hOP�A�0�c���(�t��Y8p]ML� M�f��'���
��d�|�s]�n��ɖ�Fn~��CȠ��'mB�	����ū������ 4�>���|�3))��Hm=�@t��7,tv��;#/���5mDmX��lx�pp�LbJ1��D�}���)���_��Q��F� x��PC�o�s�H�>�Su�����UkS��&
�:����=@�$��O�"��j=��r+�ZwI����Ew�a�N^<��˕�QU^� (�W�842�����Q�V�b��F	>�&�����m]!���HKЋ��尊����4�1��ar'�ݮT,�GC�ƭf���Q��gD-�o� �v58�2�m��3UO�+�g���
&#��/���+UnH%��&�ۉ�5�����t�����`�����t
�/�c|߾L���]�S2uQ��t�l[���R�a�U"��?o�����c���2�e��yCPE��.�O�<���`���]2�-�S�@�C�_�����t޿�����YRaa�=�i�_\�O{r[�q�d���i���!v�ꉪ�\�#P�ɠ�7f�v�[�c�{S��q�WU�xn�76��O����ۙ`Z��.o6�����N�j[��B�xK4m�&�������%�A�]��39�99�i�/�m�(�ׄ��®�\���_״��qa�G��Tۅ���;+�]aa>��W�M������|~��#��� SiQ��l�����_:�E�'�<�pz6�3i�(1*���@��x�Xtf���=��f8�i��^��Oү$�!�?N��+��j��u3g�hQ7JU�v���I���W��.tfӰ��-��2;y�Q�õj$��/
uAӪ���Rx r���0�.t=fE:ddunϩ.��jb˥1��k�q��q�K��U��#�$�[
�ĳn4Lb��]|�G<.�{ƒTw�h�WY
�&��9�N�;�M����ҋ�	����I��r��ǈ>���F�涧�f9`��e�d�ȶ���u~]V��?�����	�o�V�j��#��@�;�B�ݎ?�|�<��Wk���k�S�5�iBn_��+���ȇC
����ʤQ�����DBD�X��PV�ia.�J����I���t���;�RhZ��q[�� ����	YnP���W����?"=�f��� m��3eEfI"�/��	70D�{�.�[*�4�r�Ct�$��-�6�����L(���B1�zڋ{��c��Y�EJ�6!�[S�n΋��)t
�� ���/fأ�m�i�[_���/q����u�$��7�u��^��L���|�B]�sCg��Ų����v	����Ll�Ft]U����)��n`!�l�S6���5��6�#�j�9��i$#Ǭ����Ie��i������kl���%˲��k��Ţ\fmͼM,�T��7P��!��@�:�QIO~(|�VＴ�p��ž�����Tm�m�l�4:f�� cFL���^ 	��N��|�1��!�8�I��]Zd��Bz=W���I��{N_���Qj���&���>�b��]�w�<�F;z����0�W���$fy�T��/�K��_t�ɝ]ぽ"�	��0��W~������YO{��| ��B
�,��c���Ǖc$(&1Ҡ�M����t(nM�5�_�O���>4ؓ4@	�_��f�TE� �%s��Y�1/�=���ػ�;��,l�� ��� D�DV:�,�	B�OA(��Y�#�M�D6�C&BT
�y�vORD=�T�#�3��	x�s<���O�>�b;ǳM	��Ԟ��	zV���*�߯�>��%������Bl��O�U��A^o�8U��6!:�"���b]�m�ͼ	T�?�P���@�V��-6�X��h�`�R[��T{o�px7:9L��Σ�S8�;n`&oC���m�'�ےg��l�AK���{�(i�FѪ�/��Oe�v�T�t*�X^����- 5Z��3���:E� ��DC��I9���$�g��.}@���E�2T��p���Ż_(ڵ2\���RƢ&�?���+�S2�
`�Z֎*),�O[|���寏��=�`�%���Ŵ�IL,��n��ci��~���)�z��Ac������ģ7�>~s�s�Y V-z�CG��'#.��%OЧ[�g����u&<��Ah̝��%��ur�!�ʘo��8��{��0�5>��a|���G�n���o*K�WJAe��}��`!�4�o�ٝ�i��Wt��I	��{w�>x����yܒWm�4M���]�^�a
���D ��	� ��V9d2�o�f��VlZkf��`��J2�r�\
�y�,1=9�B��p p@ȯ{!י���c�[�F�����5
'��=FT�u�&�9>G��v5n,k;� �o�A��
O�=:�)>�~k��{�C��ީ������`i��k���,��Hg�{^���=q�3��#�cG� 7_��2�7�A�YH�%��`9��NV�T4q:H}��=�ۨ�Rֻ�+�CI��u��-�1�j���t( �e%���"�[KK�F���i+2rKrCx��{!���f�r���#�����EOGn�m�y%t���#��z�MJ$��F���"�q����-���mFL�Ū<��Q�@1�>�55�%V���2v2=,�Y��=����@�����
� �lh9^^ʺj �'�r��UP<�z�0�L�x�Y+��{�psh�V�	dC&��E�I��Ƈ&��k��*O|�*�!OY��鶤��hЮb��lFF~���|bsfv[���|A��	���YU���ɖ
�������|��O��7`4ͻx�i�<i^�Us���S��d=�H��U�v�*N��9�a�,[���&j�^��s�-;��e��)�GL��$���_0>T�O��pi�ҟ��9�G���Aį#��y�<0�OUZ?!���M�2�EpD�(���t��E���.-O�$�1�����ۇ}�} ���'��雱Ξa�n9�ii����p�zaBy��fȟ���dm�_i����\�|���~��,C\��ћ�]��4+��s�Ş�o���M�����Q�/�e���������t�%�u4����k���[��X�&rbsIV��'�5mP5C]V�z+B��1�9�`#Mk�A9W6���'XuZ[4��n��I��&6ȖO���U�j�+��x�y�{�$J��`,�=�U3���HL/����HV%�a8��vA�A�%k8k�Ԡ��r�-�5�H�;����`�K�g�R�C$V�y���p�&:D簳Ra���*�s����s�M&m����#{�\�KW��jY�ZI!��,h傲�I��^��ԅ�7k�
������c3-�J=%H���۩��0W�?�b,�^�J����P�!��'o�N��1X�I����y�ۂ�@�×hĝ;�Ĥˤ˱$K�c�@�Pz�)��
�����j���7
�l�� M���FW���2��Dg8'�cr�M[�\�(/�>�W�����f�T��?����8hu8��	 x�E�w�W5G���7 '����w�m1�3W�[m9�B���v��4�1*�@V����&(l�W0�mwilcL�� gI!;=^��?p������grj(C�x���%��ν���	{�ń9Mf��&� 4�M�߅O�i���jo{�-�0L���ۢ;���m�/ߪ�.�Y;(�&�)ˣ j\�����Cᇬ,׎p̖�#�Vꄖl��t��َ�(�/���� �������ї�E�}��>���"Ψߚ��wXz�s� [0����U���jr���5�8�f�>�ir�k�-�[�#-B@�����ɞ>֚<.PFPw�B�Q,�Ꞡp�)���+�������)j�.�\�y�YԦ�L�`p��B.S�I�	��7)��e������ Q��sy�Bs�9����)=�� P\߮�� ��>�@�)�����b�\$��6`���c�X�L1f6���gZc��IU�fT�����ONG�Z+U��W�lkM���^ժ���f6U��"��qN\������o:i{Y�{���z�7�+%�W�y%gg�����Dۣ��Ս��6<L�Z�����	b�y�V��B�ppp]�QLP��(�D������h] ���Qe\��p�՛ۃ����"巚R*ʴ�����ЮT���6K<��8-��"U0g�:���$�,A�rU�=� ����9�+���;����ʭ�Sj����t�{�6H����-��S���a���˸X���
��O����I_��{}]#� b�h.��~<�2�3V��C1���7�l���Z=�@|U���.Ǣs���}��Ea�f������<��˞4E$z���5�̱��J��I���?�"�~3y\�k�^�M鑠�}��wҾ�5玄1�v�_�'�/��}�;�G�tc�5�����rl�,~�'�_��*�#�/JP�Z��=�@�˶K�8�G��j-1���P��z{�T'��(�i��qVP���`ab�R'H��̟�/���?�[���U��b_��y,���,Bcsg	��k�����O-�|K�Q]�	��5p���2i;�����-��9��8 7�f�D��H;����Àտ9�
2l|/�#(�"�<����;t��x��Lž�<�J��\��+��!AJAzy�ۿ	��6ì��u����3'3;��R���aL/	�~�-�!tanfz�K����J4pX���*̐�����0!+����P��|�����Jm�<K��Zuq�S�ed{�_ �p��ʸl���+䏱����l�%��X;c�Kʎ� G�r�rj��*�^����0|�Z2�λ�4���a�XLӦrSf;w$˝8�=��l��CU�`r@j�����A�ǿh'�u�WfM������.� �m�ﰿ�ή�	�g����%<{0�x�hx��>���e>�h�$��!VIO4:#�y��_'�M�*���\V���A�p&��P�0�T<�ӲF#�8Z:$k�(�c��2B�R��1���-�I�R�2MT��L#�9�.�0���A�SС���$#(R��:.=Yp��|�6zah��Dj�j˅�8*�hI����vuAN��Б�C(����항7�	`J���o�P���ZZ!U�yu�]�ˍ~�(�?��M�y�H=����	��y�O��;���Ʊ��Vk��S��&�^Q�d�|-M���$ˎr<��L}�b�bɮ�L/]��҅&��"I	�I�ŏ�)$��r��w��t�Icj(�.�z3�Zoj�=���6��W��!��k�qc��sܪ�Q˶�{�w����b�j?'�?��M�gLv�:͍�i2I����YGf1��1Ӄi��=�\IC�E�b�����xe��ñv��cDSK���L�N˴x=q�<|Gf��\�Xa���y�:"�|�y������8��tgh=���E~�,���+�?k��W��0��-)�l<cs�_ր)��  O��_��K�Q�w}/�2�eD�c���#~���8��%q�M�,#�z(EE�xnĺ�li��sN��G�ȘFʎ�a�ћ�X�v����HLp��9��� f�D�U�l�Q'�.��a/y�c��N�7j`�S3�XV���J���v:�sv��4�s6�<Qy�+˨h��I��!��4�� ��[z&���T���Y��Ɓ���.��b� ���
p��g\�jW��
.�NTyЈDƺ�= ����<�^�Y�SG�a`��[���v��K	�b�3oww�6�YP���໹a��X�?gu�J1���i����U���y�E�Td$�ֲIF�ZN������Q�z-��G�����͙C�Z|���O嬐;�C�8c����� =n�>�6e�k�Y�9����
�[|�(�>z�W["�v�&�|������a�*.�p�h�a��;�l-x�j��vA���CU}R���-��DE���.��LNw����S��?�3r:xU�ehH��{�OS��[����t&ܖ��1���d	�|�]K٭�\\j��] �A����\O�	�N���=FƼ�J�r�35�u܍�ո�A��jfq��|,���s���S�:(i��`�M����s�ll�������U^s7gג���L��N}�l�d������@N�����0�U�j��i)�O�,�����JY��X�,�y�Ҙ���rѼs�����.T����>^����#%� ]�ԉ�K϶	�Fl��"�����Aɒ�ji���C�g��*���	���-f�Co�������}ʡ<�W�l��x�����b<���Z�H�Y�5�4�"��Qc$$�X-j#UC�����{�w��]7�a�54����Nwꖚ������5�A��Njl���gl��;i�*��_]|��*�A��V�:�+�1��Ѥ<a#5":|Z- -W �yg�W�5���0�X:� ��L}���`LS�h!{�]���ۺv�6@�-n��eP��_��;k �㬆ՠg|�E2ԇq��|�t)�J=4�4/��Dw$�Oˍ���g�	�Wc��n�Kt8��<KG,՝g�h�S��)ֈ�f`9�o1f�7S�\V�U�gA�c:�eCv�QC7���W;�!Y3�B���J��ASA9N�7���2����P�DS�����K�����G
��Og0�m�j�4�!�E'i��<8�9]\��f������x�m'���Y��v��^�)O*.I:�/�4,���(��M8�N*�c�s�6r��/)���F��Ĩ	G�E%�6�Be�1�T���V ���I%�fp~� 0pZ�j�A�p���TZ�ȝ�'
�RY!Յ|SԄG�i�y�Uie� ]�%WU�d�!�a�g�E	��q~J�������vp\���>x
7_'̍�3��)ޘ�t~Dr�,_#�o�p�ú)�8+�d�3����ܮ�&���q6�e�4���pF����%�Q�"���Z�yN嬘m�Ac&�LFw!�����#HI#V��8u���f�+]r��p��di�M�h
<��x��"tO�=9���>��y��	����4����ʫ���*WRYJ}R�`��F��W&&�Bv W�	��� l���{� k`W5��������'������T��oP }omԑ�TK��jgᶖ>�WL�hHx���[��#*�㇓��{��p~�k8�g����l#�5�F#�]%+�X�~}"E
:ʋ�����\%��]���Y�YD����P�Uuw��$̓��TW��C5�<�aP�ᣝ\��7��4IAW9_�5�=�'	v/�E��t�SW�Ž�C���d�{��,��� ����e�#��2C���q��u�}�2�@<�Ȥ}"EZ�{+�� ���&������*e&@N��S���h�e��VI�!�A�g��}k'kۓ��j@�N�'+�Q���qs��a=�O9�*�:���j��NC�V��Z!�-F��h��d#E)'���[Q�Faַ�F���A����}���Q�ll�&�c�D��JK�hzg�XO�9i�Q��V֏`�J#�S]"����"*.Bi����R��������u�ЂG�&�{?L蠀�|��������q����ס��G�?FGOl,OHҚo��nD$[~�-	���!�'/�H������q��(��r���B"pb��8�d5�gGn����1�8��\����`8�P�E�H�2���L �2������~�%2LG���qdvKg�m��P�@L�q�8r��k_p'���P$�z���I��ӫ��2��Uo�!ө����P��zh����.�%�����H~�~��tP�/hO��ѯ�NB�U.���e���g�M'�d�P� ����_2]t|�#��G_����,�����TH��G�G.3�M-�8����\�.w2�R���@N%������^�Kg�8��d�dN���=�Ę�6�6�0UW?��,����3P�Z1ٳ������0D	*�X�ҙ�,8(�+(a;c��Q��˃N�wD������?�����$�'���H�\:�<�yum��M�"�O^m����Ne~��ި���	�3�`�r����R���$8��#� L;�U�Q����Y"8�Px��N��H�-�"��NR~:�v�K;gG{�����1�XH.�������l���\Ύ�/��.֮G�b�*�<���F��m��&�ȴy�~�ݨ�����Y<��W8W%@9;_����4\|wFs��xpy9]�?+��%8wt!��BL��=��n�Wtޭ��ۀ��)��9�i�F�����X�9"a���eo�q�z:<ιx�+��:�G
˚�5�F��n�I#H��9U�I��1�T�}ۙ�wd��v��H�߱�	I�[�}|u�j+��B$��a�����o�/4�w�M.3���qW*I ��ٙ���	���y�3���;uչ��8���EvY�&I���V�ʾQ��SW�Y6�e֕�^�UƵ��0��+:����<�M�޳$�s�_�u��)���i�&�k����lיּ=R�%����R�����{F��a��_�?��a�_�������Ikb��p�{�4?�`i# Ip�Ǌ���4�Z�m��B�yiNu��	�1�Do�Ua�_�t;�y�Eςr��<���zK���Jp�T�����r�����F��yN���m��7�pU�3)Q��w��3�=L�k�36l6ox�E�2�U5!��a�Ȓ�<�\?+��u,p�B�1X��b��m��
�=8��jy�I��+�J�U����3ݲV���lL~YY0� �M�p��׀��@s�F�����	��#|e���	Ǳ5��l.�F4�W�N7�-��V�:f<F���ƀ�]�b6��ļ�����׊�h�-�{�,<�i��b}H��~���-Gh�`N�_�����Ҙ��EIw"�nxVcW<�� 0��a�l6`�b���.�E)O%�F	H� �Î�Vʡ���6_�c�x��.��t�<��*E7�Lr��� ���nޡ����i]��+-�&���t㑎���Ϗ��䭴&����z]C4S��`g����s���e]���'vz� ��̆X�D�
�@U���ԮU[
��q�{kc�~�vP�o��od	e{,��u��a�z���K�m�n���EK�V����u�Q}�6��=����U�[�(h����x�'�Sّ5K'���%��([yu���.UzM��z�!f���tT4T����`8"���!r5i���A́��3���JBzB�B�j����e�?��r�k���-����3�*�8����4�K�ʟ�'���)>�[���p�QR��܁(�w,+0�6!]����L���y�F���ƍ	5����g�0�*�蘨@҄���:V�r�*:��9�i� �>�Dn�wCB[^���Xh�h�
�[J�J`%ш�g5�}�GE��w��Jw��ԏeP����gN�P{N���sQu��,� � �=�?��>{��""�zl~_��j�F��Q"1��d���Zd�4������ٌ�8�1��9���+	�a�������٥U�G�r/�7m��V�L����و��Yhdz�'�ϵ
�l�"NbԐ��́v�g�����E��44�#�I����vm���OzO�t�ҧ��g�e�w�cG{+�3��0������o
3Im>MN��� ����,ՁC�Wr=b�
_u�E����`����o\��) @N#h�6�)毪6.2Ԏl���7mF68��+��':��T
`���$U0@�{�q��A��9����%�7ojܓ��q=J�2{�5ő!��I��	^�&��$�rf�b+�D͎��0U"�RxαN��1%�ݑ��?��W���_롛|��R���<~��!鰑t�~:!z��&�ɗ�����P�P�6��F�\��`�8¢mUi���S4*K�-[��zV�&q���^�����W9fBm�<�mϨ��pcu��@mX�C"u*��a���1M8�u��<������K�D����,
�ڗ��r�e��S5T6�r�܏�%>x���FH0���&	|9m���t�94�ǰ�_��:��_o�FS�Y�Z�^��*7~�g-c���|�@Q��[e�Fv_���X���\���,�1oIG�m''�|����5A!aF�bڑ�U>6~Е�%��{���CM���_O����i��H��TB�yC�w�Hw���w��7�P�҈)s�z_Q&Nt�6�3��p�iZ5����+������7��1ؿd��@l���}��nL�~��%�݊r�G�OΞ���%*��Ŀku��!j����c�ᾤ]U��:4���e�ߜ�y���ݻ�iR�|b88%�.��I�����#槟���(�tR�����:���c�a�gL9C����R�)�Yn�
�1��߃	઎�N��������������r{�焌?�R?,B�+N�%ǹ�x��y�v6�;r���B�g�'ʄ�NT�Rj �є�n;$T\l\����G�"q����W�]2�O�N�G'iz���Wq�B	�bIC�#�-�uPŠ2�5s�^u��@��h��y@"Kz���&���������>1�9\a���4q�;�1+�wm���hd(����z�<Փ�J�����v�UA���ER�8k�A"�#9�a���b"����!ni�@cU�K�ρ���X����:ۚ�,?��᎗t͸�H��-�穝��#w����fu��`!�t�96���/�B	��E�xEj)4Bt�
S:�
�R[z&���3g(9+@��3!	���6�ީǞ���Щ&�hlхi��)i�w����M���m6n)�J�A���MyZ�4`C��Ws�k"�wU��㙢�I���R�遚,���� ���f��֮&<)��w�.��j�1����6�� T����,�dK3�i��N6���U�����<�?U���3])���[�H�P��Z7����=�V��o��|�����*g���'x�>8�j1��b��Y`u��>���α�I3<9N�'+�<J����gA��_vT/�w�(n�h��Bgq#���*�ECb����Ԃ�y��;|����B��զx��]�Y�bcFab^y`y�ϣف0b�'�v|�A��1�P�\e���Qa�	�3˩p���'���i��cg��o}͙|�jv��1�s�Э Qbl��59ca���jD^�c�@�*J�l�K=؊F���!�,7� *���ۓ����I �cw�pK�h賉� }E���sUn�-�+�(�23����{;��-Pnb���&)����i?KP�G�wSf7��vqt��@�6�e�C���7�S[X^�l5~cI,j�Ө�v�%���D�?ڲ�?�����(p0�/������ɹ�Q�l5���f�%^�UkF�-�:�Pߍç�~w���P�ƨ,=+" �h��f$B����P���UٍJɂ/�!�F��A�����,���Ҭ�B���w�����v]Xuӌ���NE��0��Xt��6��m�|g ���
~6�볞�-S�E���ޘ�� y�Ҵ�9��$��ӕ"����]�~��]�n��U�̌c�SW! ,2�ڥ �ｇc2^q���k��Z)�N�J�U��� )��}�8OҊoD�T/���>f>|jes%�:e�����+}kN�a[�Ӝݾ�}d����\#���]�=�6�.@��Ԇ����������VM�/rfA�_9��ߢuá(�ĹRi#�Q�������R�a3y�j�Ue@��VBZ�������F��7�Aͱ.v%�4����{����V�9<��Ӫ�s ��	S�ח�w�j��p������?5ar˘w�f���e�z��h��=��؊���d�g� U��L���>��pB�A�ǔ�޸���S8�20��Ȑ�W �Y�<���(�|�/�CY��0��GT�^�)� �#ñVH9Wt�vv�đ��u����c%OUl,R4>deѕ\�<vi<�Z�Z\^�$���h�@YF��p�^c���3�)6/�Q�] IT(7�b�|!_2)��Ê;-*`�Q�H�
��ElK"��é���*�$/o�d�I�+����&><ݕ�H���Kv�K�,�W�zd����se�ΊN��;hn]��`b�Z�5ϴ3�38#��r��Œߊh�yێ�F�!��Y����^Rj�|H�rz�ZV�D���A�g��*��~࡝"��}M�c�牐����rI*
�Y\4�3Su�f��pڹѿf��g>����g�O֌n��-���Nu{�Ĩt�r1s 8�g��0.�q��W6�!�-02�����t�I��<�[�w��X�N���AW�k�}b�n�o�;5��n}N'J)���Af�����W��V���9�tK�.Q*a�)���S��S��?~S�
Aɻ�BVN�dV��ct�%6���/��K��o�k�P�j�K�HM`B6�*V�r�n��9x��Γ�����-f�x/d�
1�Hg-���b�c1(Q�zh��u�v�X�Tx��`��Wh�-]N~Vqb�)'�`�"�02Ԣ7ܹc�P��s2���,����'-6���U���#Y���X�J�L����&�S2�(r�I��W&w$�:{I�=eF��,l�I������ϖ��� �'v�k�L���]��9ݧ#�����]��*ہ�a��{�� ZX*��8e�YX��Q���a�B8�?m��0Jn�0Z��8s���;���\e�+�m���k�Ȱq�~s�0B�u��-'J[~����ZBJ�|���v������YħR��K�R��$~�;�{���{h�z�� �O�K�l.�$�p<2o^���R�9��\7$�t��ⱋ��C��A�@������_j�y)i�gp�Z��2\Yf.��D��7�能~::&ߓd�H\瑽��̷v�����F����+������N���5F)'Ӫ6�����lw�b�d鹩���?�8���ԕΰL��{p��*u��1��L�zuߍ������<�o`�B���s{���ټ0S�D�6�<]��g2�xH��%�(��9�E�(�����M*�
E���G��ۄU�Q��Ғ)i���/���/�`��}X�疞��
fC����Q�>r��>Z�B�D��J3�r�덬��_/\����SR�P���1T;ъ���1J_"p�,�X� �NF��"�#���4����w��f�S�Pƛ�X8q��=���X$w���;��L68��~��-e�Јm)"�Q��|W��f�̨c|�d%bm]��<����Cğ�3�h���]��+�ܦ��HI>�%%C�V�^�U���m��n<��֍5Q���'�S�$�D���!Ko/��[�:��g`* �^�y��`g������;A=�F�(��aѬ���etl]�
Rp��d׀5�����֌�Ϊc5�ƭ�����q�~������K��+9ЃH�+V�U�"�O�� ��?(��'�j�.F�q��T�43x(ᵀ��l�V���`i�Z+��,�p�\-�2v���Df086a_嵝g=�H,�5��� ]�Lq��:��w�2�u�S=���`]K �/r���Ӏ/�W�.�T2�Mp�>pI���[g�nj�]����>�Vb@薛H)���M�X�ݓ�_���@mҽ"�v�e�&YD����m>��Pr'��\���������D���uz��5��2�)�n�c�_�L�G�-{)����z���N}+��:���8�p��K��X= �.��`#,
4hF1PvT��я��j ��$�m����X�E��1v�sjVה�J<G�=;�N�`�V+����]X@^r�/M��H���2�h�8��ہ𢁲�U|�&j!���ܡi�,j=�k����P�ÜH6�8�uO���5N2X��(֜pK-e�)�a����D�ŕ��Zߴ�£��u(�]�D��ȩ�ά�9�1��i��/dw0q60}^:m��\(�?�^�٪Q�t_+2c�V�Ŋ[@>|�O�P�J0��Ek\��>.��՟�J}��þ0;�0�=��e���Wt���n���,r�n09j�Z9(�@�'�+#mn]Κ=5}y ]�?����ӗB��B�J�j�"�g��n�H���3�p����J��Π>B�#����]A`�y�Rl��U �"[G��a I� �L�D�;c��F$�|�f����EvL���WeM����[*���@�]Q��9v�[�2�r�K�us/�=*_% ��C��c�i�fL��}\@��I�5�ec{�j&4�M�+�&+ma^'�
��,dv�	�N̅��X����ױ�ȲdD�v�3-�},�2M;��:L���EnKM����~ʾ��~�0�[�Z+�Z����p'�,��%����]f��7Y�Aΰ�f0SQ?��b^��a K��9�60��J"�S(�ER�<}ޏ�-��{��x�~4�i79����-j,z�Qd|(6BR��@�����f1�p�_�
��a΍�pVU�7�j�I��[�{8�8�M���)kV��D/���o�Z�de#��AQu,�K���k�Oçg��g@"� ��x�v�{�未��
�uf��a��-79F_���܅�03���"w&��4�F�x�����)Z�����M'#y�NN��2��M��;�W��^�p��&��RYu�5	-�d�a5)v3��xD���/O#��+��,Y *OQG�������)�T=ɖ$u�b 	�
j0.�N	Giφ$��׵�������'%Y[vu��5X�Ko"Gs�uk�4��e�j���Ȝ�+��LsB��3��A�h���b�7/��[8֌^�e�����}]�)�1���#�4ZV�8,O�Ы�!���+�����򥼞z�ʓ��E�	�����?a�8�3?P�La;�f�gneGԬ��U]�ŏh�ig�T�&�.�6��O]��0�d���ĉ��"�+G���ܫ�@���sm)�i੍pe�p��y,83�=�K��b���BV_`�_���[dyd�d�$d�(��x�,��|`�:�{���iԓ����MW��&���P4����l�Om�(�������}CЇ�R����E4K��XP2c��H1T��� � 2���5T62{h��Oo#$xY�9�0�DwDM�T䝬�L�HH1���J�[:��5CO����ק���e����e�V̈���F�;�{@ik�1��.B��*.����	kiI��W��&K�"��hS�o!t�.~SG���ֲď���gҼ(�zЀzqx�$k����b�M�n�k�BI�=R�*f�[/5mI��1z0z�S����qM��R\�Z�A���d7�>^���Z2�h:��l�s?������@���+�
ј3���$΁Le��I���s֎��c�W�����Bwq�>
Ҏ��hC�f�4�X�����Yf�
HV�F�nd���YG�
 l��S '���܎\b�y�����$0�\�L�i3���_𨷏�߀��t��74YF��e��(����b*a�7�]����;���P�
{-p�h��j��ja���#;+��cz��"�nn��j?�1�qU3���P����x]
���#{l�F�4��_�����mie@�yQ^�P�J�4<hn�ˊ��^��!�{;����X
2:���:�+�t��Mo��Fu������:3��"M��2n+Q�2���A*��_2�@��h?���h����w�O�3y�5q�;���4 �'Ŗ�
�F�dM��8����E&�Nl�ƒ7�|e�B��]
U��z�\����R;�Q=i̬�{�a��mz��6j	�8��^�u&o�:3E9"t��=�|�C�`���;�zǨ����q���=��AǇ���0�ŀ�`�.R���*��x�g���M�`����~�h�����W.Z�R��빡�(�/�F*|���h_��l�����x���R�"���%�� �mjħ�ō��`�7pih�iQ�˷Q�$���I�n
X���x�U�({5T2�%�uB�|��E��߷�����ya�˖8��v�(�	�o$r�N���_%�����>A���{aD5Kn@a��u���X���g6%�`�W8�P?�`1�:�Aj{˚�z�l$�L�F��m�t�}�-��3��Sm�9��|~���O���4,s�y�M1ª�`R��l0m,��<��ֲ����� ]R(�S�iܣ��0) ru�F��'�7Ik��B���� G{�&��F�O�{�����+�c��U��I-��H�_#��Ha%	��v��}۸l3��Q'_���ly+�<�
FG�D��*�w1&ns���솩����JHǱ������'�������6���kڔ�P���<��C�A�KÑ�t �]�����D�(s�P���j^��Z��jktت�].��L��Ő�\�тb��G����ո�S��F@*B@�7�<���$���b�)*U��f+�`B3N�õ��̧�W�ו(�?	K���j�R�e�ef�>�IW��;3��F�@Y�~=T����������D�Jڧ#�qـ�'��95Cɿ܍|�̟/�~�`#�� ]��N8V�[#d�
}e�raެ~j:��p����.?q6z����@�A�6
;�R��"�?��>T`ɋl+O������`�ˮWV��Qv+ʉ� �֠����;�D]���o�nD�e:[^7/�TH!I�հ�%�x��_IY[�1d5F���ym\53X,*���B��\w��Hos����,f�%r���>���eҀu�6��&~J�+4j�����a�o��H�i\��ɴ��%Z���T�[�������]���DBV}t��lb���X;�_��裔J&��w�T��]�eQ� ��Kzا��y�Hc���(�̻��8�>�?V��wZ�����˃[%��ӗ�&ѬV]Q�s��H($���m�i��v��(�]�~�1J�mF�i��t��
#�2�oi\c�zVD`�����ύt�^����H�壣�#w�c1���*��7�W��w���x7n��5��2�!�u����%`VVb�⒬�#��,��z��+93��8�x��_H���p��W��I��౮[�9����
�ky&2ޚw�#��D#�)�[��50c]W�#ǅ�ai��A�$��,V����߁�gv��z㳧�J.gB�(@�� VҦ��B��P(H�~ӇX��B�N�'k}1�$R%`?���'��P�Ī��7��x�u�%�#^�E�PP%:������?v1h�+��<�&�XW���UK��<WȸHgء�gwpMO��i?�9����3!�N/A��+l�5�Iy�y������������4�@���w�۪�	�2U�G9 �+�޲ںP�Iֵ���
�p��+¨}0���6Jy���7yE�L�w��A��2�D�U`��6�������^()�h!��V-����������\��/NԜÏT���R/߸K���Ŀ���Ҏx#���1r�&<u;�.�_�,Jւ1�ȵ&
� f	��c!��׬:o�␋�L�C���so���Ђ�˹�h����=<�WÂGۊ�����������b,Sg���+]��D�z�x��������fG�&6Sg�<����
��etz�����<�*�nI��BD9�Vd ��T.�Uj��_���ĝĞ�7l���Y�W��nV����H�E׫&`$K'����a�N���k� ]�s���.�]������p��
��y�0X䁦�,2�Zv���^0�5������|H�:�U����_?hR�qAb�����rr?8#�ٱ�t~���rEv�M ���d�P�[�7`��7U��,��9��� ���C��1o^�����q�A@9ژ$%,bYN� �@w����*�����iL�_*��$y]C��w�:gj�����ӈD@�/�>�92NK�OC\���Q�����~#���q���h�`�ޒ���=S��aj�i��ս�&{�_[���>u�nd�]�k�!Z<��v*m�����q[�)���2�:�eJ�ʨ�	�͢׊�;'^"��H�C����sI�]��}�U��͈i�v&t%5Q/�/��ԏl�Lh\ǹNgM��@���wd�VW#1��R�#�.��ě�,]�ct�{�$;�Ǒ��͏���T�P?w�����:`+o���!�R������O �&̠4��K0�H=v'���K�&�"t'�X�[���I���ikS�\�5.I���֟���ƿ������K��y`5���J��&f�/��R�b���!��Pӈ�$`�� )<�y�i�F�Nm�kG��U /�֭�B3b���"+�o��P���sf�}����ž��(ds}�/͍'��_��ȯ$�9 ��8o�KA6���fo����iLX���M<b��x��W&�M���+�YD(��<�3��<�
6�z�S���R�T�rH�[��Q�$L�vw%YM|nj�<�Ae^Q8|<D�K�3�����~(tƼq���g�"wk���?j3&�÷j1��΋.��{CՉ��;��j~�nL��i�|g�sZ�����u%�S)4~��QC.��CZ	J���X�/�T�_񁱬3g�9Ii�f��-c���@��+�g��1kjm����pˣ�k+kSs|P�V��ʅ���=_�'��e4�Fj�߳=�`�>N�{��!�;�+i.؉�e!���{�Hf��f��%Vsn�Z�6��g�=��Ԋ'���=�H��O׾�*;Ή7�	�@_�^���g_-e�����ͤ_Q�ViSai*�]}��_ϹD+��mU*���<�?�ׄg�W�ϼ�/�B��[?ʴoO��I��$4���\�'�{h5{�B �4�U�����R��(8�1��G�PB�C�aw�`W|�*��R� �J���x!�ai����.�`2�3V��7�-"�p���߿��?m���n���ݷ��C�`&(��Z�\��(����Z�k�3�`����Яk�PA�-���+�-��ẘ*��~϶p�	.a��SPb�B[t3t�/]ް�/f���i���C�}T5)� ,D m�νg?�bz���nTG�v�A�/�gi-�R�ɿB�0śa[y��������]S�'y�~����t�U� ����NT!2��>���]���>)��s�g��&GӸ[� t�蕽+ii�i㛛:kJk|H���c�eǻ3�;Wn��7z�_��6�|Ѓ�^(qÒ��և2Z��2Z�u�퟽#v��&�gT'C���Uw�
rהL�~k��7�����eû��n�����c?kO
C��Ĩ����X%\r;�|�/S����nF)rB�v
��ƽe0/$䬇n$(l�߻�'}C�~�>t���x�߫̈]c�S@�Զ�������G`9�+v�};T��%53-��Wґ[�j��T~[�6J��Əu^��v��퀝�^H��U�#YcD�o� �[�{��Ȭ��5��i�v3�rk
�F����ԡ����s���ij#�vkJ�W$YxO�{z�x➂f��tf�E���+Z�c֪Ŋc9��	�;��#P��q�{�%9*��w��YvF�~���UZ0��3�w?�A��z�9��RU.�E(̦"�i���{x��Y��Ql5��튲��+e���A�6�
��`2@8<�6n%��Q��D��󴱉kY�I'�=��#CV��9�l6��I�9l&4�'�O��:�jLD��'����<���L���p4N�@Iȗo�-�.*�%�"�ga��V�TV������������J��q�+�]@�+��CC{
��oB";8,,8��x��(�4�������)� ���v�^ V 2�Y�%<hpF�EN��_��G����B�\�qUV���3#U���U֛3��W��eR�Th-绎HŮ2�Z�P�V���k��lo#K�?֓��e*�a�}g$d����6�s�ΐCLv��`���I�$�$j���c�ԧe
�Tފ��*�\��,JE�]�Ґ� �}ِ�V�Y֏�� �d�6���������\�o�����6	�X$'�D�,sRd��z�!҉
j�ݾ�K&.~�_�kÁ7k�I���P�^-�)��:�|�R5�b�a�_��be���6s�+w��_�_��?�(�HG�x͆�"�f��^"������L^o��I+�i+@֥�T��T�	�WI�F7[�Y+}�D��aIT�� ��D��38L�nitІ뜬7�F*����hh���'#	�[g���Ivs&����ahQ��p[���٧����jG��v0� 'P�h���v�²�&���s:�����)�H��`��©���`���;��B�.�n/g�j�c�%�>p�)]�1�EA�ޯ��E)��,�k�@q`�� ��3����a�q�=�^%�y�])�I*۟�O|7�m�T\N"��������Del�(�-�]�`��0[���V����78v��o�U��
�̴�^��߁c;������fh�қ[�P��AX�?����>o�����h�0��?�5����ɥ.����G�׮�vW������+��أ���~�vV�����O~�Aυ�XМT�<������ )5��M�Q��7�H�U;�.ܳTO���Y����p�ڶ^�ʫ�ql�����,�� Z���܃�=SRc��\2}5�bXz_��T� >^��g��G|zT�n*e�7BeuD��"PC�U8z�HNQp�|V 0e~�J�%v�e��Z,�/A��!���%�/$��@%�D-�]x��j'�=�������H�����C~�d�e��u�"�W
����<f�c������L,c��y��#E,���#�@�Ϩ٫��J�oo�Gq����2J�q��D?���q�y�{��F��TH�|�GI$�;լw��������[��&�v~�hȎ�s������^��	�ĂAb�n�d���ő���w���гG�9�� -8p�5���Fk4�4�\��q�9�W觲��ܶ��3��K�ky�\�z���b�.������$�������KA.��
14TV���N0��K����O�������^K{@���|�o�X�į�cG#�5��$P�?�6�Ԩ? �4AfG��5bÖ?3�.�k���pPL-a��@�[�}���$`���׮�ح�yO�d�(^���"���ze�ٲM̆���ʺ�R[\��CQV\�I!(dsޚ�{6���|*Uj���t��uf��P�8<���������@�^����j��p�G�SmUʡ˸\�������Y,D�'���N�2:R见�a�
��{�&����m��ֺC�itX^|bi�%wO�ZH���X� B��z}Q��A�a�#�ϐ�O%Y����(��U�8#���@���(�>�ׇ%C�}N�:J��kav��g�r���c.�}���L���9�����I�Ɍ�?e �5M<����]#{Wo`��ڇ~b*���2������9��9�h���X�V��VX[򛙜��'G�^u�~�e����4W&ciDj�_R<�S-~!��P;��;?���X��`���Ur�I����ϖV����K`��^6��J�F�z���m�(1`�+�]٦#&l�1�����d9�|�/w�1iV�W;	;J��|�0X�J�[h�ɼp����1eR��gQ�����.�F���3@1��,���=���F������[�)�������b�cC͇����f���_�G���K:�UiU^`�&s�M��D���˃tt~q��u����iҩ��J|d��oa���G=G|s.x,+0LJ~��bR&C��&J��aJZ����fbm���o��g��e��JI���2!��V������y�rL1n���$Ftu�侺���-r�pi|�q���FH�\�e������6��4x�A��wkOt���w.�����[旻�f��i|�7a����)}3�>�Ƙ�ܪ.v㼞�jЧ�0�3 ��$ں���U���W�e|8�ߒ��+�p{��'�Geм9ר��o�]�H�4sO�����q���0	IY]�R�?�?�#c/4�sڲz+pQ�o�w4dڂ�Z�u<AL�_��BFEi
��"�sE���������ג.}����3�:���S(�>�S��'//�)*\��iw��4���O��K�E&�h[
h[���f)���i���+���	�z��T�a�m����(r�k�!��a
o�@R���/.�C$���H����Q���Ig[i$#䠇�N������Мʲaky��[�+�̘�f��ʒ[~�'	�Ka��R0-rs�
��v��|^u�y���0o��`�:J{SR�IZ���-���y���3&���&����LI���Hs���`f�nK2��k�s颾��8*�~�ш��<��M�Q6���,< �4�M�`L����O�^n���1y���R�.���x�Q�w���1כxda{�'�h��]�����n���\ m�7��]TX�4[ݕ�A�Z{��so:���i奛 ����ǜ,��ŝw�6	��e�|M�vv��6�~ws/J����2�IM���=f��6ɘ�C~Q��'�T{šPT���C�����\()7�����|�岥��0L��2�\�rǜ�%���-�w|��!�q�IJј⾢u1����:Q+���K�PϟG5���ɯgA����\,�i�O }m��#�]�_���:�����ְi�b�fo�˛#ѿ�2�?k�/@䡭ܷ�D���<��klY�Σ�����%K��F����vI�!h��I`��l�Z�Ӥ'3O�;! ��1}��1W�=UVs����I��<[��ʍ_�e\LR����"WI�n)����%����2]�� z����a#�����ϫ��$�26�
���j��MjA�c�qe��K�`4E�|�c�~ʠR�/�jvN���-�����!���Ö�k�
`��@����w��a鸙�,r~f���ff�V����"kK��fJ�ժ�F�S�������� �\���1րW��ۨKN���t\�̤��'�΅EA���{-���=��t���NE��.�H�/+J,�ƚ��yW=U���2/��Zp��~z���݌;:��I7�S�}��'Roe���(�%���FL6��9m��S��M�uQ�ϒ�Ҳ���kC ��6�C�x����lU�Je����sC-&��Y�&��F�+5�ƴ������,� X���:�Gt��H��}(K�����Mw���r�le�d��@W�_R!
`�NY�R����vΆ|��^>��~�m���XJ�o�h`�8eP�9�kNk�j}_���D��BV�L�tˏ5/v��+�a�R�=�kS����3��<�W�u�fV>&��7�_����X<�@�J���[�������۱|Ó��A������h���|@aR�|Q�_{n�+#��`h��wԹ��]̫�VF}��I�%�g�<G"��8��>J.�+��b���`��4��H����F]3�u��'�������] S��͓␋
�># �8+Ut#��
0o&v��k�̘΁��Vx�9�P^���S����l6���.�Zֿ~Vm<8G&,&)p�E�uI\=�z��k����У�>��kV7p�I�D��p��-��esQZ,G�$d��u��1e����c�R�ݟ��*3Pꍂ�߄R�g�n�d�$fjP`�r��˟yq�R闖㳳
͆SE�*�Ԫ_�Zh}hs ��7O���"7ܞ��ƌ���m��t�9�x7?�?��؟D�G&���-�ا�Q��'����!�ŋ���e�;hz�*�a���	��s��q�7�mb��C�cJ��ۘ<v�]��c�>��Y[�x���������~`������2�Ŝ����=Oƹr�Qk�nV�H���b�li���Y�k��J�ξ܋�2�<i�m�v�_B���J�����I�����f�DI�587Q&��a0�G�&sE"}��*��¿����Ƌ��B�a*�Bf*�<�T��˚IF��	�� �]�����{���<�Y��e�X�y�?�]�F�&Ua6�-+�Vw��3�%��S'�)0��'UP=��Qug$�C55eܬ��3]`�R`�H�f��уPF(Y�D���C�O'���+U�萱4��8�&�&q$��5~����V#��"�ZX9����g�L(I�$�\�;;�������D���$��s�	�py�揬�`�S��)���b'{��1+��!��W��I��\bg�W�"��@dt��y����|)�!=�G�	�]Pu*J�Wҍ?e��-����tg��S	�4���ɯ��fA�z�8�[./��	��Nꝸ1^����X �wV6-5V1��+#-���B|˚����p�"�*���AlR|��

�_9=����o&���`��vaɧ:AU��.���N�x��F[���� 筆����D=^bF,�������n���3-{V� n�7}��H����܃�ֵ@B�j]֒��#�a޵EVt;�⾣Qg��6u&�H�\Zn͈�:�QeK� ��<棱�xz���+�j|�������k1�?M��G9��Ʋd���'� _:��y5A8-����֚Uw,��G�81n(��A��D��q��,Q���Հ>\����	���y�:��X�����dt�M�[�6
�+;[w7�ޱ��W�J:��������S�{���A�[8����� +vw�XM�y�V�"�d�0@b�R�,�����;P�ΐ^���>�O��͝�[�o�˪Jsx��^v:DR�G~���C�iRs���fz���V��z!����(��}u^�G��\�6��3�Dj�#\T97e�,�]cgq"�?������X���R'Aw�a$�:�P�|��:o#�ik,+t����*϶��=��:sA�1��l-��&���b�]��l#��x	��s�M�\�����y�ᴄ^���,�/9CA!r�XB�B��Ь���w�y�enZ���)����u�؝���|�5��M7)�k��м4����F�>��}�@�C���ň�M�1�RT\a`�
y�N�5���笏����L@�\�N� �����K�֭:!�z�oo�V���ME�����&c���֌��f���E�7,�n�Q��Sq8�������Џ�������93������H�SEQ.��˛��p�h)�Jخf<�+�9��V\^�LzY�9�����Bn��r]�+韷Ds�J��Q:dRT>i��#]#��i���~_�T�T�b0�H�@�IQ�3|��O�fb�?��j9�M;�ݨp�G��N��M.��`�K��������U����>��>�ss���Џx�nZ(�����`w`���}ȥŪ����P(�'I5�S���/�V�<݀NV�+R�%G�z�+�m��u6:�̰_Sn"-Ƣ	F�}o8S�~�;ٖF��>�ۜ�j7*�w4��k�:�܊=̪ZE��'$��(V�}-�|wĎe̲Z���E˙:)n�^ϸ[I{j�u;�f'z���h٧�M��@�뼽��M�!�M\�䃀���m��%q���Z̈��N���:H��-��;��>��ȡ�nΖS�-.��?�����D��1��$��<2��M��d{k�.g3��i�	�
�Ȯi��r?f�O|��%ۧ�HN�R� °zݼ�`h����=����g�	��І>J�dE8\���-	�'3�?.������S��vg�������$Z3�V�� iZ�HC�z�2ٰ�t���v��$$�=�@�/��o&/Sh�%{*��:ɝ"Ā���*2&w!/.��J�B��Z��C�D}�Q;LU��Qt��Q��ti�����o ���miTSk"�$���_�r�/���f�>ݍh��0S��7��dX?"�m��C�M2	FO(8w�P�m��6���0���J��� ��T}��Y��K�H�`
��(HbDM�ai�Sn��R���iL3; �D�@6IOl)0hG@РY�p�QW�۫�m�$�Aj��r�мf�,:�>F�}��i��*7R�B4��1������`���­r9)�6�L�)�����p�G��K��w8��߉=N�H��E�����7)`�*"�ׂu�o_&��^òTXP�s4��ZF}w��7�͐JIK'�ٗ0���m����H�u2���vRg�z��C^J�i���3���E*��{r�n���"7���jj'љ2Wڧ�?��'�����1w��
�-E����0����+<R���^2R!���PK����e�(�>[�4X�ƇK֚T�P�^JKp�����䅜~��3ߑ�-HQ�����5�[�����Op�S���:q�:4
n�d�y��g�e曦F:C*w�q��hY�Fۄ�����28������W1�B�K�r��t�歗�ue����^�}���^��ށS�`�u�
�dq�͊��y��Ë�Q1!"^@ŀ!>��N\J$ܜ�o!"�d'.��Q�#`K�H�'���2���سj:��e-=?�&��{����̬�%O3Cn�Vn�^���̩����:@���L^���d�x00"�5�]��W��8��0�q6~�GoC��~�������l*��3�J1]�g���E���cH# �?�<�i��6`��Q��_���er%�Q���(�kC$��h6�,3R#�y��BH��V�Պ���M�*��=�c��j�R�H�;G{�K<�<�~�n�\91�C#�i�??oȑt��D�r����A��*q�c�Yu�5�&R�M�uy<�j�����߉S����N!�L����#�f�⃀1e�ذ��wqa� �f#�#/N"�bE�{�,e�G���a^WK]�i[�A<��dwjmǎ��N�*�q#r��[�ő�icJhu_Z��+�*=���o~Y4�>����\pٮc<%��x�B/�d���G"��&�v���)V������9Ǜʵ�7n�q�O����+��V�07�8�vO�(r�(]1'��QD$���c�!ڭ#��o�w-�v,�f���_d�5Iþw��Zĭ���*{��W�/�_KY�G��FW����b0���VC��b����#h5�}�nK��4�A$$cc��j��\�F�1sSL��:f�e o�T���?k_��T^�?΄���r&8�yV�k������ܹ	���W�x{&�;ر٬az������T/U���$ة稪�_�MF̑�v��,�@��kh���i�:Y~���;V��.��ɂ�}%7����� ��O�`^��O�:�|�+}<���`� H��It��{�g �h⑰�q4̲����ީ���@3��~|lL��@���~�J�s�|\ԽD}z抄
���,��
��R֧�"%}6RZ+�36ʫ:�y����\�����O����-w��́�ϩ�ڸZ�FZ~�: n]�U�rw�%#�2��,5�2��jL(�c�ѾD���SdyND�J!fS;�-��3�P����H��w��$:����퀛���Ƒ�qbj'o?�e3�xB���S��=�
/xXk��s>JNoܞ0i�����yc�^���ђ�@^�A��~�z�um:�Dֿ�^;�$������?ۧ��Չ(w��h�iX��&V=��FA
�?c�r�A�W=�7����{��z�c�r�O�� H�d�,C35'S�j�p�${I�yc$$���I���	Uf֪�O&��(Scg�Z?*�")�<#����F��o�~2�BJ�6$;[DD���>^�;��d��hH�0e�D/�W뜥6�Oѝ0}�JT!�h�P]ʋR��,�vb�3�JSa�'�/c�w���?.����� ��@�n�X��Q5����\���:�+	�qm���p�d������X#J�9q*����Oƛ�����TE��B�x�L�[�b��s�z` �`8�e¦ڬX�W�t%bҬ�ZM=�M-~��4ON����E/ �#-�{]_ci�B�]*n�Le���YM���4t����m_�E�ԋv�0i㬁YHG� !�IY�*��x\1�����~��p�W�{�rkߋ��߅ozSu�0eJ���,�\I�Ok�cS�.�eة�	����PY��y\5+��H�H�'Go�:��dAr�\�c'E��Gz�:~��s�C2�Jnt7�ܤc!�
g����Xv/6�,A��O�"����#����)������?�W*H͆	�!�G�`h�
��0��Ma,���q;^�}�_���`(�Q؝��4��G�^���=X^�Q�*sÏ����Rm�e�j�fX�aǰ!v�ʟ�S��E8ܙ[	��t��trn���{3�L<В���Up��+�rj��'GUa�T��#	��b��]m!����h�+/W����8�[(�,��s�i'F
���$��hݿeHK�G]��E�K�IM]���(��#,��9��`�F���=d0��Y�g�%�����J'T`���ޠqo�����up�3��q 4�_�o'� �7�F�c�k��q4����}����F�2jb*����?l�ӌ�M��$x�z�hKR��+#B4�𷯻�����G'��I�;�=�rG}��RZ�l�oJm�򑁪HG+��-�tz��z��^k��-�C�j,�J	 �$�_�o�� @�Y)�g�1���<�oɅ>�&lVy
�<���̥�[w���	V����G�?V���Z~rPLk%?5��<j"t1���,5����=�՟�1`�qr2	u��zN��MS�y�cm�B���!��q��Q���h4�����#� ��ӭw�[�a
�f�!�S%��-�h=/��{=��T�������3,�^���(<����Oj&+��NlZ�e��Xv=��Js��;7M�b�}��&d���8e��z��Cw���w���'�%imP��N|��:cb?h��L��/���4�_y�YFX�����I��ɯ�U��U5w��@�EK�/]'v]�]��/s��*�q�57���~G���K��f�'/��7W�!t�t�y�����Jf.s�q�:}5['��և&�|1�l>\T��ר�	[����������_�SNd�i>�U6p5��D�C81�6䘰���^�Ϥ�)j��$�6�q��'�<�>ik��G�@Q�����l������s1p�Y��w9���2`H:?�QxyyXe�3/f���R�V��:���sY��������dU�����dpu�&!+@tF���6��(���픉�4""�5�:�~�\���۲���K���?$Ja9Cר�6�?�$���B��l�QZn�4͉j0Ip��@ZD�[��i�fT���C��?��l7�9Q�^@=wk����|�ف�#����jQ�%��B�4�rѨ���"ȿ~�~5�X�L�^V�E��ry��p+����X��AT���S�����C�����k�q��9�j�o^�ki�\![y��P�[��Օ+G���R6��q���,ƌ�;~��'fKS�M�|�$g���N�N�j�$}	[��f.aO��@��yA}Z��Xc��b�}��W>�ps�}�x�����/���U۽��9~d�hڭ�R���F���*g	P������bD1�IH8Sjd�nl{�b����5�C%qa!P�=g���5��ڣ���%j(`Щ�"��R�%q�g�P�)l���a�+ƃo#�ݸK?m�U[�U�����x��I��9�]�>ǭ������.P��)(��;i<����&��ʆ4�٪��=�֍��X+!�ss�ۻ��|T����5��ֈ'}L�
�Wz0� �mb?��<{vU�M��ԙ=e ���r�b��\h��0{_�{f^<��O����~�4A�FJ)��ؾg�>`��>D\�ż��6�b m�L�y�����!��X�_��g+)��w���P�I��)Ͼ�VT�am����K5� �n�/�D_��Ŭ�f��٥`�X�@b$���*����� ~Qi���g�����~��+E�4$������S�a�b`�\Sb'�����[�Qt����ѾK�f�Z���=��+�*��n��������5�N��D�ݟ^
S*�/�[l�.5|G��|�Gq��	�Ա���4���s?�Y{����Qz�A}r����a\���ͺ)Tb�j;?�8�:�nԦm�᳙���o����U��
�B���]7�9�F�o�h�|Jo�h��,�d��~���[ï�ܨ���}|#��'��Ջq�S_�Ga�����$�&zaN���ʜf�)��@<��Z
<X���ş)|'w8��ϼy���s\�^��JB6s���nl��>�S���%��v�Q]�[�yj��կ�'���P�mr�2R��H�1�zI���9�U�IS�r�j���W�w�1�{�\�2�N�*�)q>�o�#2�S��зw@�[����FS���6tk�9D�i�c�9��t`.¬HI� Ƃ}�~P��$�0��WBT����p�٥�%~2�f%�.�JX��o��j_W=��.|�"�۵W����<������q3%ߝ��ٽ�����W����O���O[�UJ���?�Ɠxv�Yn��+�6��L������:>MH���ṛ�[�u�w�&W�G���ם��P���B��}��6���wn��ǻ@�@vCv�����hK�L����S����J�\�}&��d�D���$1��8���vl�!��&oq�P
Z�E7l����ӵ�4��|��'e���p�&erqӀ���/�nH�RU����<���ϝ��0n�J���T�p��Sl���aE%�ES�n��Go���(� D'�g�wN#W1a�&�u�#�G������1���ރ��S�y��eX1 Uç@%A�r��w(@Jk��G��{Q�'��z�an|8�5��G���(6H�E��g+��~���vJ��xrE��ʿ��D9|V4 �^,1ǼP��i�i:5�>&���\Yz����?hdBw�Q���;�h
��%fUOZE�����}<~1ɀ|����B5F�v��n�v�=�]�)x�;)�7Q}-�'�3)�2����ΖI.�!�pL�@^Ib��;����4x:I��6�7ul7x3���ոio錦4��*�t�4����6���a�4�c�����.W��[��ojJ�UD�yQHLvs�Uf��7������
�VdT����o[�֗n�k�t�B�x��ӑޑ�������L��,E�V!�:�|�o�%sw�X�?GKU��w��