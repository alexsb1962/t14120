��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~�J@#,�Z!��4�Um(m���7,9��c:!S?��1t�Ћb2R��9h*Vկ� �h(*L\VU�� &S��=�����SX�s�3(��[��pe6b]��CO~�\�B�����y1��P�,O ��n��Ϲ�ܡ�dNе�ul�ū~.ʣ� t�����#S����b�

���}��9tF���| <����5t=#wQ8	��7��m�llt�}5�s�Bϲ�K�%�K�a���~�Z��N�C����&rYp���g��,�|����@�g3
�A<M�(|�S��0e�@�f��@3R��/�ޘ���Rf��=��A;����״(��tr���6[���H\�S��@�i�HQh�"����᪣(���/VG���Ov^�Z�.E�ə	�~�ugEӠ����m�-p���8-�d�hz��[��hvG��ݫI�jgK�t�������2b��p:���Wnt�{� �g�W�`v�c������˩ki�&Ua=�������"�"b���ަ�M�rs�8rbm(<�����~5�9jh{D/�2��Q���aX�,ЃB�;�@Ag�R������� X��>.< ��G�)���|�H_5��w`JK����T�aJ�Z��Wi�#�0%ۜ.��P����,2�L�/����B��hi���9�Z�EUE�{��z��捜i�ɐ�f�g�i�N^����He+A�tT�>�7d�F����<�~(��ǌ�t�}5t��q�;փ����rJ��/�-�3zp�"�7^./l���(Ѵ�K-�NY!�';c�_�����=��k����?���|N�#����4(��x	��~KR����s�;�&�v+k��&4�'�JU5�C^�ލ���X�d�;��d��'s���$�D�S�=8\=sa A{���Yr�O�uc�W�z�)����t�����{ ����]�|.Z=*�}�ݭ}�#i� �<�JZߥ��Vx@?�����#H�����Õ�tn�@�ˡ��m�%�"�F0"���z����Bۊ����C[R��k��g��j��0s;��I�Z���1����
p3<�����:�N�5����iΧO�Һz�;�<2T��$P/�VFM���0�]���]����h	���z]~�3�������c����O�T�v{P%�j��U���b��:@��cH��{��I�C�Q�G����#-՗C;�ӄH�|�8�����1�� ���`#C��e\�=���!�E���a�Ǹ�|5x"����X�$J���p�Ʒ�'7o��� H,nH'�Dʢ&�@����\�8�%v�pEU!GtV�^
HYr]��]IV���9�R�����-	�?��Z�?�@qE�&�Bj�G�UG?m��e˅�� �M��ɓXex�3 Ai�{�&��ݎ���w�ʑŮ�f'�w�Τ��f�����y7
J��KE����i1���h�!��¯/�"�������Y7Ѐ��:��v�K�8^��,�]�nt��6����ъv2@�ѧzr�G�����A!�0��n�t|c�PX���7<��P��i
fe^���9O�N�+���z�Wz�!� >�l�2���sם��XS3'��\�Ml/	�֛#*��R@�$�H0�8u�K+�j�az�J�> �Mb��ǷM%B3g���K��(��;̙e! �^���̿��Q�A���խ{�/�8GG���0��K*9A0�{���1���F�:����ca|�|���,4қ�O2���?+�'&6�ҧԟ�����!�fⴌTu�(^&-T���3��J՗��Ǖ��҅h��RJ�v�=��?*��=�h������?����s�v������Z5��t�7s��`F�P�]p�+؅���siʬJ�nܪ�T�M�#olz�<�����4���h%�%?�!�S�]X�c���yf��g4�u8wM⺈Ț5�MO%�v��t/S���Wa<B�.K��7�A�L)Gl�Q�E�dZ�2pj�=2Ǘs�s_��]��e��x���>�l��?k����`p�)�,N P�,�2����I5�SDyB;"fZ�ASCH+?�q㌇�>��_Z�+:��ȁ��宔"�R�Nl
D2S�҃�<���O�_�2��Mw�m�j�+2������z����y����#|"�V�����)�������TS���(l���2��/<��b�0(P�@Vu�.#��7~j�?�%R�� �[�'�{���M������~�D�Q�[Q4�}lܺ�����͈��E��̒
��V�:�8�!��b;"�F�߄���R�ٯО���1 �"��]�*��Vٗ���;�'.H������?�7Ϊ�3t�<�]�yPHCDo�4;����o�!釬��UhC�B�����X����)���Ѷx�qީ4h<�q�G���o�t�w)����+�4�y��ԣ��J��%L�Ķl�MT�j��rS����FmH`��`�,�/��u�	�N�p�"шk4FM��}$��  �L�3nB�UL\�$Ⓐfʧ�!�M���#�q�c����܎���Q��a+��$XT,��+8��h|�u��L�E ?�~.r�]�LL�0�Y�6�wtuvc��������kD�P���>F>݉l�fPZ���� 5I�c&��PQ���}~��=�QU\c!'m����5��e���v��pa�L�Sn"	[''&'�o��J�Ma����Y��h;T))�����8ꈈO�Ҿ3��<
u��}��cnOR{_��G�����sB�-�L'6t�)*��R���Kό��ʣ�8�i�ɭ�>�z���Vm5UJ�B䎠��.LŢ������V�ť�\2�C �g�˳�|I>V�;	�Q�x�yC���Ǖ��ߋ��>^U��Y�5�����gO�P�>�7�О{0� zjU��{�_Y�7kaf9=|�(	v0�O3��5�z0H0q�0s�$Q�P}�|�:��-�7Ī�Kj��Va
 #� U�U�6�\�Z������j�e��ibȏc������%�l�{c,��2�!��[9h�t^�y�S��m3{�h�o���]��8h�Я��@�]�S<$Fr?i��ҿ��8�Ԓ���,f��2{H^���M���/ޙ�S��]����&�磍OAE�{ Ŵ�>uF�'��L�bb(5�7���&�=����	�J3�WU�*�g��R���lkh y���=~��g6��_r^�$����?^�W+��wg�&��~�#]c�4i����Ȅh����:c~�VE���U��M��!��x�û7��������K4%53�j`6$�"
���;��D�
���XڼĄ@����{ջ<��g�%�g���iOW���0<llc�L������3�c��3�ɉK�0}��	f�_��Jf� �0�#�j�QD�Y����Fa2]�/��a�Ez� SI�ZZ4j�;�8����'m?�b:T�m_x)�T�~1A_���x~i�	\1���/�?&�w`J�C���vCQ�	�Y�~U�<��K���B^��V��5�=<g�E��o^�ꡒB��v�Fd��Uj�*�붶CmH��L���T ���S&*f=�V�=K�q��)Y�	�o�=�&�r��˒�q,3��dLKK5�
�v�oa�d�+�'�70|��ѯQ"����׶�8���ADB�!��1LD�*J�ya�J�JJ� ����
�՚YA���|8���K�ïA6����z�I	Aq,"�,+@�J���D���#�})�5��*�e�fU�i>D��۱ �Q	��oFM��%1����[�Ȅ��k
$b��d�-bN����NC"X+��oʰ�� �j��1r^D�
���BJ��A���{�.���V���ǥ����B�"3T�P9Y�?��99p`���Ρ��������rlj�u�Oݽ.��]���O_�R���0aQ�Uu*Q
ۺ��^B��z}����/��ڹ `jk�
��C՜��j�fm���Z\ϓ&-I�����D�,�{4q��8�X�	sv��
�>���Q�����U�Y�kt\t��T����I%��t)3��H5��d�@��~.���tC��^i�=��_�ʕ_�	"'s�
-�3~�����!�+܌H�x#�u����h����׆ao`���<�F�o�E��*ͅs�&V�Zv��f2��@A�.6ǐ�_c���:�t�ӧ�8�f
,#�h�%���O�^[ $�����J����� 27A����K���V/���0ENՌ�i����CXA���P����!�����ŋC�}Y�q ���{��������6��mc�i�}� j+v�_ݬ\��v�/�ħ��#�R�i�^�Sz��|��6;"��
�N�a%��i4裩�<?��A�<��\=�Z�%!��7Sݕ�J���n���?��Fc��~%@w�]4:iW���i���Sk9 �]E�k�ɨzF�=���'1�1�^239��f!����ºW^e���ArLӧ|�'Z�m�B��cKG�l��%4I��i'�P�trSR��%
�B��JCuQ����xt�/�T##[�H+��}�=d������*dÊ�&\
|�io�c���l/W�F���h���r6i�&��}�S7ys1s�>ի��6�ṮzS�����ӝ��n�<ּԖ�)�Ĭ��:zlh���"->T�Nj�J7����h��o��P>A�R;�o�!���nh�J��j<Y���j�k��9wF����1k`��Լ�߇�ވ�7�ͻW4Ndy�h~�FϚ-	���Gɯ�2��k>���x��m.g���w&��_,�W�Y'�����'����� ���G��}/�0unˏ�nĢq]_�Q4>X7hl�{�z�۲���*��g��A^:K{�9�E��C�R��i"�\�d*���^/:�Z�lF[�g�Y��R�1s|RQ�*��ʠ����uNV��ح�� x����@���������AI��aZ�E��U��k�E�<�T��tÁED�o�D�m� ��"�����r}�/,��]�`�é:��3�a��L�]`����X��o ѤvSΗ���+��Y�yj�n1��� �
c,W�RԻ2��.<��"F��A��^W{$���@`�)�Z�Hgn�'���LBe�Ӯ�`�/��h��;x�Z�zެ��M�_p��)�.�L%�d�7��Z��U�����:a`�yV�ܥ��M�.�rZ�!��g�T��&�78�A`8��8����8Sgq-�)�I"\L�u��+��
��\V[_n���âL�jOai�ڸ���e����m�8ԅ���hZ;�Ͱ��'16ѩ�SP�Wh�#��_�dx�����Ub��yCs/£q9v(v��'P�&���4��U�{�;~�"$h
����^:�S:�����_���W?��|W���0��䌔����+��S��,�e��#��7k��Aw�uw���Y�Yɺ�.4`hT��{N��R�&?�F��`�椹��N���4?��=��S�	�wPK	��9���?�B�G&��^~�S�G�n<���PBA��?q�_n�`zőL���J�7�zrIr� �J��#�q�J�hH�R%��{3��V����"[�~���6�Z����gn%��t��ю֬>¾f6k�U� �+����x鰦�&��;�B�,�Q�r�|.ʰHglV�O{�$���AC�-t8��H9ks2����v5��r����1���'T'�4�����������T��Mlr�J�]F|��e��Lu���¨uะ��\���6�L&PMZ��z��MM/φ�U�A���^��*	+{!C���V�p}6�ߩ���#�}�y�s��(���*�t{{䂐��\BN!en��l	�����Nw����+Q ��=5c#q-;�0I��v�[�Z�p�e0y�R�+���Ǫ���7�)	ʨ��[��&yٳ����I=���Ҷ�JH|�?���7Ń#ő'm���۹����nNN��� �����=ċrrQ�{��]	�v h���,���V]�kh=�L�fN���D�t��z`C�