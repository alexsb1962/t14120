��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*�s��W����*��%3R8x�l�a[��_oS�3���
�hfAX�A��gF�k$N!�_>�Ł�����ߊ� 5"}
���I�L�VB�y�(�hf灭X�l���q��c1[i��Pa"LG0K?7�<���5��F��nuӰ"룏����
�M�{W'v�,b�C`+��+�
`�ȵQ&�3+D���@�	�m� ip��m�Ms}LYv{Ĳ�����$z��F�Y�|�93�B����b��z��<u�|&0_���}��x|�ߦU7ip`���i�)� �9r��NeX+2k���5�A��y�m��M�G�B�<JE�w֩�B�yYO�[=U�'���.��g�P�^��.�!�\9=���?{���DL׻�S$��	u�
J����"� ПC�FP/P~K���4M���t�2�g�O|D����dN�)�f�8o��T�Yh�l��mSu�&x�����;"�۬z�: )�
b!����6���Nn�;�üh��q;���2�$�&�{�]�7v�m^��k�I��ۛ�{�P��r�Lkk|n��H����=�j%8�v�Bd,�G���Y�ʻB1$L���ݠ47:j�I�c"��j3%���|�K�!At2�f���;ם�@Gy4|�U��mZ� B9&a��\4&�I�3)�.���*Kg����ڹ�h&�벍�48����oΉ?�1�ٟ5��#�h�%ʁ�R��h(��?��OC�q��C�x�;#�������&.p^�iv�1�vjY��������y�Y��@O#V�ν�2}�ZIV��;����Hal���ܽ4��P�n��E����c�:�ClP��f,gJ_\U+�bP�Y�%��Ҿ��؆I4e�ۉ@��L|���ĸo6ɓ �u��W|!6>ť��D�
�dIr��G� (�7L��Jv5+Ŋ3�:�#��)�L��� X�et�1��֌Y��)�t�G�qE��tړ_(�e��S$�ypXʧ���x���@*��G6;���B�f4P>E��C�wnv��s�|pv0m � �I��ׅ���xhd�u��xYE|{b7t��x3aƷxYf���l���g�"Ç�fr|QV�3k)1��Dj?'��i+�_�Äj��Ό��CX�#�0w0�+~��=�\=h����`���B���sMa�?���E��a&���҅#Uy��7g{)��w?����U�X�u�,vI�P湼����P�K�4r�N(�A�q�
��u�x�R&cK� �����bR��p��ndZ`�Ii�R(�d,��<�I�P�4!�2�J����TV��Dw��}�x�,D�yK#nY-����C�nx��4�Mo�N���rpsr婴2z��r�E��}D��c���e�WF4�p�Zk��un\�����F1�}�*��q���H�Q'N{���ȓA�M"�)�2O��[��f��Im�X��iS�wg��1&kA��/�X��J�"��qbؙ�����kyL��^�}i�����e����OU�zW��G;�zR�+�Z6�:j�[0d�-&��p�'.��$�~z����Kg�J�>����wD�LV�
�"Pi���W�2A;���R�D�M���n�]�����խq���2������vY����b�Z���(��7�N�My9%�5UK�s��̏������fŦ#��"E�,%�?�14�	<M�_"^h-�����8��c��?�788�3@�ӳe]��P�`X���xNE�Ui�;��۸��F7��
�j���De��r�}�Ҍ��!��[dk�m4���b ;��ȶ�vVM}�J#�#��\ЍF�ѷ���	A��b,(�fD�#c�X�zk�T���Ŕo}ݘ���GV �X�jQ/EdU������v� j��ZR�NH~άV�C���1���]��M,����4up�.�����b�7����+%e�<�<�\�a<e]&��n�_�r�N�K�A�3�أ��*�̙����ɀ�L�S9�l�����hh�.�(x��s��!�zj�AU����4PQq�������0�k(8]lmnTe�Dų�ZG�'kb�|�8�&���my�"�p��1�pZ�ϧ�3��<b<� �c����(o��|W�k���ۊ���e����"�3��W���+��Y'm͖��eV��l2#x!�C�>��:����̎�zu�wvنwCK㧾���iRɲ^T�XCT-(2�V�!��jf�$�A���3_��d�4�C��=��P��%������_�S�%�-P�L�&X-��q�� �OoOOj�H���i� �W���F@���gTi������߾�r�#ϕw��sX�x$��5�M�v̞W�!�:W���$���cy��R��j�v�N����#NZ�B�p��
��Y�
���H^��m���z\K�(�`�4n��D�	3n�1ÉaKEf_���42ȿ`�"	{�@�#+����Gl�U]D��ʱ�Xu��D��b�s�9))�桴����br� �2&<�	5CMA��?�=���y��A�fb�v�
�͇�1X���iBa�%	�AL�sw��k���˅�cgmfE��~�#a��q �el�FF��5�T��R&����gB���jI0_��ais�|�84|m��K���l���فo� />����K��O��0@�ϓ�43�A"C�`���:�6N��!�>�7߸2���$���`��t�3��.���?*J¸8��QsQ\97	���I|�ş�<�=����>�A�~k�8�t��~M)��ɈG�q�rx��|XW�b볰Ih���II�S=l�F��h��l;])� ��&�W�D˫(��e=儖_qY�as�W��k?R��R�]ˑ��L�2�j�>�y������G�I��,k�_���ąIq�{����Z2�(�@�w,P�({=�l_<���#���=���(v/7�h}�ۥ�!ȁ��T��8~󅼤�#�X����1��d/��i{hl�ޏ6`Wh�vqQ$�vVr�23�Ks�}��s(�q�2�ci�`����ؗQRfE&׺9,f�Y���֑ocz�/�,g��]�T��ь�]!W����C�8= ��=��b'I�9�ܛM�V��Z��9�\>4������;�J���3z�S�K�<��:���V�����]�V�����s�.в�.�)@_�M��Y-��c�ZY�=��#�Ӥ���,t�q A�t����_
I�t7&?CS�U�Z>��"��擋wR�E*?�:��)�p�{�2pNT����$���Z�8�+t���g_�y�����D>���{��u�|\�3u���B�}�cLj���H�n�?�����$̫dN���x��d���������i�͌z)w҆�'xZ�Emަo�i��V���=h��Ac�s��u?n�T�ln�j���B�l��3��`P�*�Ez�j�[��B��C��2P���a%mwG�Տ2&�i���қlKH7\&�k���:w��z�7�������P-��؉��ճ�ȱ���-RZ�q�>�E�Q֤5P*Gc���ɨ��J�p���[��e�\�Gu�: k�w	�����Rb��.Vm���FO�,��8K� ~&�ڌ� ���Ʃ�h�	R���,���"�g6 p��Ƅ������G���|���]+�����<ZԤ�d����w��k�����~����s'0?�Z!(y��{���+OD����ɕ�aD'�/�Qk7�14~R��(Y����I��1�@6�w��Fp+!�E2Z�q�ЖG���$?f4�LA��C��7�5�iX�,�|��8n�?����	vW�/JmZ����'br�����A�̕�c�\�� �f~����<��FL��������c5�S�F~�l�9
�2Qo�t�L:�ߪg/��|�
v;e5�R�1�\���]{(��|J�W-�:r���񩟹s�Xi2��_^�F>){M���K��Zr�T�E�N�+��ud�AF�*-b�oD�8�x��w�	�O)b��C��^��8뚆�CE�oV̢Τ��j�p7	m�E��K�.�?��K�)���D8+������I�!��PV#���o2g?�@��i V���W���[t2<@�z^n&����ɗH6˰�Jb=t��P�#��E�<�<�n�ِ����Gl����0�˹먴�{��2�l?��q�y_�����__
��M�ۮ��q/4L�'�\PuIܮ���+�ά��T-��h��D��+�U$~2EX�X��!��M�� *�a�W��Di�����d�:�$��14�a��״��Uc�e#�}SE}p+]ك�s��A�W�!:4r�>J>�� �9;5Y��/�c,�Jƴ=>����d`o,Gc疶Plg5�nj�8��)ۭ�S����q����ߏ'�HHh����Ɇ�^��X���������^��Pָx�d�*��T�� H�S���*�$
-�m<���S&�N8�Zmf���c�#���F<�����PU�fq9���P��6$���#Rc��1j�긟����䭔�*_D˂V4��3�0K�Θ����綠��ۄ����'����L�<���׭��d� b�5so5
\��:MG廀�4*��v^	�q��!��q�Q?�
�B�������p�/�ၲI]�d�y�)�:��F��Q�I���mq�[fX���=���?�޷J"���w��K�(Ú	o���nT�5*���z�2���G�bT��G�-"h��w`~LxK<H�x�-�ǟ�αC2;�P�W#��bm��'&5�J�L�z���؄|��]�:q����ղ\BcU��uk�Ke
��Ï�&��/D�|fy@O����F�C$��۳ݢ��q���B<R=�	%�I�¸��vU��N}dWF�и��a�"/YNeF�Ҡ�g��Z/%��u�_9������W�Iˢ�O��[}�-��<]�b'�Tq�苊Y��(��}�'��ѓOK"ۚ��
�����9.��]}�W�i$y����+&L�I�*|������b!�Q$,�����]�a�щ,�cO�>�ZP�o{�אHs)5��{�q�9��\��Rl��X��~�ְ����nD�~�� o��Ҙ%��$g	j����s��?����WP��zqPuy�l�4bs�|�' A��y���|��u&)��y��=�|�[��5��b;ĝd�kv!�0@6���~ae��x�JE8<w�e0x��ȏ*���׈�4��?IŪ��>��N��V�Bl��:G�
߀�i�KQw�3�+��;��})�~'�������n�,H���`��3�_�ll��� �1�6zgLs�~�b�z�(Y/���R��x����N��ʃ����u�Z��S�դuo�����,Xݣ�>�����,a�X�h���tu����h潊����V����	�U�ɓ��L�,?���+-~#y�X�B�z\����L��0�8�Aa��J;�}�QR�؈
�)C�#x��;���P[�;�i�a�G�p7�	o4���`r�£���Ő��;'t�/�i���Y�k{�n��{�@ sK��ڰh���a�1��H�yH�j�7n���kU������0��-�e��.��)�&��a-1È��>���Pl��"J��ϯ� �R�h�m\��B�uuM��0��o���Vu�`o	�-<ߚ\��b�B�6�m�<�+E/�$���vUXf;ɐ�|;�$E�ִ����w��1+�@:�h��E$�}��E�$!	�V:},|KM��z"|%��X�c�#_m�c��� �Kiþ���{V֩a�l�u��	I��ۛw�Ӵ��0[ƒ��3���M��%�B�4RA�D|[�|ftJ�	;�� �/���2Y�+��Xq�� �������Ӈz�R�����.^���Q'������H��FF U���N�Am�I��H���x_�"��Ѕz#���\Js��tI5��҇��
T"�$!y0±>Z0��[T�T�-KC��v�;v�4X�Y��Vhys��Xd[UFh�G�s��&R𒯝������Rw�６d �>0PlF��G�f>�6S���)��3P�1mw18����|u�[f�9���Y�Kd9��W�ѩ�gv���.�߯E��M����G��br�u@�ٶ�p���6ʭȄBR ��-H�����k��]v��].��x5��ܼ�����VزfۗW4.��p�<��L�ڥ���wה�)A]~PڭsӺ���"�笎v���,yJ������g�v�>��&��~�e��L�AL�Zovr48 U�M6�H��{��)��U3e����kg�k��c9���k�rݜ�y�]OXH�}�����9�H�Ï�
,�J�zJR��� 
̬��mR5P���'�r�tzW����x��Ό��gE�Z)t�?�֞�g�`\ B%�������x?�=r� $�Hz5���I&X�TD�{ge���h��C�j�����3����)f���0�Q^��Q�@1�f��X���\�p���<�d<���ب�8l=�5	�$�6����ZqW�Lc�����l����k7 �C�Gӈ��)��씂�g�"�A/�3���|=�5�;��͸[0t�9ܳu>zu�5�2S�I����"��
���d�6�~�vۚ	Q�H��h��<�;R=nC�%/����J��4)��A�ˏ��=�ȫ�m6^���(E�h*}285L>o(�O��<�Ƅ�;)R�g���ƶ��*�{�<\��_�����Y�q6�B�nJ��������-�	Y�z���2*���HQز��.i��또�d�D�c����qr�Q���2�ѩ�0��v͒�B�<䑞3�j�0/N���!���[+ihH.�(xs)������*k	��.x9��>5#���[�p�2"�΢X�?3,����@�����{�߰�s��Oa���)㒱������d
�7�q���_�[!;�Ni�YY'��A� 8i����˩#���~�Y�jؒf	������i�S`)I:����"HT�|���u�]��4�E|���Z���c��&y���0`t� ?(���4�A�~I_1�=T/�^���69~�}��U\	�2�s~ŀ�'�<���ởyf<W"��E�v����^�x��0߬: E�ւ���I�-�8��5Q�y��+2�Lr`�=���nuY�l>Е�!����(���[�uI�Y�4��#K]���'*��t���\�v@�� C`��:Z��'����}/.�;����"2�\2s�t�����n�/�����M�*�O��^�8�Լ�T�o���]��*[uBg:�e��F��-V��o/��ST%+���]�w�cMD0ݸX�}�dx�F��D�xq��5�p�t'��5=����Mi��s�X��yD�D�_h��8�A�#v48����Xa�h��''�N&�Cj��c����� [��b�?[���g�W�~H�B���ϐ��Rʝ����4됳�h|�,��|&?KZ������X��7�[�I��Dd�K�x~�(����SNv���S,�R^N�� /���{�@�.�H� $$6�a[O�=��P���u�4`�1E���%H�>���?*�Fׯ�+�~��驏�8�����u�m�Z���[���"�-?�g#���c��E"?�x0*����f:V����#R��]˧i�#
-����j�d�U�(E��D�8S����!z���Z�ևp�7f'����>)��E�n��2'���\ʡ��8�&�d_���-^������
8�=�U2	�J�`�m��c�Ϻ��0��hbp��}��|�h�����{�c�D���[���ǺR!�O�#V@v�k���4i�G�P�Xn��}�	�<\�)}����b�1�Z�[���T��C�������?��K�	�\��-���3�G�@ߙ��m�~�~_:Z�:=�:�-/s��7��9t|�!\]���y���lcn8��,�W&QŐq��ik����o��{d{t�%��A�L��aʛ��79p�������O�P��d������y�t&:-�KNjTc=JF,��Z`	�'��t��;"F�FO���06�G�v��A3�$h�,$�!�r�5hp�b
��qz�9�A\E!i�&E�,� ��S��t�g�6g�&�dݭn�7�_Md ��[������_�'���.��i�ZH"OLF6� �����X7��s%�͕�N 9ΠAO
�Wbf1����&��$��Te)SlgvH	a��Q	�����N����N�HW�d�{��S���q͗ʉ�U��I�������(��Yz3��le�)��`[ا�P����/=8/Y�Xw�I���g�流1=cI��.�̧
ά�it���5�3c�񁿄��#����
���U�Q��h#�x}:�bƓ����9f�~Yز$��
�Y�!X�8O�^R(�^�����岕B3L{SK��$Ts�Aɸ2�c���y�;�B��6\��Q�ó�� ��(|��T��׉��ܓ�Jr��d����ׯV�S��o�ۋh�i�u�}�/FM�J��c>�.0�� �o�3s��kg�l!ޮ�*�ty.�Կ��)W����&fB��s[�	~��T�tQQ�ZiN4��Xݸ�[�oEZB�m%��,��|Pk��:z᠊-�H�G���RǧϏކ�J3n�M��p��Y���$҂'�a4��x�گ�2��N��~Uj������<`��{܄����Q&�W
�-Ǿ� Ԫ�B.�Ҷ���~�_����X��4/��7���~B+6i|0b��{\�GR�a���m�{��lpGp>��6��
ijAJ/�����HA����H�w�cT�u�x�Y���9���'U�Nv�7�j�o����f#xS���kۚ�<�c��H����#��:(N��[
��}���v�1���´I�7b��=g6�ӫ/K�p�=�E�d�XƵ����?��>5�c�(��{��:�8-��n��-���?� ������L��{�?-��Q��p��Ve,.y�\����jΆ���!��(����(��5�����|(��1�+�N�澇CI!����r��3$n�<�%��yv��aM(�>�4�L`�p[',q㹭��0M��p��,���l�NS��'#����BZ6��aU���2<�G�D4��3���2�&@c�҄�$�ԋ����ui����-�)��� )��_�j4��d�R�
��zVa�%c�y�*P�&���a1^ +x}?�n2%M�����IqC�׻P��N�������@B���Sp�&?���Ml�P�N
FKn9�fq�0��"��2�=xNh�@G d�A�F�������P���F�G���PG�� ?�����Q�P]��)���(,��2���"	:t�l�*�@F�T� �I��'J���&�Ϲ�c���֢�j��a��42Ơ����>Y�)�LƯ��G7톗Np����(����HQ�N����4+Q�/G�jȇI}�+�+#�p}?f�%YU�=)(�e��y�Tο�[q~l|��]I��MW�{���j� v�B�@��:&a�(3P��uN~(5�����1ӝ�H>����!փ�PgKB�d�hE�8@��À��Q�K����-p�1:�4^e�%�U%0Y�OǈQ2g�Wz�{X�h"sH�~��� ��� �6�N��h�@��`�دc�h���Dc�(g'�i���h'h��s�;:�A���f\��oז��%�'��L;�w�6�*r��ՙ����7p���ѾwK_�*gc�aҰ�z�L7��,+1�
�{����w(C��+_�~Ւ�coL�w3�9n�<[� ��S#��aR�x�k[�z�B~�^�ԀART��A)6R&Z�Z�0K�t��紤š��MSiѸ�H4�W���ufd�E1��u}pmI�J��%�cyM��Y���!	��F�<�G(k���6�G}�>I �+���W�rZe[9�S��od�.f^�bȌ�r�"��!AD�u��6�L��Ɩַ3~��;�8�z��Uq^~���V������:D�� ���@��KCYw��&:�=�pN /�Z��vc3��ۓ-�:&n�:��)�_��p���Τ�U�T����?�ڙmp�I��i۴�,���^�'�l�y�0�7�����@h�l=Φ!���p5������L�	���;�G&o�t�������.�ˁ��7|��޳N��*f7����s�,���� �	��V�%X%�\�������74��O�=�'թ:��|�?���^�hu�2�����g�t����� �2�&�DJ�#9
�&Z�5�#��lvv~$(�E�I=���z9�Cg&w�`H/ �ʄg���<<,:�,��0P��Y$�u���a���k�M ��x��u�tr��'$XA����OA����+H�OTG�Z�և�3��FZZ?+5�����L4I��~��V�X �+��$|X���������T��L�KM�3b%��L8�;},�%!��'��5�mo�\���x]������Ix#��E�z�^Y��1��c�.A�ݟ5���$�]�;�n���%��0W�D+\��¾�׉ۊO@��:���^n�F<�4 ���*� ��`�'��b�v�H�_��;���T�n�h}�������n���:O�\��8�CmDfX$XΨ�����3�
�g(�٦��Ao��ִ���]�.I�*p݈�nl��-,CW0\��D��W.�ȹdȆF��[4���/$��M"L/�nݟ��>�i|
u[J� ]��z�}X�Fn�L�$ߖ��3��&�7|�ԡd��� �b�ۥ1���=&�
������Ë���F�*�Q�/v�{�*_�<�_�u���P��0�`������6l3�/��'O�N }8[K�@M��H�
~���$B�T��[��-�b�S2�>$��"z]��;�믂L�G�$��8�E9����5$��A<�
{"sp���U�b�[�����4��7��㿐�6�4~�u�qe�[tW0�j��S���dž��Ӫ�U���d��7��V�<Ųn�%�@3��ѽɜvؤ���9L�L�����F]����L�tni��tl�ɺu��F�1�lUp#@	�L:��4	��܀��b��d(1����Y���(�AŴ �<���$J^����ޯ���d$�Ҿ
��5��j��r��m���h����^X	{���܊{
����^�'�X��o����ƞ0���|�c�(���oY���wr�I!k�N�`�c}�i�W�:yۭ��a`N����^�iY��1��9Wˡ��+���Bw��+r;�zNQD)$�1����;8*��6u �脍;�Gz��}%��O���#7^Ԟ�����n��RC�t�v=�<�`"!sMK����k�7���~cGֳ�[fS��wj�	�o����G�q*�4�ğ�N*��{�ؘ3�����v�#t�#�W�ӆ�+�F���238E4-�㸢�s�2�s�C�%��̒z��]�6��-�e�7�1�M���i���w:�UUgl9e�9�:;�8y�F%3�����=V@�tu�����{��:Ǡ&f�d -�%�[���/Q��U��|1�w&i�6_�A�5�d�@Ƿ�Y#�G�:��� ��?"?�E�k=�c�CZޝ�u��S��:d�_O�ҍֈ���䌥�~I� "\6�y���'��m
�������d���<E�Ҫ╞bi��?�c8���ӛ�^�1O�hv��L���X�X1c�Q�3#�ۧ���#��:����p���J�`�K�d�t����{<�",ҩ̷X�Z��S�ٓQf-�Ǔ�i�AX��󫘤�"�~�Tawg��/W\"+	A���&L�+�y]��O����N��BN�?�I�jR�%�d#t@*�u-N���v]�}ғ=�ŒØy��.� �k��t�ٽ����EWFb;B��4�Γ�{k�#���`����=���q"C<��MJ��R-u�2vR��Z'5��?�
m-]<MlbF���/�����m�
��0�qԧ~%��x��K҈��:b\����f�x	V�XѼ��Z�0�Q�TE�R��b-.z��&��#����r�s��h���hW֡3�G��,8�!G��
M�wH����F��KsG�drK�����bŵ&�@Ԯ�瞼Y��W�	�]޶���sP6�\5�����^���i�md���>���>���v|�(o��R�T�q���Nِ)���e(J��v5��ј�}S����&I_��c��r�e���9DΏ O�5v�D���#5E���{�r�to����s�hϽe.�?s����1��O$D40c0+���ή!
��%Dp�U6��/�.�%�y��P?���0���'�j���b����Њ�ȿ��q��De0��}[p����˫j�����Hy�=+HQa�
��y�a��M�w����]��ĥN�9��ܹ�g�u6aT��-Ο����EW��yWk��O?�<vd^1U9��*��2=@��Ȧ� �����s�Wdd�>\���n� �8��Y�H~��z��˾IIQ�U�vG̭���p[b�h���w�5sƝ��Ff{�926��&f&��
jϖE0F0%�/�z�V�ZA8��b��z��@��d��K��:RG��5��>��i[���'��=���n���&�>��p�?�S�B�d�&�s�͐���Wk�Þ��C-�Xi��u
d�\_p-9ђo\뾘X�1���TB>���m�] ��h�a�g,��g͊Jf���e|�J����s�^�!�6J�$>kjeS�>��¿�9{'A��,ǡ�n؞�ah�y8w�t%���Z�9�hi�_�����B(�w^��JWM��6�c�N���iU�Xq��[���U��3!t�O�����@�~��&���`O�黲��mS�O����^��;l��c�f� j���!����B5������߰��9a*�x>0�̔^R5� 5ν&eGʉ�~��^��n9�X�<s���_�A�H�eS���B;HQP���x�z�%��%K�OӁ������`c}�?f�	�Y#%�.�ȏ�)	�i����%�?����S�K�f�N(]+	��9��g}N���ϮrU�X�;�h�c��[$���Y/V�fš�VݺN�&��݊K
���EJY� ��(~ys�-2���~sJ+�� FY�{�Pֵu��j�1�����R�>�L=�j��E�N2W��O�e��f�X����6&rD���qQ�:y��� �"���\�Ebt�We�Ljr�D����V~,�"������*N�͠�e{v	;:#/�"�`f`���D\*��{&lH�z��:S��@=d[��RG�4&��1̻�e�-a�D�y�!�tƃ7Q����[mB-3#e��L0(F�d�Cs���9�_�}&��^ܠ-V��2��8!X|`���:Ԅ
i�������Qk���p譿�p�>,3[��n!���A��ˤ��������m0lt.������������D�aK`ϑZ��8�L����MX�*��e
5vk��<z�-�Lo�s�=ȟune�f\6�8���V`p�"���X���ο�hk�L�?pa����n���q���@�N��Abh]�%�酕_aIh��W#�����������d�4�vB�b�]�N�QG�RZ����9^ð��
�gM݅{ˮ-`i*A9h_l�a��Q�4m؜�*�j�?��+mn��`!S�}&��<j������͕4^���}b��&�2ߐ�w1َj>�=En'PmЦ��8�@�����ޱ�՛�A��l���G'�?����В��2�r_�u����&��8�-M}���м�ס�;z<,\�9<�U*�A���gyYs�]�d(��� �T/X���
L4�Ok�dUR��!���{������y6_�syۺl�	����1@l����}���C���3��_ޱ���^���E9�湗F�+t"b0xv��'I�z�h��$7��,�ٷ���+�*���I#© ���B��FG�|����$�����LN(pjA2{�>e��������`����tȑ��|��:;�Y�,C*0��=6�}+��p�Bm����Gh��^6�xY�=�涴�"����C���_��M�t`�N]�8�|�Y&}��|uc�Q0=!��Qb;ⲝ�J�K|�"!�h���U%� 6Y1.��
��ڳ���l��	��v�K�|`1e��_g��=��41�I�j�RE�&|V�K�1�P]0�����:=!����:�9@���Lo'd�!Ah���֞lR n�*K:5��
�X�£��A�U��ڋE�Nj�
�Ԭ��Ԉ�
*>�i��u��ݶ��Z�)���gU��Ҧ�UtU.��쐎�Z1G"_�'%�C�B��:CF׊$��-�����c�M�*�YjA�����uE��p�Nxk�A@_x�V��uh�u,��dq�#���d���4}��i2�~�t����<e�$/�(��Pl"f�4�D|I*��0xB�;��Qye(5B�	,�=f�1�v]d��:q� �oWH�@ֵwG^��,�����,B�{-��hV�<x�t���(��e�lce90h	����.X�\���((�-80R�z�~���$e� .��	��f!��H̯��F�g�A�i�9���f�t��aX�RW[�\�D��$��p5L�(���c�jx�FH�/_�F�,;��N�<�˟~{w|���Yߝi�.�;��eC��nP#����_��O Hn8��z��ȱ����Q.�}�%?+�i"֨����;���6�1QB�ŏ�a�%�4�#��T�*��,W��l��_�b�>�w/[F|���4RS���,��=^����m���_ރ
vA �l�z~u�j�)�ܿ�W_�!�r�"
�M�]u�3A�d�4����'�0�j�i�:���{0I�Û�4��U�L�n�p�tpo��X=7&�>
��yd�mÎ#a �/��B&"�J_���X�Mr��B��l�$7!��P�B�q 90�Dd� L���3Ȍ��xjA�`xz-�I�O��w�Kg��E3��o
��Օ~�TW�K>�gI�T�-�Z��}ϱ�oc�����6��M�W
�.��0�@��z-&���N˕a�!�O>� ��'�0�A�3���D���Z�C7���Oj�=���xq4半��;t��]�%���+63� ��P�`�g+�=O_`�ԟ��X��L�.,r/�e�+h�6ꉁ�C3���4�:�+e�Oova�Ql�ǩ�$>e4
�ӏ�SW�بm�O�៍��	W7��/ؼGI>#�XXhh�1�e�X�lo�:2�i|�z�ŝΉȩL�
�/a�����[����PG3P$�fU�j.iT���>�k�D�J0�(�?����3#�+V  g���"&v�� �N��]$�mS��}�OB5��
"m��u)j��=�㫘nL�3Qؤ�̈́PC�(���m3��}��,#�;l@���f��1�C?Fȝ���E̴��j��և!�V�k�p�Ãn���y��aǥ��Ԡx�b���ʦ�w$>l���B' �:�C9EV��t���X��,�O�(��=�2X��{��'���f�GdIvG��9ƕ�wJ��w�RS�udE��`ٙb&`7R��L���ʵ���"S��Z|�����%!]�W��P�pf.31O������P��ԍm��$b�/X��*��H9�X�x=����	u��0�^8�Q�P���+��T����+��[�7}�h߅���	|��ɝţ�e��C'��Y��nU�����ٹ�-/��-#%G#�����J��;�_�����8<d BT��Q���o8�J􂒩�BZ=��CY���ϻZ���8�\��U>��]���/��#�C��ң�0����$��%g��N���D3�Ȳ[*#���I��L����o/�4����'�ô�dv&���)LE�	s�=���w�'������-��3,}��z��^���k6�g�;���W��6O����v-?]�����{n��ƿ��#qb�֐�E����ǩ��u
_p^�+ ��AE.�zt�66n�d�eT��������.�	x�S�~��b�W@Q,����t'�K_*,iY��Ih����-�� �N��*��_�$��4�R��=9"�"-Ǎǻ��"�L�9��^��^0���Ȍ�'e�ˆi.c�"�b^��X�ڡ��ʙ-�`�L�n,�u#��Zd�HK� �&VoPA��ނ��ڣף �_�H@<�w8�HN`<I��巳۶/1(�G��6̞�\0֚3�ʥ��0Ҁ�N��;u�N��j	�7F;Ua4#*
uy�G�G{��Y��]C��-�y��ܩ�uI�+�öe��7��e���4�!s��9�xX�����jL>� [�g�����9�܇]Ø�����3W��WL�@�e�S���1��a�	��f����ÔVg�E����"�O������4�K/<�7N'f=<�:DY��S>F�%�C�ۻP^�����
o
�h�5+Jh�Kx�
���=��<]���fu{�K�.l�b7�}��6�%ˑp�Xg)�54ǒk�l#�6�4ޕ-z�`AV��*�r�=���d����Y-P�DO]��w.��0�i�J��{���x
�E�uX�������c�Nj�,2.��Q�L��q�NeF�`58�\f_� ��Z ����s$���y��	���2�A�) d�o��D�6:R�a���FKQ������B������,�;�h
Nb��\�K7������J �D��8-����հ+��;ĸ����4�}7(_�~e�1�bOsᤖ�Or	��B���pB��E��*�.�YtX.�)/�F���{��r8{�/��݉���*yX��oJ��-+�����j�3w�bG�v� �*sh��E�"��"'H�ǟ��蚞e_����g$.��p�4�|n�kB9�vZ�ԩlj���<�н�
��"l|�ұf#Ǹ�.��aɝܻE!a1�� �?��P@؆Ӟ& �kB�����\h8ʍ#�]E^+���f,�QD:�3HqEWD�pu�<���
H��_�f0�,�J����BJ���1-K�c}#z�ku�P&��(��Fvx%���<���^�� R;��,�U:�"�"ڈq��m� �J���F�{Vh�����(�og8����#�U*l����3�<�dP���̽�����Y��/�=���.i�.uO�TK9��'����Gyh�3�u.]�:���S�eo+~BH1j����fĮDc&hx��F���
�f�v�^�/�H�	0��q]H�_`U�69���4�,�6)R�a=�\�*3�I�[2�р�5�Ц��s�p�Z��_�7��o�n?�~�Ft�;[��n:�"���+�/�T�_��U4A+pX�!�Dp����bzw���^�T��/�������Ɩ�����"T��7ۦ��s/Mq�#t���g= ��:) ��9��wg\�0ڱ��:���ܸ	7\���YB��M�``��d�4��k�E2 [W�( ]jR�wR��@|�n��uq��p��&J�צ�,n�����﷘�����C�Ƹ(�e����/[$_����K��GUy�X���T|Qp�;��)�r�4�����^���R��&��sT��K�jY�A6����S�h���'��7Xe�f�*r$C����{~K��aۄ^u�b��;����\�H�x���l3���}%���*�ů��F�Lީ6u�;���]������z�3euh�$k�O��sFɔ�~�V�����ٶ��b�r���	��{���Gູ��t@��DC%iՉcu��i71nz���b��\�sB���KF��~X߉c�~�Ј�"��d(s>mM>�8~�v�{�"�����'Xr�u�X�E�,���!������7s����kf~}�!�C��	��$ ܔ�J���P)��/�M�<��E���F�;��z�+�ZI9>3La�� �;���^�D|�ki]Cb%�X��^rY�߭H�a��3���8��`�:C�,�_�5ϰB���R� �e�M���l¾#Z�K?]7;�2����vfry�l�SFD$�|��B��Hm_N����Y0�*�@	�Ĳ�N}u&ũ̖�E��C��{�A�n;>$�va���-�!){����K6�'��1�u=��2扒<X��-�t+<U�0�P�]А�i�RGuFߛ�ԔS���_פW����f)kK�b�>I����}�N��րLݹ��zH�GF_}����R]��kճt����`����-���%@��>�b�g�皒���[��9W�@��-�	s��6B����swAd��y0�՚���B�|ۄU�D��D��"{.[����<�$0'�*�wɚ�Tj/&(�j(�hI4.�?�U�ލa@R�Z�^i`�\�}�:M�?�:H^Lڟ�"D)��W���on@+������n��]��b��vD�;��u���YL�XZ|D�6���l�Sַv�j��kD�'�r��a{���w�h9�,���01��B�����ξ�T�eZK�0�L�'��V�R��P��%�>��~�����}����Z�g�G]j��2�-x�h���5q�Ų݈Ѳ�"�[�+A�̛ˣKo���O�B=����7t`7�{�<3һ���Esk+ƫ%O�z�h5B���ҏU.����* V���~r�5!y�&��DT!�-N�F+�R�kb;�W�������<ݷ��##
�o���8�i-�L�����>$dD�����J�Kq i�l�É2~��1'��������|�uL<�������b�TJu+�#BʳB�_�
]�-��ܛ7���qZ-�K���bk���PC�H��=
R޻��$�u�	OT61�镓ͼ'�����U�?L�F�Յ�s��IN:��	���ifz����ODv'�9Nh�g9G�*�ۮ�f�
�O﹢H4T���w9��d��-�%5�
��J� �h�%��C�?�j���$I�����r(w�<���$AR��D��;�m
�[ȡHY;�M�;��Z�yD"�,C�<����~)���ݬ�]�a�U��i]���;Fl���O�Q��laʩJ���g)�+:��fX�̤P��?O�ɷ��S%jYA�q�ɚ��K�y�u"o�CT���xx��-�T�C&�` ���p�##� +%Q�>����qʣy���T�pX���tm˧��~�!�x0d��W���ϣ�5�y'��� {�m�e�󶇾�$J����8Ё��ߍ��iy�*�}I�]	�Jcǵ��{y�:���x?w	�D����y��h�r�w��j�\�9��}�B�����ة��Ik�I�G&�
� �v2��]$��`jf��90�NĬ�nZ�Gd�M������P~���f^�s:pE����8]zt鞫D�#�)<1#�\�<T�����^�>T-�� u�P�q�+�I����@�v� E�Xk�1��m�X�HFlHODu4x�A���T4�Λƣ���f�1YS�-�y�r,�D9ǕQ$��2]a)����s2PGH��\G���^~��:�z����7��B�����&��8�4���;���r8�w���Qo;d�+"n���)4���f2K��8��ԙ�F[dH�Kq�YU�����c���T��'%��J2����g��2��F����[!���r�wK?��4���2U��'�%Q�&u�w���	rq(������t Pc1��V7j��Ox�L�����?�oX��h�br�cv���v~�m�z�?#� dG'i�;;��Co�q4��%�)>kx/&�g荑�r��s����rr�5쇤�C��}��}�'*m1����ίж��/�����y(��;[)�9� �ЂŔ7� �U-�!?�6�����2�O֟�d�x��
�(7'�.5TУ�l2��~/��ZEU�b��&͡���S��X>�](��UGR}R�e� ��@��'#��A'
���*��R�$��]?�`h9q"~�\L-�e�A���_Bk������۾J�xs�}H�[�k��Nt�V�Q��w�Z�7$�v��>'�7�q�'%A�>����$����"3��ʙP�����dsР��@����\�oV�P;UuXa��#d�G�T����יG�`(D�H[�<5Vˢ����I���v�ąk�3����ж/�_��u]>[ ��ʒ��V:+XkAB��Ql��\�Ѥy�=ݘ������Ia=�����* �d���8��'Š�M��T�R��_�]X������K�b�N�j	h��T<�d���� ��K��g�������W��������nYk$,�]Q��H+S�]�N"SM(��JYu��6v$R6��H�}�h�e㉳r
�Z���;�s.��15�*킜Ph��)�S�hu. �B���i�Ն4q�ڡ����Y�ú%�Ȫs��Cn͂�s�M�>%��<|{����j=2yH�Dx�a��E�����Z��>f�J��nѬ�B� ��I�'b�_�V�ܛ�gf�k��`�o�����qТ�"�z����)E�/[U!t��*J���
���-�q�m�Q�+�s�:<�P�0�qw=Tkߢ���GV"%{a�%��$�@ІQx�0N*�F5��oy;e�4�QH&��#c,�������F�;��6�T�y��}�o E�?n�t�9�p�Z���m�������\U��i�7?�\�eͽE�t�[���,זg�4�%���ߐT�S.�����.�q��z���&5�˴���Tݾ6ov6�.)���⎠	C�A��t��e@��٣�C���Z��jc��ռY���z��51��JsT�si^�3��z=+�{�/�ø�-ͯ� ��pְY0c"+{,�0�5"vD�=��j0���@���Ԓ�R
E�St����A������z�F*���W0������V0&�aRlhC�"����>��;f��r���D� �(�m/�=,�pmgt����e,���G�[5�>Po�m��$�o�"&���,���|U����R٫Qx����q�N�Gb?��V�QS��G��V`ړݝ�L��c?�6p��e'?Y!'/��R7k�S��֌46?�ݥ-7��J�v����K&�҆��_L�l���D��b�e��̭[�Q�G�
!��K��<Vab��2���`q}���5����?�Ջ���X$d�>cl9�~�}�� �bB�V���Ϛ�� c �z�?����"4�HU�6;��U�-��}(�zE���+��sٍ�m�����H)>.�|H1c)���(�Z_r/����X=����_�0.p�HS	0��ci�F�Б��$�M��c>WT���)�m��a���V=����%C��`�>��Åg�[����.�S2k*�p|�s�W�:��.��=�/�*y֧�9�s�a�cF�Dr�)�ppx�|�D�?��1�+K!����#�%�8:n�:Q�A7�_�)�T�hg�)8 5�xsx<p�\����1���sK�H�(��]����^�`�T%���%1/<�ژw�:�Q���
*���A[��՝��_�ԕZq�':�E3�@�H�Ɋ�=��{G~o�@21�Ь�F�kl���|�*J�w���=����6����+�*e�G�$:��m��@X@l����i�؄��n֖-������[�G�*�߀L���<V:��_>������{�8���ٵur�k;���2�ב�l�a<�n�5��i�����y��vvڒ�+Y�N���L�^g}��&�!ʇ��+�F�t0�� �V �Kt���c8���MI��=�������Kv�<�#�O�8-'�0�]�"l7{m���s���\�{ƌUԤT�FrѮ۸~�k�y��h����EQ)�BZ�
��μv�͑�mj�HX��mV�@̿�"����`�WQ�V��hygHD)�q�ΎA��R@İ������2�ܺ&e�r~$�v�4`�z9����� B�!>�P�ϡ� 9�3�ٔ�(^��E�����c���a���*����w���u��J>\	���K��4��[��__���9_�FEu`e�2�@3P��\̿���>��+����"��I�U��{��
���L2buM��
]V�T*��