��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�Eݹ+@%$ѝbNs>�%���%c�M��e���Չ8Q�;��0A)֟ &ȩ�I��=�N�q??G�s��ˬ�}[���Qα���1�-G:!6U��c܁e�O�#���P~H���n�G�O�C���3��>��:��Gҁ�>"@�9��x�[�����u��}���i�d�A=dx��>�q�At<�l�y����Z&�����/Gb"��?(�մ�/TM>B�C�Њmz5��̎�#|������,�������0�x�$!�N *lj�U��ۍ70�XT�ep��5Gb ��e?�l�o�lZۂ���^OJs�ڴ4EάPWA$�
U�O��孡��O�%��+nȰ��Ⱦ���Y�g�c52o+���`�M��_��&�=?9g�3fܽ��b��ŤG�iMV&E�"=[��}jvɖa%?��ԝ�SJ�7��X:~��e�$k��^��- S����J'@�^��ܧKQ
�y?�ȼh���y��KT�}��q���t���`�ԁ١x���Q}�����6���T�fH�ى�ʡ�m&3) �J ��?�f@�#��5���T|����O1�FQZ=�^��鋯:Y��_�Q[]��ߛHn�����w����Zl#��	,vѮx����a3<P�}!�:��б���Z��P�����J�Щ9��ѲsY�*/d!��$K����ۂ�Ͷ ukR"��ޖd��]�Y��רe�t����:W^�Q5'��`0w��q�q)J,ݡ�Ia���ӥ���/��
(�w`&[����W6	:,�LC�y��p|�?�LEf���Չe�	:+��4�{��ԥy�*��8�z���ll���p�R�^����U;ȹe�E^�Q?�qw}-J��#$���v
���E"�9��H���~p
"�~.�fi\���=���WB�+��8�i4DgE�EA�j��m���IZ��X�~��<�Jn�@��	� ��-�AT܊�W#%6��G�F揈w'A�GT�T���"sr�H����8�"�x.�E��z��>=U�NZ��I��G�U%y����Drs,<f:�˽g;���)�'VT����,
��	���]��2����N�ॱ��n�Ix���N��NO��G���4��8�I_Ax�ῡ�ۺ+�K,ߓxN�3��Qr����*	;.&_�ؕ�M(bZ(*Ya�E�b���R�I�2�4m�a>xy$�@7!�d���ϯ���G-���4��$��!���(���n�6=�����Wc�L�OM܎&E��q�l��5r
�y�LVpg$[õb���*����U���4|�O���j].F�"{��Q�`���ʓ��9t1
�쭥�u`��e�9����x#h�Q%v���8���̀��E+ʽ�`�,�!��|�8g�y[�
�m�X�ha=�.��'!OMc����5�;����gFu�
'T�m��J��,��2�+=k���c'g� 
߷xWd ��k7ŋ��K����"�u0[j]�.���yУ-���,&t6R��툣2�%Mc��ł\K@���(��^/<�:;L*w���%�,h�L���T+�\J�Y7L��#k�!��%+/Mx�ڹP~�m�@�Sϴ�§��Ϧ�q��}��o����ZwTL���q�,(�<H=%8%f��`�'S,�V�л��Ul�Ԯ)P���od
퇿��(���K� �~yx�,R2���v�+�����\�4�/��*�"����_��A�%5�E�ʍ�$d	�֔Z3p���Y��l�Mv3/'����ܖ��uĒF�Ӿ�'��6��B40�ݱ`�R�Ź�a��wF�"GLߵ�0�D?j�[
!���1:6����2'���t�'��m�(��ܧ�%f�9�����z�$�7�)�v13�.�@j��~��8��F̔�ڒ؉��V6��8�W������MOi�)w�e*�*S���ղ�6WRӺ�˗xz���q�<�����3E=?͖�0�x�I�56H��
<M�-�q�6�b��O��7�V�Ó<���r��f��x�]����[9��jb
�'r��@C��p�A��訰��������JW�"	��?2���=eX��Ѩf�Tw���'�D lg���́��%ü}���c��&oL�;XЂ���u!�ߓ�FI�~ j"� ��g���&�2+��<�[�!�N�l���ߣ!6���sgL�#���C!l;�ԡ�K,<��;��9#�1f���`���{��z~�.��L��e�"��c`��bp~h��#��Ŵ�}�{3V=礼F��P��㈽M!�aaL�yJ?Y[�i�i��L�es�������&M�p3�׭��a"�k�_�M��պ�:���Z��y�#�ev���c�L�r��Eɳ@?�ׇz���2��9|L"�5c� w�i����6�?F?����WK����䶇�ϸ|'t���KSq�}�9^Z94k�A�����Ù|�����V|P[� � ĕ�s&;�� īd������?�e��5���8�>vS�����ܩP�[�έ�x�G��|�y�׮ǵӣ9�/�w9~���/�E'�\_�Y �����C������I�����j8 �6v�a�L4k�1�FTy�[Lt�n�rp�.�S����p�Z�E��/i��"Sm��B�p�ϰW��JJ�l~݆+�N�1�>�}j������iT~�Ԍ�5�N��>�D}Y�i�^�I-$r����9�FG�X.f�K�Zp���:�Cj���)�\J������G�K��b��ew{=���Qڿ�7��7T�X���=��|xh@7uMuZD-�� ����P#4�x��	%W�|�G��Z�=i N7����qsh�u�
�>�ʿG��b�*�ķеp���ƈ���l;S��[�����҅��P�©�R�f�J����;%����D���L�,���	�N�M�Hv�$��-��[t:,��q�hM%O�&��e98E�ͫ�*�["W��������3�l�҉XQ�B7˄0�-J��ҝ��&&I��#��Ofg~�\���.Z( {b����y����9qw**�A���E�'����������x[3��tr"A�e�,?�2������d�pg�NjZ���'Y�:ҿ1�/�6��|���K&:��I�{���T���9�\���9��n_�-�l��`��id@��t��G��WO(�W�Ώ#;)���[���
��+G%:$sf:͘\��d���ȣ��0�1����� Le�J����鄎>���;���ю�q;�]�O����T�{�N��Bq��p��������$�V,[����jL�E�.�!%��f�ψ(��dG���t�g\��*�mG���;�wub����Ul/hX�֕7	4+f�|l��aa��a�f2���۞(ΙP��g'SŘ�p���cM(�� 1��M4`�ә�݉�J7,�)+����vJi�g.������x(��԰�p���K�� .4����/H1�M�� �����.)1�s�)>�80�4�-�i��:ۚi����r�m���tx�$���X� @���e���pu<��f@�t�ϻz����q"g���\Ӛi�n�^���1҅�F�g���*�i��ح�"�S��+�H�d)�iFZ�s��Ų��~-���c�r����!�Ip��\Q޸�J��B�Z5�`���SOpD�ž����3��g��V�nR9����� Q�Ӫz�LJ�k�p���.�R8)���O<�%|���@��Q�U�ж�$w罺��g����" ��P��Q8��������KH9!dw�`շ�{
�� ��$��wz�M6��?pb���
�j�xO�;�~�ݍ���x^��C����li�CM\�ӿ9H�̓-!:	�wT*�3oYil��_�gƾQ��,�z֞�,ɰ�Q�=������Hq]�:���u:�d�o���0蕙��o�9y��l*��e-u�Xw�5����8���Ҡ�H��D��hv��p�7ȌB��{�즖R*�rZ���_�6�x>�d�|�E�~�brr����"*N�ݗr+|&�Y&���}�,��V~`hɬ
S������=v)=<q���}gɶ���9���8IXn"�M�@�@5t�]�'>&p�����ڰH.��'z�����^�A�$ CFm1]ܨIE��	垦'��h�4q���ٔ^��%��|S&f@G?k�z91�9�#C��
��X����< #Rz��]��zλ`���^8ܦ��e�#�����[�[��᣽e	�h`K�*^�-�4h�����1$���	�O�2��h����@,;j!�%M����)x.�!@��#<����t,�T���"C*ZG�_�_Bd�^�=Px6��J�[�0�y�f�%���`?�����d�d�x�����F0B�QὡT&�S�I��� &2d��#{ٕ�r�P�tfqB)j	�"�&U��y��p����J��9p�e����da;��J5�]`k�� ���g�sGAfznI̓c��.�Q�\���q�k�}�����YOl���E�0z���Q7��F���-�r7���T.~Z����drI�\y2Dρ��Bݨ���$|@S�w*c�+պ�2�Eh
U�rY�Hc��|�@��=t���j��d���K�x��14F1)ZF\�YV�Dw�@�3h�F.�ҹå���!U��x�p�X��(μq�b�����#�<� .�k��*�3Ѽ�.V�BK���K���ݟ�r���eWL~���o<6�`쯨�m�X�1�H6��%�b3~U����Nf�!H.Q[��D�cm��z�F�Ko	��j.�q��B�_+�]D�ս��i=K����/Y��y+d20㆝�|���5) ~�A"���N�_�Kˤɯ6���L*�Fl��5���|��gL�3V��ۓ-XK�����'�c�|�Hx(�Y� ����>_��z������L@����"ǩ%Bml�&�շږ}K��2sYH�#��Z�r��H�"�J7����Y�֜N p1 �����CDc'��-��@�w��=�& x��r��H�?�3�T2���]��?���҂�k,6�n�s�l��y��Y	)a׿L�ܐ ���c���4����z��EzY��SR���7[_$?�c+��'IU��c\�i�"�'<��=Xl~��h�/,�t@/h�R���8Y�0��J���k��6�j��(Uܧ�����m��1`�C4P���H�ɔ։ls���j�޼(y����-������r��������%��x��?ਟ�Fp���/Z�A1�u`@8Fre�C�It���f �G����Ef�	PSJ�ѻZ��������
'�z�K��8�>f���n?�N�;B�p�.��:�i@�+t�p��0B��ϵ�t���5ŵa�d��'��)y쇷$y}!柙?O��|�z���d�x���\sO�&��K�,����еߵ��Ÿ!�'|A�wt4A7�����
�R��C�&W��i�,FJ�_�o<_�Q���R^>:�L�.度f�K��4��7_Q�O�'��H�	y≠�q�4-���K�M[n��6|�����B�#�:��� ��o����1��!=��TXi�A� ����4�̎��di�]���^�/���b���ȱ��C��7���������t� z{J�+��g(,pߺ� �u������a�Ϥ�㤄J7�"���n������i�b���#8��׾$B��H����3����z#��Pv�^�����6�kzB~5��#�nl��6Ы�G�XRx�u:��c"pJxڱ��"�w%���AsX,T4���M��l#���I�c��8�1����g���]���k4F(��>nZ|�ΖI��YŻ�A���=��_	@ap��<Va�j��^���e��d��� k�1U�KL�z*?��q��YQW�y���?�r("s��.9Q�X�x��}ˈF7q���g����:�#J�5,:�^ߪ2�;�`�0�� N� �c,^���)�Jc��i� �'R+�'���Eh��I3oZ�ŉY�b
j��2���E�f��h	���]ֶ�>UJ�dl�F�4�:.���Ð]N�Z������&X$�5�7�H�S�"�0Et�9�c����x������;�gh����	*f^@��j�]j+�FCn�#Uvl�uq�|��
����KH��'����Q)�Uuj���-~�L��Ԗ��M������?�I�A��ǌ���InOs�& 9�a����k��<����yL+;��Ic�!����2��
���䱉n _F�ݘ�՝F��wS�"�6%g��ݱ<��@�B-�y�?F�Գ/t����q,;���Hۺ�=����ڧK:l�W��\�h��W�x+��n�͆��q ��3����ԉ��
�G�u�݅.�&t��L2o�T_y5Mnx�0]=o��1�;l:��S݌!�:��{��7��9��i7�g�0:�-*�?؊���pkRkl5����;��ybm��q��.Q�dnj���i*�$��E��(]�V��S�>l��d&D�y�hnK���0gi�;�[i���k&J���Wd����u�Y*+`�;td����mH�{o�ҐN�ۦ'��)��o
n�|�.�=;q,��51��ʔU&� ܭ@��ɵ9��/��>�5v���(�I��CH�_��S� �5e�'�x)0u���ER`G��=
�I��]A�~`���H�,ܨ�DL͸��1cNrTC��x�sԉ�	�FKVdk�&�n"+L8�V�qq���T�΄�@
Y�&����E[Rg6�(O�1����ٚɀ����n����\�ӽ����0�0̌>Gn��*uP�j��s��\��D@���F�p��oj���<�u;{���g��H]q(�������#� �G��^bhc�@�Θ{m-�2�Q"k�t����˶T�p*�\���!H��[��9���<{���?�cyHɲ�p4V�5���D��}�2����\h
np������Z?4p#N��U`�&�����ƚ���th�"'ԓ��U,^��ca4DL �i��GXR%q�{n�f��s�K�ڧ��aD��[��N"`VL�o����<:H��*��5=$�ve��׭
^F� Q%4�>d��q�ES2�a#vs��oBE2��x|�� @�]lF���y]�\"�X���v��R~=��w2J�գl�Ų���%�����-m��Ұ�&���85�ذ��ӟ�ƨP�a3��9����#�n��X��1���/��ߐ+$��U5����%�%��Av�v�l� ��`�Z����V�X	F�l��1!�eX�H^뷙ϭ(᯼�~�"f��c����|�pc��rs�&/� 6BM�s%=�(�����=��`�iu�PS�cM�6�l��x(�d@�<R� ��-8=>co��.���Ȋ%Jb��^��6K�ؕ6��'�e�:���Yҟk������,�`Qk9���QU�{�bV�yW�5�ѹT��Y��Ok�;Df��2"�F���N�^}v?�هG���ٹԿ_�� ��్:&��ћ=����\u���{D���>��jv%��b) lJ~~�w��!j=�9��,Unoڭ�Y]%�p-�F��J�~�)��&`�mU�D�ju����Z![���H���j��:�u։-W4i�V�Aє��y�h�L���x�\-x0Psf�,��Jє�4�餉�R� l!��k������������tL�B 4��Y>�!��+�����PgJىՋ��MX�xT"���+R-CѴ�+?���h��;��a�|gK�3L�;��/!һSᆎ׼�%�$����X=
�<�C�MMD5@�?iHh%��v{R�h����mPv1K`Uꕤ*��g{d������O3��
B�tkHDy[��)����(��E�r�%6vy1�#��3|�k������°߽�ŀ���C���~a�X�����V
|�+�����tx��Tz��X�52я5m��7[��1W��W8h�T���8m�qEGU�hw�u?�cϣ$fF�Nf�a��������U�b�(�Y���vO!`<�!���4�����i犁�Ϸ��Cw��r&�p�µ�lQD�5NAB.��?��#(�Z�Z$e$BÝl�b�<HV�|і1��уp/G�AO)�ɜ� .�'��i?~L���P��js����b�������^����#(�8��^�GP�b�;B�k(?J��s�:X���܅!��t����?/0hL.�8g~�pA ��iR§����Oz}Nd�� ��@���@�;�X����D�5���n󱉢�	��R_
�<8��/-��]���Y�� �°��
��K���#���^��a(���?܌�W*���Gl�8m��Ɔ=�[��Z��e�X�ot�<w(��lltM*ZI֦�94=2N�X�M!#ގ��_�K
�z��~s�uB"]v`V��S�Rf1~�\}�x_}	�ہN#=i�}人�2�3�U���5%k\�����8Yd?,a?�Et��@�r5����C!�F�諿	 c~a8a�p��>�z݉�4���ΚG?u>�H��6�C�˩Ͽ�����)�� �RLL�QA �7���
È�UUk����&�=�Y���*�4�m����	�m������b�]��'��!�j�W�)�V.'l3�s49�t� il�4�J'��<��߶<�JNXYg��mU�63qN��C��͹B��Y�,U��Y�>ڰ-���o�@e���ϡv,��%XK���$�����yNO���.�D?8��R	f�IdG����ހ��JU65��E7O�L f�'�_����p �e�si�?ԌL�_�����x׮~�cP��Qu�֪�^���A?�H?Pj�Úނ�B�v՞�X�酋
���O:j ֓��B�w�����@T���1 8j�R[e��$<R5�L|Ზ8kr[!D�p$�y1�Z���$���&P��/�]Î�t&��(���;ڙb��6_��@-���s�X���Pݡ��<c��G�'jG*��mt!��˞��>i�nxR��!��WM�w1��X��)�;��)q���pC����a�+�]�)�ew�M� w��	11柎E�S�S�� P\ƭ�s�WԻ
��E+/;>n�1��CiAhT�~��D[_G�2��:.Y��L�R��ݧ̞u����<U�A+kvC���@]�����Хw�χ�`lW����TD�[P�:��<�}��Q_�*��_���e��]�r����a�����]�a��x��v'�<��HMe��bM�/v�̋�oS�;�E��U�`Z/}YoQ�W鐒Wlu�D�1Ԡֈ[���2�N25��wq<����vEl���sj���tL�9�0*1��d��?Z��4VЧ��j]cCUI���ȵ_��:�����z�x���D���G��!� ��L7>#R�*���H�*� �`�"��� �[�y���'H�������{s.�'L���F����x�,3�
?}Z�}�gIq�*C�Ǵ���!�����$�]��d��i�\�b�L�?C�rȿ�ӯ��N�s`��:��]?IP�౱��Y+�k�{⩴,�Cd���Lb1w+��]��
��ل�f	��P�UMS���F�k���$����d��K;J��R��p5�t��W���`Sƾ�����@�u ���A�j��m6
��r	��z| G}���Z韻�5�ɦ���`�~�Xh ��U�xF��dQ���H�u�22^	sW����r7͒[�S��&�>g��+�<��i8J-������q�#��"�9q�;�������|��o�s;{Id��x��)b�5p�@��gZ'��!��ۜpy#�#��<�0_,�yTϮ��+��O��@dY�U�tGȟH*�Aq�=���X5��K+5Wxvc�[�8l�ꮾ��ѹ�a��h#[����Ӣ�2Jb̒]�f.��r���u1����ӈ
E;�$�/�N~�#1�'�޷�c�!D�mJ�aj4�ą�:a��Λũ��D5h��3����닫M=����3[�5�?����i%�m���r�d�;��%M�
����������/�dR�"Kf<6JѠ�aj
������8߃k��	��D�(��� ���p'.Ō�n�x�?$ܕ��,բ�&L�DL���y�
�%(��m6�t���p-�t��&qPv;�B�=���+��<��
�0ѫ,Tп�;W<���e'�J����&϶�=a�����ƀm;O���C���}��|达���h>ݕ��P�
��f�s��P:��L���a�8Ǹ�֛�ݙ��!��/�� �lb�ˡ���+�Q6�����{y��&:�X��SJ��kZL�aĦ�@a�ʬ�*��X�$mf�ώ��8�Dd��.����q$��֎�����КY��c���{2Vt�e��9m�P����o�x�_��<e̓q�3���c�������} ��r�4��e��A�����`�O`��t�1p@��^j?y�D�w�ù����(Q��lJ,���y���En3$fL�`ބ���h��@��A��2;(%n}B�(�>�T�b��Q��<=�JN�ozJ'�C���P����)�,�&:@hݏ Y�PQϤr~r4�V]�Ϙ�T?:D��:!�7��+�\�_�A0ȥ�g�# ���HEߣᩍTe	�q1��ó$7��²�ʺ����������f�ƶ����__�	ӏ�AR�4�(�[}����lm�
V��p�i��l
$3��x�k��ls*����P2xY-\�ƙ���z�u�%�ƨa�_c<y�a�O^z���v�3.6\v@Ľ�6!	ḋ��Iݼ��؎o�xrp�0�'��MR1��_����jc�)螶��$�z��n��"���+�o��z�
�U7p�i�6~�T�v曤ܟ�v��\�h �	��#I�K��d���2Kj���ܧ_v�EU<D�-�U.^[����xv`�6��"�j���B��D�m�Տ�t��j�]>���e���q��ׅ��Ң��F�4���]���GwQH*0�'���:
�y��-7�'.������n��:N0�Nᖬ�.i�>�m%�� ���M}�����P}0 n��u�F�;1R�/��-#�+���¯ڐeP�u��:.v������HO������g"��WN�q/�3I�]P�V//�_�	l8nbO�q1��\��l��N�E�ldA�c9��P��T��{@��m�o�B�8�.<=k�&J�g!Ck�w�gV@�����u?TGy<IGt>S;��q�|��W�S@�����E��G�SНи�������h�6��r>��3~��k�;2�*Q��~^��h"q����]��ti��tl]�?��,L;���ƮzA�n��둳E�fFCm�bт����3�ͯ�9-���3��ۊ�]��Y�d�4P	��U�%���-�0�5z�6j����P�-�>����HH;\�}�VbZ! �ԆL��ee�ǐ����r�!��L_�#l���z�Τ�@���"��������oJ���s��TB�5���IPR�{�}��h���;�L�Aj;.l�{��z�M�Hm�VNd˞w�s�6<J#8�0�:2o��+��	�[��9N���C5�C�@�L���.�1��N�����������^a���Dr/�dL�a�{g
��ۊ���g\@F��$��>Z���+�r�̛�%��7��n�!B%^�P��ڣ� Dk&o�M`�Jt���)�)\��m`��Ghf�<������R��	d�]-I�a�����6'h&U�����I�&
9�}�;�TļRr)/jܽCA�&R��
����4�	@�����*�L�y��?#Ϻ���9��ɓG�]u ����[FB�ӡ1b�l��|�A������N $=/,#o��J��7U}Iӽ���(�M�e~��K>f,�h>*����\
!��#�"�t�Qgl�&I�U���]��(���r�����h�@�4��.oz��|�d9S���'��C�S�9DW���NM��V7���]`�B�z0	�6�S5a3J`x<cif����o��ַ�v?�ȉԏ���hLIr-k�\�b�!ҭ�^u�.���Pݮ-`t �Ѫ���)n��W M|��W�i��&$��"��3nAF�D6s�P�a=�O<iИ�o<�7��!C��[�������g����D��G��y,JS��ICv=���H!�(�K
�4�zU�@Z� :�u�%�~;�\l��7�ͪ~β/wU�>"dd�H��i�2�Ry��A�ӬG�Pw|
�����)/o}x��]z�Nw��u�ɼ�f��	�N�&�m�:�8@¹������ҭ�Ϋ7�=Ѱˡ��u��ep�@�1�R�,��&R�iʡ@M��&:���F=���W�a�Z(��-�G$�FB}t��u�.o&d�/C �j�əD�Ξ���������Ws��R���J�=0Q��99��l�7�/��w�m�c�¡�iR����'n�4���H���O�����11]�{�FT��d0b��Mu~�k�I�I<��|���5<�7|��Ev�����O���n�䍖j~|��A9�?�K�.u����h��A:d)���g�Z�(|7bI%�%���`]\�d^���Uf�; � T�BH��j�2f��'�̥��`�r29e�����G5�@����;-0~熅�i	+�m��V��ƗJ��bZhT�Dy�5��
 ���QML)����,y��ofd��1��iy׷JNk�j���zٴ3��h�4�_ݾ��I"���S�����/B[��*��{ZN-䗡^p���}��9Q^M�:���
��]�l�hsKL��(ɂ��� ���0�"�=��Qa���N���~I�>�KJ<d�*(���n���"9vu?,V��`$ޖ?�g�&��>������&vX�}QOh"�֪}�����gR�#<[��$F{���A>�`�y���ZUޝ���׬�_�?��M��Mms�����y�$YI�����ٛVey�+~���e�Xx�����/�C�g�r��֑�WT�d��nP��(�>��ѷ��h��Xk	���Џ�Q#��~�N[���Z1>z��R�B��տ8��h` ᱈B��{R�0��	5���rt��|��K�e>�$Z��3"��j��(V�W����
����E�1��C��足_.-P��j�Tp�ܲ�|�5���I1��"{w���l�!	�XI���M*�,��u3
qc�S	����F���G1�辐���� jTE9X+E��*�(�A6X���َ�n����M�>���[r�� i�`!O����o�_���iHdn'�U����C�Nu;%*|���m֮4��6?���>(��O�L�L��p��T��*��,sy(.im���ܨ�kٕ�����R�&�4v���s��v�T�H�ôޖr���r]$���f�:���^6�8��#tC�ao��hI���hoɀ&����ʉ2my�A��@�Ss�Y)����0-�]/d�zv��	��R�'0Pp��Y��F��V7���/.�t����iq���K����H@�qI를:p���og��X�8+��3`����\q���Pa�7~Hڑ�n{Õ]�M��{���"/fh��L̺��<�����%���Z����E=�-0Q|�|��۽*-�xц_.�������;`�HV�.m�1[�҉��t�N)��� �0�Dzvt�Z��^[LvH�����7J��bi@��"9�S�����Xd��n@����Aٓ� ��MqF>O�(<֔�U��7����{���
����,9��G[YMf���͕Y������GW��k����N*;�١M~ ���s`&� �Q�>_��B��~��U|�7��1�U��p�EPj�X:h�4EOC�+���8��-a�?|�4�NUS%����uO(�?ޞq��qސ��1���o�Ͻ��hJC�K����.س�W���-�~ްi��u_�r�:�CTP��P �NP:�<�9�p�S��lY�`�@i?��H�ė<ϫ+p�b��.�{U������{Bd�T�-����w�1|qe���� �ݭ53�M��Z������"�y��h���-�����1�m6ٻ)���$To�VO�=���wՕ�-=��*��6��̖h��%��gh8iJ���L�,bߖ��4g`��P�]�t"�?�X�;15 �2�Թ�c�S��0+0Q��'�33��S(���o)ԩ+�6##CV��
��~mO�����#`�д���<��h\f����������ø�j66	�8e��n��~��k%�����A.æ۵#������Y��v���?>����g�2S�)�jV�y�G�$��8U� ���Y�'��E'����U_!<"�SH�5}Ihg�%9|f��?QP������Zz7,NV�?���p���:�[׿s��Ю	�th�Tx�wOS;e�����=�D��"�A�~�V����W��H�p����?����n��OI�!Q���<�jv[��P2-Y��^�8_q�k���#�5�� F����6y���.&�H���$����#'��z��'֏0ZJ�)�R���7��Aߤ����3	~��Z(F)�F$ǧ;���D�:�_G(	��)�9���`�fy���Ż9��i���?O��B��oXŇ��Q	�7<@�+�
�F�@Ylϥ�$���2�غ�UO�4`*���<f�<������j�g s�+�l��z�6Ud8�M�oݚ��*D�WǸp�k��h���\U+�T�#Nh��un[�(X�q$�M��-b�:�ϒYFܞ�j����'�VQ��f��6ꉶ)8�k�Y�q7p���5罭���O��4��s:�����5���2���H�����7�Lq�c��z���/�=�<[���}߁{cM���%Y�S�MR~�w��g9�NO!;%��$6hE b����
�VJ�|(�כ��+��g��5,X�7j敽Z�6�9��y���C�KS�}���������l���z����I�.ǚI~t�H}��"1�P�x�TҠ�-��ow��fL�ՒxP�L���:��˜���ci�s�k��<k��D���Z�D@?v�:�P���k���Z)�a�.˰B�v���'E:�qŋ'�J�z�����A*x�����9��h	tŹ~�o:ĺ0_%4�#�0��Ό�Ĵ�t"J+y���:�(R���c2���3�/�ņ���i��.yK�i�Ü �5�/�R��ª�����to���>���J����mK����fяs\����929�<�[��.��nK,k��G��9�D�F��V�CR����7���Q�9�� 6��nɍr��_X�S��Э��c�!��/hw3?w�zǉף�5_�>����,�T=�N�����v�f�v�-9d헝Cִ�+��qI��bB�����THd��%y�ƛ������go#����~3�8��k#P4Fp�u#,XȠb���}���P�T��ySd�y�o���bA|Sa�س� {3AX�ePX�+�i(|�ƱR�ic$��44����� e��|n6Z��=��-��9"��X���/x����.$2��}�  #�-��]�wa#��'�4{L�>�zK�}a��Ux��>߿Z:��!:��t�f�&{
���@	w�~%xD��b��u��u㨢�!��1�&�IEO��;UQ� Hs���tEY(sa�1�[���%1ǘ����;���~�p�xc�-�<���[v[Y���&/-���3@��E�����]��4�ԯf���`���_������)����#� ��蝽(����K�}%�����x���u=��U����0�����w-f�a�.fߠ�\(���s&2�ݐ�N�7MI�cH��Y������sg<F��!֥�qT�́�Ƶ��$AbҞ�� �Pa�e��B���t��w ]�'�s(�ltܔ��N�M`����A����>��܉��,	�{�M�O�y�"�j�#B8Kj_��P�5�}f	SL�1�ˏ� ��w�Y`������:F�6j�*�ނ��^��)s~�h���5�,�:��v<�e�����b;?f �����z	n=Y��М��Y�2Q�n{X���ւ����8W[����rچ�ǹmyۨ��CW�p�&�ow�[F�{ߍ�6�L�<o�k��=؀���]rJZ_�E*b���nNՊ�_R{ApVѕ�����\MD�̩2����$���!�v����*�ű��	g�:4QP�-{�Yd'P,�vZ�?e��>ou�VlQh���L:b�	i������N+g�C��iU:�����z
y��h��f���G��jv��q��\7���7�
���ġ����Q�`D?M�Lg���cm/��U7����J�!��Rl.��%�'���Ր'8�&���}w$6�@6��
#��k������Q-�K�F����]�k��ʹ��h�
]&$�OB�+XJ�̾O����<c���O�A܈�Ki���G�c���ω�����{%&-YV�/Sc��i���𐸨dp��_OmQJ54T�B�f�������V�>>r�ݭR�x�'S}���{?TG���Ff"x��f�褃��ʏo�'�Ǒ %�@�P�[��~�'!���Ҙ������IE�J�=�A����`�\aw�����@��o��n=i�l�Gb
y�x�%|�HYJg��c��Jg�NNbxr�7��j�_�\%�y*erp1.+(��ϒ0"�'�Zԓ�0���h\i���gm��7u��i�l�ݽ�$�?|
�)��(O��}�#�IdF=2әm>	��s��{�ΐ�:v���]m7����N�!q�rA�09��1_|���p�A���wF�.{#����фc[���(��#�RF��2��8$O×�ʔF�g���1��6G��>n�B�.�ף�i���FV�j�T��ƩمR�z2�T�G����(?��g/�Z!�xw��v���3dg�tb�,<G�k�w�״��޶��ʎ��G��������.�<�񥗔T���>�M�5�:"o��k�Q;������Y�G�J�(�ϒ د���R��=�V7mD���%� m���G�N�q/+;��[�a�1r�����e}�n-a3˔Պ�qzR���З�UNd�>����tj�5��I������-�;�ﵧo��ù���D�v��~�M�Nvn�dN��F��o:d�ti��R��r�����Y���/���������~a�}]�b�`���` ����[3z^h�g�d �P�٠I���k���WN�""G�E��]p߶ ޘ��U"�gy�e�|m�2S{��Of�Yb����;t���v�\:��"��Z&�I�t��<[*�C��S��\�go�:uѧID�d_D.lF�w��C̤�M~s�� eb.�희1��g; ���J�J�s�h#���(��&mYH4���0�F���zi���`/���ʌ�.�p�4�y��!��"���h
�N=��W�2?2Q��ˊS4z�
zbqD���q���g�[1C��u��rcCL���#R;i�!��&�d��>Tn��W�=�US.H}X�G�k]3���5½����*(�'b1nR�C��-M����UQ�̜�}:�}������W�H_�� �(޵:	���bBt��n@j0su���J�֋�%�M5��h���ׁ�:Y�w,��A��	Ȉ4����=�[�0�<>!��:���P@��K�=���c~6��쾼���?F��8��5K(ߠl<��U
������ꉽ]r��w��5<�#��Nwg?��_��Ӆ[��^�c�R���/�Tq2��.�z:�^���*���� a��K]d\���l�B�p��ȡk����7;����N�Ǩ3&�-L0���ڢ�S�Ng5b�Y�V z�!��#TX���8\A�e���|n0�Z�hקJA%�ց��.O�T�[M_o���4�J�83l*����F���H	2?���~_@=V,�Y��9(ZT:'DÑᤡ=��'�
mѪ(!nMe���Mx�X��*ple[��O}zPR�j�X42D7s�,@�ݙ��Q����5{͛ԑ%��
��#7���fuyo����sմ�g}����R��A�J�2��������<��	v���Ĉ�Ā3�^���U�5��AE�u�D��� �r�sq�@�X���6���o���F����j��3���{d�j�Ib�{�����`���7>��WV����~e�̖�R�ڽDS��N�ٽ8թ�3���tR�	�F[���&4�����l�S�N�B��� �g�<�K^��aXܠ�ejX��R����Ғ�;(�&���)E:e�ώ��`�7���z��q��y���xP��{�y���53VgN�	����b�g�DVJXV���$�D��77��\s 9���y��E"D��X�_�
����^R��ȯ��챢���ׄL$�J�O;TIpIp��:�p��y�AB���ajN��;�9�f���N�}�.��ꉇ�U��O�8���X�0����tJ7Xp��ͣ[�bER
�Gb$��B�m(��K�8Q�#Qz��Xcߓ�,Dh��,:���.�(E"��5�H*E�ŰK��������ĂU��A�Y)�܋���a4��vpd��"GPٜ�Ǐ��L��I������3`p���ҷc���UD��L�����n١KB��ow`����X�5ݹ|���eS�'�9�����nd��w{`�lТ���J�)�;�����H�\�Ut_���H�Q�:�^�g�u��G��=�g���'A�%D�EN&)����@>�`l�tIn�ßQ���Y4���QF���d���pP��)���7�2����N��灦�.7bz��l��˱��Ƃ�� �-U�j��؏��C�8�0H�ٯ�ƭ�{[��_Z͡[�*��un�=�9u1�OA���	�7�D2|j�����k�s��^��� !�Pӏ�G�\�J�N�SL\
gWiut��/G7�2�����(C��0D~�tޡ�(Y?���!8
�l���|dI�޺���]nw�$�'�J���	�Dh�@��EX�LT��.6_pPݮp���e��=�h����{��Af$@@y���/^�����Ƚ/�_����U.}��S���M�C���^i�pa�aۏ꧷��^�r�{YRW,�� <]k7��X���
�|w����yɷ�;�O+п%�F�. ӳp�$��>� ?��L�Vu��?T��܅�p8�1�|�w7\,���4.���W��.�0$�ꛗ%��$��%��"?%��.��n��I�h&������/��xJ����;�`�Ȇ���]�
㠥Ȝ�o���o��+�uǵ�k	�̛���Q��ؕ�y�����_�K�o�T=���hų�F�r��lf�[��v�H���,$�փ��KN�U���7v���gLB����4����>v2 s{�wg�w�y]����;VB(��6�"8�]���3�pu�z��*`��RM��ϿÄ�:��l�.�@�M>��,b��`_��e���-�����mˬ�Z�*��Q�ԇ����Vߠg`�2B�c�C?��67����A8yX%�_b&�cX�� ��p��o��j�����a�ۖ2����r�I;�䌗���JV����hGGP�8�*ݿv����9����OہG
���ӓ���#���,T�����P�Zr"��,}����^�*��폚��ǓhK;�s���v��?�uAVyY�I��{VqG�I�#�SN9f[��<>��OZ\p��K������-x��P澬���jΝ�jO��.r�D�]�^���_�5�1e� ��h�`g~��3"���Xk��&&��a=��Go'������L��%nv�m1"D����G��ޛ�="�(8T��^O+�B,X�g�s=|��.���e�������+�#��o����.��F������NG�V�&��e�rY�>`L��p�Z�#qL������[�����+�6������х�U�H�n�	��ؗ ���t�
&i?
�\���U�� ��[W�X��bc��}!a��/T��~�R��r���XDI�X=樤Jns�K$za��EjT.���#��0B)��i�1�CK,���I�7�N`_e�@B?bݴ����B�IsQ���Q?jB׆)����o��G�'&��_Ѱ�* [!Z�ֽ��-9�W��<�j���I�}8u�[w�o� W�&�P�q[1 i�e䉠[���%/_��Z��s�A�Y25^�*�~�w̸9�Y����[*�u6��"�i����$2��$�x��z��w����|�׍E�v\�E)��Ϙb���R[Q!������L�r+V��o���Y)+�]����\9�'�p9���8w�(�`��$�#����%��~Ś�<Z�����81S'鐡)�X�y!׳
U��(�6�n�Φ�b �.r��'���s
w�Q@0�б�O<}ʩ .�0��EI4���Ccy��s,�`!�h�SGq6%w�H�-�:	��*�'_��'e�?�[�}�}M�ئW�d�*�kꡙ���lp���
K&AH�xC���|���n:�G����7�FA�7"o��q�U���	�!㫵d���Ά��[�=K�� +�dc�۴���V	���Tո��2�4�3��W�z��8ET��Oi#$���G�������nT��(>H��ڐF�8�Tn��C�V���o.Ԃ��~U�jk��:� ّ��B5��-�lPp� �0��b<���X)����&HZ��w���Fɀӂ�CT���
��X9�yc� ��L�ʎ� t�����a��Se�ӹ�	2w��y�ә��������/�"�G-��TQ�o�Nﶅ���bH}f|��tz>�W�B�i�$���A��=�����%ꎶ���u����˅f�y%�w�������Y�V����eтB� ?-����,`�{�������,xP%:���>�wN��GҲ��%��E���z��.�e��/'B�e?� �cQ�|�d<3D��#+�˸�K,�)}X�H����`&��]�4) $����d�+Aޣ[C;��|W�IX�r-��S�BO0����p���
"��9aoC/4o`�ۡ�3K�R�O�Rpr�Ӧk���r�}i�����X�#z7yZeBṷ��Y.v�o��0��8(z5|��;�.8�Ux-m�k@B��8��r��(~fݨzh;|^՛_DB�Y�wԲ9今����|��G����Gj�>�?7;mN��M�W�.0��4+ȪƏ%���ԙC5���ٱV�D,a��i��Þ���ͶY�Q�d��©�/�f�s�qz��@Lg�?B���>W� T=T�U����:�:�'rI��9�m�i����X��`�=�O �������6���\z�u�:d�������4(I�|�[¿��!q�������&��p� ��}�����Lk��l�6Wi'-Gz�p�~Qo�CZ&�\&��*��;���\�%8�D!
��Z8s�ݶc��rͺc/���V�Q½	��EŻ��U���(MҸ���'a~��V��aD#o^sQʢ����V��h�@4l,܅e�.���0��A�P���2N$e�A`�y�m�0u�m��Q�L���f���ly�g0�pHSX��}�zK� Уw��9�N�U��ʀN ;q~��%ל���O y3N���sS��?��f�v�g�Z�G@:x��N-�[��%��|�$4���םl�6��
�&2��!I<&��,��>1����R��
Ȩ��!<[�>_�/�$k	�=��l� cHUG����iV�;n,�p�$�����Dd*��)@6�:�I�B��i)���,�rۢR~���������$��̳����8	�{Q�T�IO��M�edѷ!�%��(�r�)��@|��;1��4v�㐐��\��p����c��'�Ʃ5�b͔��q����p��:�N10�+di���5G}5@�]�Wlo�������k�۫�����C�+gM�%�#Y�'4B�Ǜ-��2����z�����~�~y��s���x&���]�rE��c�x?x	�Z��x�z��P�C�&1<�k��v�	�p�esƆ��pw;�7��iV`�����y��������#��d�J1J��ġ
�\��G>�Q�NX�1���D�������^��Y,^�1��$4#��t���d0j�"A��?�'3]H�wU�)b��º$8�OfD�����l6ߦl�@좓�#�@13��T{�vY���{jg��-�p����ha�+��V��W"��� 2�`m��̜�gooP���GYiD{�<��T6�S2stьd~�j#������|.���!
����E�[�f ���>�"�@�4��f/��Q^�������[�򉊾�T��:D�($���˾>] +�)B>C���_X�Z#�5���i���,��
��ś��c���)�M�T�DP��Ч15Ǡ��u�^�E��3�|cL�RA�\q6�,��G�eo~u�PQ�/W-eִ�-ŌC�j�|o��8s"�{��
S|X�(\�_)S�|oA �h�VA�����rm�&��.�z��X�&V��U�!Ci�����$'H��D����ο9���W�F#FZ��mAu��Q�F�[��
�����ͼ���9[�s�R�އ����!�:^Scw�����O2����	0ڦ���$�<�� u�S:q.j�`���������D�)C��I@ی��� ���ь�Ӭ8!u���������gMz	�[H�x!�z2Ǯ�M]��.I�D��Y�P��`��D�D?>�K_[&%dv�+&7U�� C�!j�`�@���ѯ[��,)6�w��7!����r�/����j�@`շ��^?���i�q|��ޮ%yc����u �5�&ʧ�oG����2��-��׮�I�,8��\T@f�2u�"� EnJ;S�:�/�N*K��]Biid����9�1�D,�j%�p��Oo��w�:E�#,���_�q\x0F��݇���&����[]��(�ˈk���T��K�Ј"�GN��ń�wN�,dBd\���A)g���d{ـ%����5)hAC�Q�_(`�xX!`��z���Ss���n�{ߒR�B�l��G��{��g�z	�09�v#f��$\6T���ٷ�l�
����\�*-�eҖT[\"  �'j�,G*���g,Bcj%y���-W?�܂,Z���y��,�KWw+��)�v6i����f��ne��/���ST�L�xz'�U�W�'Yc�b��c��r4I#_#Ǩ�|M_�* 	S��Ҋ4��ս-!�ɇ��hx�2���b�}�\��)��nd��)�ܐ���O|��E���"��6M�D/. �Dz�٣�j)��s�j�s����b���sM ���cv0Lg{��~Ƣ.�0�=~Of�/H���2M��ds�er�+E�I9�(˲�^�8)��K�$�KUB����[�C�;aoT5B�A�Ҿ�!\��nH��n�URKa�#�����_�M���]� �`��H�^G{�h���J]��K<^�}n�L�	�CD�x�iU�(nX	��,s]8����D ��`Y����u���?����Dm 0"6��8b�}y@�m?,v�*�9:{;��叶�Y6ob������ل�a�3�����p���$�l`��ی�Hc��_S����,W�0�O��b'�k�S�
qs<eo!��1$���	�uX��3@�6�'N8/��$=y��	�*45�N�����v�1C�Ա
DA4��`Q�t��Rr��{K"U�~f	J��s�_*x�����SH���|K�pcm�PZʾ��������f�H��F�qsw����q�MPy�(�j=��#ݚ� �J�הj�i�T��'Yɱ,q=�ʊ<�u��y�a@�"������k�㟄z� �j����>���t9B�hFf�TT�sJ���S��ÐP0c��p�3�x׍b�J\�8�'�Bل����0�!�-�bL��J�P�Uϫ��s����9�w�C�,���l���Hv/AIf���� �lR����R��a�$��*a�<���|c}[���Oz�5뼌�%�ާ�.Qyj�y�]��O̽�����[7� K�/�ić;i�����l"V�^�S�������f����E�|lƴ��(>.8���́w��Ck6�@Z\9�6��u@�}+��,�>��0�;�i��w3�}�d2��t�������7�b)Q�č��V�}�k��x� :`2X ��x9�0���i�!����>7L�����uY2A��d�i�;j���Q��֞v��Cⶨ��ȏ�<�ءPL��9����m'�Ѩ���v����Ԉ �Q�rTR�W���R�(j��a���U�G-&<o�_ � ����
�~4� �����SxՍ�~�ڒ�L� "��խ�n",�7s�u;,sp����踗�����OƢ�/���oi����1��v���	��4^��e��Wo�?U���^&���Hn����`0'�!M�ۅQ��A���!Bi/@G+r�kGdܒ Sǩy��I�\*%ߧ6��I����qVg~t���*>yO�@g�-��>�ī�WN�5�\����_��='0.�������>�)�l"3����Nj�@�ʂ_P��U��j�����*O_D��cs��3��5�T�m&`��	����N�{ʎv�Umµ���1��*�h
&���T���;��)��V^��"����i��3г�w'��[�#�,yA�,���2.7=�#���)�ų/D�:u]����p>�����˜�|��=q�r�Z<����^�?fqY
��:tg��Zu��1e�ܮU�4�F�D!�0�T�5��_ �$HiT7���٬,:��_R;*C��#������۶�J���	�Z�A(9@;V�����<؍��d��5��KZRD�
�&+����Dj���!<��� o<Y����zI���j5�<=$.^�����h4Wph�Z}f w�K�O5T��´k��TFf�y�����"�������i�ѷ;����`�F����Ǧ�*X�����F�%��毶��d�3���X�HI�
��qs���Ye��e�'�뙸��D�u���_.֩�t��h_o�d�]K|Q�q~O��j�эj�~�����\�9�f�	�+(M�V�	�[>��=�=�MNAM����3{��i�W.d|�G"D��*8��-k��K;VSY!�ֈc���7�#���fJ?�8���x�*φV?&�Q��V]��,٩9��ny�� Cu�,��<<A՞�v���!-���׹�XB?Z�
;�2m�xH3��lAw૾���=B�dF������f�ބ�Z�1��u�Z��1e?c2_�h�^��R��F��_��2n-��*�"�+V}g��G���L-��&�vP06k�|R�f"��V�4_�a��u�,��KDx6}����kl��R	1DY���~ل$���(<����󊨠���
��E�C�J/,�f4y����������d,1kĴa�����>b�����քJ�l->���٢�[G��d$;��r6���3�-I�쁊$,p�d1��.��u �u�k>�f�,�pS�6N�ZlG��!�#�	MX'�~�K�����,l���3���r?�#�����"�,�"����t��<fs�H�ꉤ�R��2�R��YPI��W�{R�L��|�ʎw�����Y �-e��j��1��j�qX*�>D�P��X!�^��ΰ�^��I|d�Zg�z�s��ÅԿ�An�i?'�4Jt�q4��cĊ
O .�P�a(���"v|�k���1��w� �]�������r͞��B����@�CW����3�B�>�#�����j�8'�����S%�m^��+��X���%o���Wn�*�!@�LWPLв����"��"�'�&�4���ͪh�Y���|˱d/�
�&j?i��C`3�R �G>Md�j7 ��Lr�g�æX1q�$�K��[qC@`��G����(g�EJ�)u;;dQ�ZP�H��ȭZ�0N���c,�m���Ŷ�.P(!�vQ��]|ߎ��4�51r��sz@�"�aW�k�o��]��ȳ��9���sd��v4����tv$7]���X��Җrx��P��������V�9A~��p�-�W�(H3P��ciB�]���r@��K��>pI��
f�����4��-V�o�h�,�<�f*��*�[^���)I+�]m#OsDw�?��C��������u��#V>9���]!�;��)"���>Ve���.���� =V�,��H�����,�m��8g ��i�&��~�֠;�, �� ������q���!�A`Q�/�'${�)y.�/0)З���:��N K�7�
��X��{	CxHCe�7Ǩ.o�"�c� �*�*��W�]J#�Ղ����)�jز��&�'�`=��~����7.M"8e3��>kmw��m&x��#-�w����8͈�t��Q�|,�)���5�T��u�sCH�g{Z3�6��z���"�;��`$�atwlV���Z��=6&F4{�ei��b�����eb#r���KuO�����Y����n6%�>^M�PT������Ա��CB�O�mr�\��CU|(2��R)�Z>Eɡ����Y
O�SQ?o�B��9��o��4��+AʲW`P�������9�_��:Sg�U[JF�.��@M k�5��ϼ!�V�:Q��(���k:�Tyc�w]�y2*jo��J��ȿZ�#��R��j�RK���L9�f��wK��VJJQ2W�fk@t
���H���-�u�(p��MUEPâ��*�Cz����KF� N3o�ij(�۽��K3a+A.�7�5����47;�w�@8��:���Fn��saM˥/���P?���l�A�Ҷ�M"T�:�5�}�U��J�1 ���`hݯv�|�%�n��_a�F3R7�� I<�[��k^���1�����]6Ӧ@Y�Wv���+͢�A��'ezf*r�9�.r�����)Ѡ�2t�Y,,ef�7����YRH��1��x�Љ�E,�j�e��b��h���g�몎�(l�)ƞlM�o�̈["��} =���ID|���p&rjW`ɥ�M��%��Ǡ�4�"�����b�f\�{����yƸ�$I��!�"����!�����O��G�rP�A;%��r�1�}�7��Ҡ��z���=Vg��V�k�cį�W8/�/6'P5S�W��W�Chh��0��'�\)��F��A�c�6��&�ad�D˅�̹-�v��[A�p�A��őrN�M�gU@%1�;@;�,iץ=�ȋ��!n|�_y��;��C�J|���"�}V(�QIƧ;G�n�[jT4�`s�*mnB)#a�8��b��у�@����{hD���7��'�� m�E���fzy�V��G���Ώ�!E�m��>���|`��L 5��e
�L����G���C�!D�:��ur�p�F��.�ڌ�ؑ��-#���R�x���s7D�����WP��I�2���Z�)�.����xX��5�[�L��)���#��R�?�nA��mY,�(Y ?�B��މiE�i}��M��ӳ���`�|���I�:�Sr:f�bJH���C�8����קB���<i��4{7ϙ�����
�Eӏ�Xx����M/� ~%��I�Ml%L	ƣj�WMSG|���L�s��M`r��԰دn����W�G�ԧ�YC�<(�U�y?,�uL���#ژ��AE�K�|���Fו
��o0�!G`��B�>��1�Y��q_��F}-��$s��ȹ��O"�1������q�3*��\�V:e&eh?���R�]�mD�:ʀ�^B�:n��,�n�x��hV�ЅϮ_T�n�=��!�4($��0�=���w�ɉ"������f�~�鸲��ꯟ�T�J� 3g�4�F�'k���6� V��t�P� H&L�FYpJ��刉�������:�e�_�{yCq"4]d��@&Ҩ+*h�/Z��%
�V��W�U<u�w�omv��Xf��y��TLH�����۞�#��b"Ū$f����7x�ʒ�0S���Rrs%ѵ�ow��R�����j����	[�z4�@%�%I@�'��������Dt��}a�g����o>��~;K%�~���=�d^T��b���;��D!��>q5�$�׿��O�/�r����Lg���cG��JZ �-P���@S����#�"��:�ovÃKW�sD�e���岉�Aw�$�����)��e	�kK`�69�'¹�7�px��W��-����.��p�L�T�ïE#L�Qd�m��L�*-C��.��.�1o^E-�8-�h�O�	}�w�\�i�)lM�!���㺴јy�Ǻr�	hcF�f�|f�@��DD��iz�J?N��6�B_I]��s��l�i��e�������HⰄl,�o�������-5.C�Ӌ	��9�gO���F�:w~F�����A�I�4i�L9�7XC䥄UFUjm>���u$oB�e�� ����Ҋ�ӏA�����ح$<���@ �Ϭ�����-�!�Nh�L]Wp�,'j��D����%��$d�6�j��Qz�c�J����Mg�'�`���}�o[�f�� ���)���Lc��Xl=�@?[�L��4�MD��֊?*��6��A�Ϫ����
?���R�>�	~�,b܈��w�9'��ɼ��w��^�t��p����3���Ơ�#��d�\� ��h���S���3��vd�^���q�9Q`��=8����!9�;L',���5�b�,�N���LR6��~-��iP���8G�%����3G�zGZX�;'䑣6 X:�?u�?�]gl��+/p4��ߓ3���F��xb�dZ��
��㨞>���c8Ѓ?��q��9�#���8㙁4 �s}z����� �>���nx7XN�6|��� =jJzBF�%�r��9�+g����ecrz�?�˻���	�~�o-���h�E�wChY�f�7��/�|y��(���������Pp��)�:n�6}q�O�̖m`S$7�2�k��ٝzr�<Z6F,��=��1p�������ΗL$-���4EBP� �S߀��}ܫ�<L�p�b)�	��?��L��d�M�9M�ch{6�[ߌq���l��\ढJ���D=a{b�"Ϟ�D���5Zd1��H�
�ye�-i!�"�
���xN`�p2
 ��Pm�9 �g�FSR9��Ԡ<��p:^�Yϛi(�5ˋ�1@%��-D�"�&�P+E�<9@l�1%��uVͣb. Z0+G���Y�1i��&�_`ָN{��� /��uLmi�
	Ҍ���`����6r��Tj=K�=��RgB�g���-�[+�&��B����J�bt�Cᔊ��M]/�������rc�XT]k&%�oNDe���t�k�z��^���+dc�%d���=���4�n`�q3L���f��F�q�g�������?w
�,XU&����W�Aw�-�tw�ԥf��T\��K_T�����l��s�y����Ax¦���r��i^C;
����ܗelO�<	�#w��$��hh���u)�Q���#b65�\~�kW�Ԋ���Ȧ��B#�A�́7�2�}�a��'U�#�'x�������iZ�{��y�2;���6	�q�vhx�y���G�����;�Z7���J����l����Bu��Og��������DA��gQ�/x+A��{�ܛ��y���2���3az��d͝�XM�H�u�LΪ��y��Y�!&ܪ@�c�)�;N��1�`��y�9���e���:�E�	������U�����anY�٬���y��e���r�[�����t����f��� ��aE�5���; ���Ȁ�g<��G�0g#��9���$.@�:��K��r>_#��8�kz\T�-�N��d�����P8E�����q���V�Z�X�,n��	��� �Q��M�6*���	�FliC}Gl.��9�5��O�ߺ9^1�v��3�f��>���+�A�ڌF��iJG���=� AsB�Px�4-:��Q�5��k��ss�p�oe�b$K���G���-K<� �;m_��ʲm3���!����Agz�xe>��F�˄
��ȧ�L�@�\{�(���k)�Y��O$h󳯄`.��o�
��/פK0.
;w�o��,�b7��9�i�F��C��`Q�8�*�\ab����|h�oH�T������	\��dʂ84�z.2?I�n2-H�X
��J6��yB{������t	��O-�#Q���,�����=�mp��_k�V���xX%�d�0��&4�k��Dk�OMv��X����eE�7���
Yn���?m�w`�"�k �cT�gX'�� �n�����SW���_�;v���������?_r
V����U!��|�a�s����a��⳵�d�!�F�)�ja���J~b����۾�@��g���Q�00�"�}�+P��0�׭R�_���Q�������!�gj���z�"��=b�m=D
��y���M&��B��~�+B~����H�' 1BR�BJ�y�1�����"�N�ը��}т�`3�d�Ϩ\���N�>@RR�c@") ���U��GR�
g�ƔJ�E���мB��h�\�8r_�F��_Ͱ@rr6����$�n��P1,���h�b�#��;��}��5'e�2\��y/�����}6$�Y��č�(c��y�(܌���u�}.�r}�IQ�� 4ý����M#`qs���]霴��{�M��>�4�#�g������������P/謹7���VC��l���h���U�n����*�u?}G�IW�f����-����ذ�E¤_����f��?��n�����G��1)�U�j,���~KmTܜ¨�#���3�� Oo�y���A���34���`�����r6��w�ǈlʚ��0�cn�����rc>���wb��_�D�W�f<���` =%�6\
��(����ǆ���{��9b��$Ȝ�ZB�v�~k�8
V���}�'��bM�T󬩰��I��2�0�1#��c^z��q��E�z�̓2t����c*�6�I���o����X(�0�&`vg�^����ߘ�z%�䝽��oyJR�����/
o�N��s�~"Y������,۱�;�)q�� ��b��?�rs��,ӣ��f����z6q�ϪpEph7� �׎0��"�B��,���ɗ��3J1�f�H�W/G�Q�ui1�QH�)w8�T�\���ō.��B�_�V|o&4�8��k#ѦgSuF�4������"����e�ܽ��/�gT���Q�j��h�8�,M�~���1٠+BϰEAC������w4��*kMO��(dk��yIj"�96%�����/�L9 �נ��6W�%�|�a��H�ts��\�3�-��N� �9|7�� >�UU�ϕ�f�� �
�����ւ������0צ�{�:#����mc�l� �Up����Y?(o�f�.B�j�p���{�s>c*"�XF�$�W�q��>wI��y��]��-4����-���S��(�[�e�ʘ�n�E�Q�3��gקķ|�6q�lS�VxԸ�������fZ����a`��8lu�<��Q����6�0��Ơ�
�B�I�|x|<!-�V\���f��Ck�Ī�	,p�L�$Ҫ��`6X�f�0�� �x�XvS�0q�)�Y�%r8��ۺs�޲���Qc�J��#x�a���3 <��)L�	u�n�7K"�?s��yS���Zu�i�]�Mg����"���� ����#��hY$c����M�/��%1ݡV�Ɍ�x �������J����?._�e�{
�
=�&P��y�L�hrD��O}p�G((�y�i&���eP����.�1-�W7��Bm
�(�Ľ��(Z`և�"��R͒�����)��E~v��
l��RUr�]��p��@�:���~�$��Q�������|�c�K�g���y�w[�F�k��y�UW�W��})�~���+�F"c�e�@f���XL�Ũ��~��4U�����v� �Nߨt"�^EA�؈�UB_,cߪ�vH����X��ޒa)���"�yix��0/����<�C�-�D5����
�;�i{�:��/hZ1��� �����B\�@`&̰UZ��T��
lJ������[n ��F'>�cyb���۽o=9H�Q-���_E�p���%�WP~ɳ�s5,� �~_S6�Jг��:y��7�T[�&�m���%6��$+��ŕ�(v{�{R��2����:�6�@^��lnFT���ߤ7<�,s��'�RF��+p M̐�gQ,���e^��t;ѳ-�	�}R;��fd
+�� �N�t�eb�A[�yV���P;���BC��a���N�^c�Sh�6����h�~R�ӯk����*�a{CM�j��k/�?��?�t���H?н�����<=��NӮ%�T6�;���R@V�c55�h����4��������kS'�/�g��o&�3#2�v��^��(�5��V�����Z��"7�\'����s9���|�XM��)�ȑ�Ǚ�?��0�^��X�=����X��>�
T�	뗆/���1�[�d@��`6�ёx&#�F����2%�2��śh�.���S���z�Oпd�>���;ΈlM66xp=��PP�&������g��n�)-��OR�	����s4FҢ�>��Y���{E��Ҷ���DX�[� �o\����<��;�d#��6�)�mD����z�]��!m=�KI�3�o]F;�iY#�:{]��q�d� �I�pu��eZ[���6Sy4pN֭�3V�__sa8n������⟪�H��5ޡS|~�!�R���5f�	I��!>{B�F䥥��ee9V���_a��H�G��5"��	~�t룩�&%i�H�>c@���{�ĲDB��=e)�H� x��8�k�3Z����¶k�>.Io2�áL~vA��y����R���7�y��ֶ��j���������:�)-PcK�.u�; �Pс4�%_rA1��������W3(��29�>�Î�����JS����ӓ�q|a�b�^Gy[�-bh��XJ��L�G��O��T�a\Y{F,��^���������J״�+w�e@�=�OvŨ���ev�4MA��!{�.��팚u�b�D۞���Ƌ��m��|�~bt�/���e�������+Eհ��B5��ĸ�Gy��L`���!��z��	�×Ff�(B�}A����Wߴ���n�|���]gAMXm��4������r-�*��-c�'&RAxiT�����bc"sp�1)y�1�Қ(��-��)0§s�G�L$�,(\3�ܖI`�A8�M$�����
�!�h�PukN��7S��WW{XZL��-��Gf�+�w%qVi��Ҳ�V�jb8?Vu*I7����~��o�(�<������ϰ_�m_��3Э��p+���#�/��J����"�2S��*$<|O�͈�a�.7]q����������53߮IgW�����E���\"��l�&;�r���H�h���S!����u=@΢D��~B��,�%����z+���j��9��e!�������	�By��s��dټ��ts����JR�N���Gk��֪f�""E� ��ã^"$��X���t�	1�0�hy��}��d`���ewKԗg�2�&�-�0O޳	���߯����n3~�"�D���N�{���q7�׫��!
�n�r��I��Z�.�}��=C_�%D'�p)���{���1���MY���ز?d!��%/�Hb�f�''�v6T���%y���u I2��[��1��U�ֽ��4R��D��J��҉��d4Vġ�`�&PW��%�0�S\���An&��JhM���Pf��SC�o��Yn��-䙡�<k]�.��F��γKסѭ��Z�1lg��_�o����G/��ޠ<���i!k�N���tv��m�:<0�¡1���JӨ���;7ݡ83�U?y�ҳ�ܖ
�s9���b������I &ԕ4��;��(���n����a�!=�G�K���Ό�� �i�U��3\z�6�ߗ%#_�$	��c�����)uvW2�J��"�H0F*Ò��Wԋ}��NM���c�(�E��=��������S�k��S����}y�B�,�}�b� �o�M�a2�x����TJH�գ�
�Tᱥ�}+��>�%��n�ue=z�k��omy��{J���2�On�Uk����?�i> �A���䜝�"�o�j���ę/,�����)��#��EB�h��"�����+'�"����7m���Ho��k�a|U�Dj�gs�N��G�1��}/��o��J/w%�RG?�+$�}�F7)O�F�5�X��	q��*L��D1����Ԕ�<5"%\rJ�N�~�<��-Χt�"F��R��ܽʛ-��)�y���
�Ĥ�k>�5�MȔl�:�>�NM�a������C:�����Z�Ӡ�hM|V�s�Ä��6����{�<���P�r"�=n��ȏ�K��m�����5��F+b��Z��aP=�K^2����ŋFJ�z�{�#�H�tN{1�Ы�(��~�^+]Uʟ�+du�J\�QKУ�a�_�����"�k
���b��o�q�$��5H<��ٛy<6g��ز�����T1�"���p�(�@!�dC<ȯB"�PB�U9�D�O����	�9�d��I�v��9� �|קx���<a����U�N�.�d8|�) IX�^�/��[$�&�L�тQ��I��h�S}l��[�h%��:�E�6�`�U�㩆�se�S���x#J��T����k�H,IX�z���&6��?�Y���ݱ�7��ӋK�:�^)�L�펫ˡ~^��TWE��NN٧LULX�=WZ��_�3>�/�~��\M�]�$���ng�zH�˰���������+�3M�;!}�5{9�[<���q���ޯ�`W��H�o�����	a=2yD5��jk�QxIv��h�%��>���i��v";X5<�ȰN��A�[>ز���&����{�Re9lC�1 �"��&���E�
��i�C˟#�9���ѱBS/uh��M��@gV~X��Q��wU�͒a=��8�K� �-
e~��P!N.8������F��L�	��j>�b ���2
��R>%ۉtܸ6��?ۮaƆ�é&��p�A+���X���?UK�^��n �)I�%��d��L��ef����K�A�(�Hἲ*���p�Zֱ<�6R�nzx��>��?����t�8@�H((�l.+����<-�����d-���$tS�Th�3+��m8���q�b�r���I"��j���e�׵/6������r��"��Y�6�8����a����ZB�I��B�e0�?x%Mֱ{��8�����c<�@�?�I����_�R:n�H��q?��a����2`�>J�F������c+����|��=���2��RڅJ�o|
R$>���w��yR��!Ԟ)��@s��YB�[� 9D� c�$�lѮa��yԷN�����isd|���0���?f����E����ߌ�Q�9]L�D\�vD	�x��0Jn	��G�	J�%h��K�瘔�3F���C�N<0LWV �.��J��u�4��԰��B�l��Z�һҁk,�.��5K�P�5��W^g�Ր�g�:�w�g�W]� ݴ	�!:�
�ޓE0D��珠Yۦ��^��q�vG�0&��lIC����O�l�݌U��V9Q<��^�Z��AK��ux���՗�쓘Bݓ��ڐ\̆5�վ� 򣵧�䅣�H#�	=��+��m�w�*YNuR���L��*��_q�$ݕIt}��X��':�{h�i�i�3c�%Nߙ�R�U ���"s�u�*������;%�>i��˒���Fm|����a�hACsb^O�a�@�'E"xYd��G����L�HD��d eb��~�gQS�XEK }'��~ٝ�UF�]��!*���Q}��k���`�4�T3/h-%�`R�s?�L(I�<���C�¸�"��Y���8����1��^Q�mC�L�h0�X�/��g��j�h+B'��=E�$�J|���ҹ������į�)�7�F"��va6�k�p��ւސ�T�H��t_� �I��a��P�#Y�#U�+��d���mP�K�K4�U�xy�����9!��)]���/t�y'�w�ɸ-��jy"?�B����X�g���7#�Ozq� _��K��^��Cك9t�{	�Dz����o�Pn��+
XZ�!���޲_��]E�ֈC������2��]><IgĤ����y-)P���v�6.��7��=�c��<�|���v�ν`#�i$�>� ������.ɩ���5D�J��w�a��h'�/�1�^#Tv��lu=�Mq��qi��wE}u�}�S�-)�������-ӧ���^�7��C��X�Ӝ/���t}�G#9�y�{�yB���ۖ�l�2u9���V=�)�J�"R���E�*� �K-[��B�b�:`M���U1�uc�f�`�F�N���&HYE��-篷����[��=H2;Q� �9�u	��Q�BѫxVȜ�1}B?�!F�"���Y���o�W�-��.�V���t&5#�g����-XM��b�4k��iR_�<����Q���X`|	W��g�p�&�`�'�X�2͉��]*����ڲ\��W]�$��~`�������:�	�t~�ƃVB�\o��/� ��I���� ,�F3{��;m���K[�͓U��6'BV�Û�_��՛�h�6ߝ�/�܎;rxC����S���\cgQ3~ ��[��	x�����1cZ��Ŭ��6�0�-�����K�C���H4�X�5��y�T���QI��*���KmpY�P#�5��I�[������[!����*�^�Ew̦U�O�h�n���u�f��� E����<4L������:��n�$ީ����X���M��9��C�t����`n'F{0�Rʪ��s���3Y�ֱ�����ʩqc�L�#f��2W�/����i�P�������#52������D��H"QQVA$�"c�7qt�#K��L�(z$��6�mћ��*d�C��v�6nLa 1eظ�+3�d�_$ 1��`i�!��)�ma��s�~�YQ�>��B�N�)p���'��,���DTc��*�y�`)�t��Y�8��MleO�T\5��Dڇ[>��m�����^��'�ѓ�"]TOd ��ĉE����0 د\����HßM�pGI�*X�8�Fq��Y�c�����hg�r�6/u��TP���j��q(1�/P�!%1�v�'��
����}>�%K"�b�z����7��ݴ��׭CB�eJ�V�@7?�S+����h=̏F�Q5ε�p�����R"�uD�I8����.�=�\݌{(��"�0-��ܵ�jZ>|�Z�+k�T� ��9�X�c5�J^4�Z"'\�q�Z��-(A�-���r"���_	�嚗���g�Q���l���6�Vҕ����X8��hĞ@+����5,nB.X��<a�T��"��?Ƈ����w,{S���>��go�o�(�
�B�����W� �G^����M����"�u~�Ҙ	�`o0���=_��|o�u@�K'�X�+�����Rsϰg� M�x�B�T;)� KL� u�-�NɣHM~]�|�#W�e?���5{|f�%�����q�:cHj��P�e�<���:�e��i����E�����eώ������x|���M:�	eap��1�A����Y ��kk��ut�I8P21�ȇU���\���4�_F
��)i80��Z:[B�/������5��"��iJd�t��������\"|�q�i�SN\�����һ�m�Ų�Dvn��4_0v�/�����hc?8qb&\p���7�4{.+<�w+�e��DYKϢ
�n�	{|�!>��Z���ݘq0�'弝�ɔ��}��i�a2��R���Wvb��U����X k��V�/�󯔀�?f�D\��'�Il��k64J@� �^��6i��)9}ְ�-"Ҹ���j���\
��5څ��$ �b�����p�sAS�Ri�fU�j9��igi�j?�M=.|�|�����_�)�;���� M��h'ǰz�M�LG@&#���~�r ������q�C|�����P2 �JOT�Y6��0�EM����7�i���W�`C2!��陙T�I��2�r��%����]��3Ǌ�X��wBFE2�`+\�ӄh�溑+�8�5�p��Q���Q�M: ֮��:�"���ͦ���:z^� w�j�I�?GY�hz�^����v,�h̝�%���3�ѱ�������:��`{^(,~E$.���)���|�]-�D��+�L�;���R{�A�c��C>��^Hd���	�L]A�}T3O$�ʋ'b�tQm����nw̾Z9�r��B{�,.y��E\����q}��)_�>8����^�	k"��"��:Ib>����O�c�x�r~�>#&L;5w$��= ��r�����X��]RpޘD����^~]�ǁ���A�(�"�-(L����@]�����GxO	F")�P����굜	�,�]��R�/Lb�puE�_�xk̒��>��� ے�N��v(ہ�TЕ�گ:e�/#�$�e�ʮ�=��t���#�ﾅ(��muq[�}Q�2�3k1oL*cp�v�H��1S��R�U5%!�Cjuđ����r�}�>��/�h(I;��i6� ����C��A��,�c��7�o�����M{��m�(0���"�O2fZRM#�4��P�)� ������Nhp6�J��=��m:"� xȶ3��2�YT���z�s����_����,lw�Q�X�"a�chN�� ~S{�[=���K0����Ѷ��C)ԯ���8��'Ś���<�3��dZ��~=�xE�N��"�ͳٱ'!�i�9g�5mB�Χ�1Cw�����G��Uɞ��Y;&��纣�Y8I�����0���q5�ja���>uIǷ	�����h��Uή.,a�L>����s��-_e�jy$@��B�Y!Fل�s8o��I�[�	f��C��G�i����l|i����d��������jR��#�����^�a����h����&��8]'��E�lY"�|]i]"ӽ9�F��'C-z��L���X.���=��s���o��7����u���� $>���&w�?d[I%�&d˛��E�!�l�f�����Ya��6�/ղ���9�
g�[��rW�km���ar���iw�N �E��=�#�&��/5�ů� X��K�E��t-e�"�jI!�X	<���eS�ob�� �vn�)�����y ~b�YS~}����2F%w��d罛�]l~��'D�z��xc(A�-�/��%�
`��BO%�|V���d62���؇���