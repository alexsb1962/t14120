��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����F.��^KN|6+��X�Rs��Be�m�.H��Ld5�g�X���3hUW�E��rbϮ��8�e����.z/���%�3%���y�%J��/Ơ:~��������D+���o�֞�����`9�2i�	mKbOh�� �\Nu�2J[��F�Ƹ/����R����x:RbЁ3�������0KQ�cu�� !X�֧��o&K�����1�>}ժU��(�`���BZɿa���8��s����?�cI��5I$]�m>+�J�Ce�{Bb7�Ե1c�u6�}�D�o��+�r3֒�̠��;����h�-C�C�/�~��cL6/��e��v|A,;H��o=��=����	[�M������Q��� ۹6�� h_�o5�Bɋ�vU���,��p�f���f@S�І�*l�$V�J;����+z�;����ޕ�i��Kw)�0�n�R�BP��3Էɏ�`����!0@@h�e��p�"��U`�k���y�L�.֬t>�Vi°�._�u��oFS_ ��e��IP���|���	�D�Z�X��r�H/�?5.����8�8���U?l���(bΛ�g�E�|����a��}:;�R�j �}�i;�fr�o�*ɩ]}�n*�{7�3�m��Y��Y|�p+Ê���*�c���x��X�ƭ����uvm.��8���A"�AM�c��`�G �g���0�'�pڜ�~u���{�4Q�G��E�y��J�D��������l����r!���x�z_w����~hZ_^�{��R�.I٨T=`s�Hj-�0�>���
U���VƖX��C�O!�W�W�G���GֶA���i���Ӥk�J\���G-A;�R��N��z��&}�V�A�NZ�tKPf���&�7^	x��s�Z@�|!h�J%�,�=i������l����"ӂ�m��M�N)�^B�9��	�*N%��T�ȼ&X:b^o�ep�/�ȃ
��`֡h�{�\΁.=f|&m��*z4�~�߹��Zy�#@[RU6Mn�&R�=�?��oa<�J��Q�Xߩ�Y����9��;ȧѮ�O���u��x&��'�s�ͪ"W�z�0Ԥn���P}(��c1gУLE���54���^����.�$v�䀋��n?�{+�z�l�V�	8VG1��p{��擛���?r�O����s���C@acZ��!��zXl�ŽtZ��ʃ��ԧ�8�����Y"̀7�	+h���\��X���0��8�P��"�����~�h�=�vv���ع�(�$W|��K��q�:,=��,�P7�΄Z�d�eũX�r&������1��wc����S�U�҈��98���̷/ǉO�'�/�-nEz����*f��!J��5-#�������҄ g� ���� ��[Rb� ������|Dk�q��(9�\i�բ�����w�z����F­�<3+ �� l�j�X�c�h/��r[y ҟg!I:�������ǉ�rvDA�(62��{��=D��d�8�棈Y� UlE2oP��&�Р
 Q��&r�!�7�&|̅'G�נ8n�)����B�s)F�Ҽ�r�T���/��S��.���`n7����=����rȉ�0��7�@H�	�D��shz���+�h���A����r��*1�(���rE��M����T��^��Vٱ ��zO(���]��	Q0�<����������&��n�GFPp��D�A�[�j�?*�ʛ4��:�Pg�~�-�4����ѯ/hsH\����'-_V_�]�ϸBè~�����5�q1hٳ���s�`D���]���2?����ٸ�fS�L���{}������Z���#�9$���3���gw�F&��]X�
�D�x K�e�^�RP�7@#��yq�Q������
�]�tDwt�C��h���:�ڟ�� ~R��O*_ǖ�$�]Œ7|�7"�Q�� �K�vVQ���d.z���?]:맰���外cT,�Sp�o+�~��
����g�a�Ȓ�i����~��Gn/P"���:v�$�^�D�˞�Xwr��k���P�bbak�PVX*�q�� 4���2��[V���;r���]c�gV�+�~��g���$�ͪ�4H���s��;?������=ֹ
$.Mנ`��;J�^'i�"�y\vA�@��,'�'��� �[C��]}$Cq��/m�r�Z�k�ޒ�Ѿ�Qfuy������_��N�i/��V�T���KT$�)����Uv���>�Q�Ր%6("D�}�����)�U���~�:�եe���V��&�0��%�'���oׁQ�jj��\.5wE����iKb�ds���8�����8oR-�Q��o8~:\�y�:��@�q+�3e�}��8� �A�4"+l��꼵��TB�*�t͘� ��W4��na��wv��:��5�� ^�Ӟ;��j�����n?�=j~y�AH��C<� ��:c��љ�8"	y�MP�D��I?=,٘�v��)�U	�+K��'�uM���g�:�o6rD"�(�f���w&1��ynM4� �5�np�N,�ۀ���FN��W7uC0�7)�T|�T���-)��۟�dȺ��S�/�?r�PA@X�<�n%β�k����I}]5;��@"�?o	�~��2�1����}9z��x�8���g[��%��ȹ'E��T{���c~�5�+4)f�r@%?"��;ɠ��N���+*2?����e�nN�|n!n'K L��L.��N�V_w����*`8�6��Z�LC������I�:�*�@j���K��z���#ڡKL|���B��?���W������y+Ğ*� p)c,�$�W�r���
�`0\��L�lN�C��K83:p�	��NE��l��Wi;o֝;����ǷlM^�ei��;�$hѲa���G Ʌ���,��E�e$R�*�5�Nx�_��܃�:�"�ƨUCK�G���Ob��Q?�vT��6��7�ϳ�9�m�w��L��D���<$s�˴i��|y��������c뙁 �N��F��&�Y^+�bg��Z0	=����� t���J墎�4�#N��K�A�D��� �[5�[I`d�E'��ͥ�ҷ|�V�JD�,����/G3)�o�Fѻ�4/v�G���#i*<��q،�[.��uܥ��C�c�����IT��7����DF�גT��Hzv��@���m�4�V`�l�񯎾��@iA\kԳ�����uY�֞�Qq�����?�����D|2�c$�v-���؎oց=~�g^g�if!�(�sM�`b0�r\-�
tp�~l�W�D��6L�5��<,��G����sp�٢@v������Q"�k<J?{뼼U���;�� Τ��_����5�����<_A?�
����_"����!X�=������(}Ɩ�(��mf6�Є��K�޲��ė|0M�1}K��	����P-б�������n���|�W�t
lD���!u\��k��RH����ѫ�WCm�\gyy�Vs�;jg)/�j3Qj_S��(���4��r�j�[����#�TH4%��=�ڻ��N2sq��4)�FN����8��6?����m�ޙ����S4�o||�V�	�3"z+��y�̍�]�*�M��W�̭�մ80���0w����t�����4��츔E���)�;�`fƽ�Ȟ���e���j�ycւ��5b�}���z�q�M�W׫�/$_@G%b��ܕԝn�`~���� ��}�C������򈘸����.]Yன��H��+��
&G�k�"c{C"t
u��<e� ���t���	 [t�5� �4g��^�*'�~�XRc�U�XX��݄(b�[??�x�����7`��9���=���34�d߷ �uؐ.��.���!f[��|_B������V`�s`ɉ>��!Q��[�*¿{�_�;��Z9�33[ܾ��w�!w����}��D��R��k�ԥ	`{�P\�d�#�ʞ�`�nR����!�ՏG�g��j�
77vsA��Bm��}ϡ69����F�4;���1�h�@n
��^L��9�<T#ߠkF^M��
��/���0[��l"F�^�MyƛTRY^
��ߙ��^6�M�u���[2���<�
%��D�H�6���NZ���~}Z�Y
6q��؇��[��5�p�U���5�[�ӌ:�إ-�#�g��48<�������N�H������C����g��qe���Ƚg{*�A�e�X����ƞ���BAJs޼�M��0n���jqh.Ƽ4
�ǉ�΂��@�~��Q�ܭ`����D����B���DO�R|0$� י5���4�:��2	���NG<�\`��	tF�{�?/�i`�S�o5l�`R��B&;���rj��v���kO#[{/G��Z�ڙdw<sp�h��S`h^��|�t��Yi�^�~S#�?	��Pn��[���>�F��Bs�����Œ���xhM.��?�`�#k��"���-g��x|�0A��o��I��+="���0�����o`�9د�:%'
��a9��(W&�!�A횼��[�G�GWs��G�5Օ��\l�x�É�G {藛�U۝O����~g�dH�Z8��G��= tW)�W���!�]ҵ��7��U��
�(Qi������4Vs��@�/�HL���ɕ�\�a�n$]I����%�J>e�a��t���U��A��۲{Kd�c&�k>�
��s�}��Dդ:��I�1�F�O��"!�l�w@[��p/a��dۄ*�����i-�FB����&l5���ԡ��<�$o������8��(�GE䮙UMH��R�V��TcN�)q-�yٰ���Ч�OA�p��͗r-SŲ���/�����5`:���Al���?���^XP�K�l�K�=����`_Ǒ��6n��S� o_:��A|C��@M(�� hxv.hX�Ū��_���:�i
�o8��֙�XBSI���R�3��H�0��P��p�ɮQ%�B�ex�{m,���4��iE�d�*O&�|\����k/04��Gx��=��/��,8�:�(�[
ZY�@ٱm��j��������҈��껣���U�z���������s� ֈo떱J�m3��x�ծ���'U;��:�����*��8�j'I�yN�:(a5?�u��n���&�%|�F[@�<ٳ2^�B�}%��`&�DDIꭹ����Vv:-�2r��u��1�m��{�#H��y��^�
:����n*86��YĈ�w�v�{��7��
���O�n?�~�fIR�m�9oYuf��ɦ�y_��"<k*UKH�dM���~l)z�!� PJ�Syd/1�~9��c(� ��������+nE����mF�|�'ٯ�w2�K�Q��c����̏�nm�9kP��!xh���kR�q�5�a�c_�q#a��������e�Ց��ѿ�I�q�T����,�-6/w��o0_K5p�D'
߲uꤙ���-��4mM�v��y]I���;����@$�EʱRj�z�-��[��!YPBW7�J�M�Ww���gTZ�q\���ᾊ3;~\���U7�^�t�*q��3wYj{ńI^��Q���x�"CNz�gnK	Wyӈ�~p&2�XR,DwZꊩIH
͌�u1���:&� g�|SF5�s��}�.�=�i���"0z��b�0������)�Rd�V�b����76ү��;����4x��DbH�L!�L��f
,�&{>�<��E�|��<�/��������1F�x�V�D\R�,��NM%LIo�h�%s0DWz.�F�P~�E*��oV��ڼZt%��O	V4FH��l�U�7�f���t`��<1xj*"<+��:�֦����F��?'�¶��]��u�FZR�)�g�I��v�(i�� ����P��|S���Q��'�n����T�	�|��l��#�l+�����w�*ɚ�:��Z<Y��Xe��b3i-&1ΝR��	���:�d,R��q���%�W�РY��n#��>\��[��a���-�X+�;���d��'ˬD�ݸr�A���Jѯr����Bv8j7�/��s ����tQjX2ruC$&/�l0��@:5�H:2��sYq��E��V�xm��*���C:�3pʧ[]�7��_�w��;Utsk)26* �"��h_P��s�Jp��c� L��h��HRw$J�+v!��+!�!�����80�)|o�L�q'�V�ay�[߿���j���hwt�r����l������~
`�?�	����I�8h�~���[���l䎅�'�A���O��|J���Z�֞������b��J�]̦4�G
�AeЀ�āX{��h�i$�Z�g���P�>�J��۾��Q*��͞-O1�Ir<��R���n�~��K�����k��X$�nB��c��()�8��C`m�o���H+ �wRBs)�M,�N�I��K'ü��A4���1�ݳ#����*�;.	!�Trp��R�z`�~F�=��?2��C�@���B(�<a���ݯ?S�!{�y�����mO�� �Y|��w��ή�L궾�\MJ�S$Ԥ��9џފ��0��ΉS#��o�N�6����l�iSD@|�m��I�o�a�ۺ~uq'HT�a��Վ���4�k~l �O�^���g_�pzъV�PӉr+�b�[�{���.Z��%m�$�ɲ��~M�bIw$�`nN}�D5u�L������/ ��xB���-���G���ĕl=�ĩ���%�ʵ�&�&��Ɩρ��3��PR�b�0�&��R������X�9Åq�璇Z���P��=sVEcΖ����{��2���Z�E[1CWƎ�zywL��}FO:�&IO�:�alv,c�W��Gtf.��]�iDȦ��_r<�9+�mH|�؟���O���Τ��yT8��U��R�u�$��>`a�O�B�>�vR�[���*6�&*��{> �}�'���M���ߖޔ�,�i���q��YY��ts�Zb���2$!�5~�+����F���NC�z�.`GO�'r	t��V}��
�C^pm�a�y+�����`{���#i�@�:ފ�:��W��3�B5��5�;@����v�f|A�A�+�a���+�i�e��?�U ���rZ��k�G��̗����ٍE����]K�sp�O�����]T�A5�����5!��9����A�%�xJVv�	3�9�ObL����T*_;��&i?��A� �Ǽ�]�h�p��l�^ׄ�~��
��V����-�%�1�u������������<.�H��A�b*�!`¥+ ܓ"���]��KkI�����5m���ڧ�鱤�~�����9�K�����W=m����Ng!�
_��:7�6 3O/�~ި����U(��Tu(��A�Ӌ�t�XO{˯P"�����*����9LQPKP��#��5	��}�4(��r2�$��>Są/�O��6k�d��m8+�N��X�&�_�&oZӌ~F{���9<�E�r�%�+�c�I7[#�>�;���%�u�{��/��>W't�OHtb p�������$���5;�߸yG|�yǒ�;>3V�[]E���`���w�t�i��{�ㇰ��9Dd	W\Sg��൚D���:&v7���2|q������p�8�6j���fE䤺��f)؂U��g���ۘ�c^�=��� G�u��)~ju����9��x�K���mP��Y�gi�;à/��R��U���[��`�޶�eWt]A��Z����'�8��L�XLʏ�y�ŀ���YjT��*�����r��\!��3T�+����~8DM�7HS�-8��O����fE�yS����Gi7Gܔ���U��;�y����B �W�b*1�\�9��m�����Ke�w�ڭ=ZYi+sL�ݴF���c���`+�:j
B \[�G���߼��]{w�����SS�R.���O����v��"U��#49�y�i-�+�(����R�E�Eg��}HJ��)���o5T��Tx�?۷vg�D�70朎�"͛�7��zi
����}gҺ�?��%px'�,}V0���f�Vvy$���3��<��US1�N����q�,��π}�h�>z�M5��F��i��+n�͡��"-b�����uR��y�Y�Ɯ�7!/;�E�X�(�QA�Lbz�'xj̰e���-�����#�\��I���DyJ-��&^�R�����=�n����RS�*e��������� �v��M'���L:���ĝ�$~����ef9�˔��1��j��d0������/=*��j�Y`�T�!V"�)	L�+���@�͇"��zI:V����b&!�9�tG�*hw����I�z"�з�5��"}���	��C��
\�(��M	\�K_�r犧A7�l{��A��n�:X$FڵO����Hk����װv�0�h��k��>a؅KAY�5��-��7�\ƚ)���)I����'�k@��>#�Q���U�/:��0/�����z���";B�����S�yk���;.9�Qz�.n�8�����9ܿ�,]�Y.�NXNx���ȷ 0�v�-�\�d$��!aޠ�!<i�o*�9{�'Z&(�%�z ����c�v�"YX,_*	�=M0�P5���d�:�X�@D�BM�~�W�v|�/�l���)?��w���'.2yt4� ��l�z�
 I�,� +�9�����'Z�W4���2�*����Rb�ժ�(8���`��I%aIѩj�ݛP���P��]K�q�v��gC��T�`;�Q��l���3m1�û�h�omh_�>O7J�Z���)*�p�~b�X�	�2��|���y�=�(���>?#�}ʚ�&0�B�{��N����yD3�W�`i�Ѝ��s���YW2�����7g�luF��e��[L5�$/��2x� z9�*[���gNU��Nj�*����St�w��E���Hָ,4J�ē�K� '�ټ
u�8���Ckp�m�]�Y�f+���~6�
7M��	�1E u)�}_�"?ߚ��Z��B_���c0�*HjÑ�9(�>e�)���p��ݫf�-e�U=k��?��^M�/�@�f}&`�S�d�E�ҟჃ�!ya��|���J'��;3b�_�d��z�|&S�� OPM��4�߅��ï���g3@�:<htiF���Pf�c�^%�"s�pe��H��h����J����!��pK��bO
lѾ�ʓ%�vc���k���h��_ �#�se��p���c�_��F�"�;"�6���s</�cd���;&O�Tr�T���y��U��{�3�O8�ai�����f��]�&�b6t�H�>@��b�;<zO��b��ƾ#HYs�1��t���yz&�4ԺD>�+L�
�2�@��B��M2;��_��t�5�Q��)��&:��|䕑3Z�"!�"~Y�U.�Ӣnw�W��y�B�L%`��A֟vIX�0���@���&�v%-"�6S�$��H�I$����+��G�3YK����FF�S����s�Ll�8F�p��9���cVy}샸(,+�W����Xt��0N��"�Y���-���dc�ImPxb�č������U#�M
jāf�0���N[\�R�P$/V<���E�T��!R�/���\h�1�P�s��X9��6�p��|d���@%����G�}�,-j�㑞1�t��Y[��M��� ��nm���A��U͠崍��Q��b��r�N�̀�O�`7EHd�c���m��Q�ޥ�?���%�Mn�T 3���Tm���aA����_�RS�_=���@�/,��k���)�˜��t1���El24�cx Oe��}}�s.��V�^���ϻ6�{��N���.J˅�OW����»e��>*���6�ƙ�HM��N�?��!�>�=��ES�
�|U�(j@6mu���i	��o��LKB������$eTР�f��������T��Ζ$���B8��Cn)��<%�)��!0j�ˈ#w`��i��8j� ���"����"��I]x��'��S�!�sv�0+ DDJ�kT]��[��K�LA��0f@j�����&,m����i���s�j����.S	8�YE��V~��:RW�i`�+#�ā;7���F�,�P �/�Ck���k��Ydk�ܖp��(`��?�,���>��_ ,;�{\ݥ u�BV��Ӷ��[� ��1��m��~,��#�V��g߷����]c��4�� ������R� �̮�K��Fµ3�!�C
y[T
�'&O���.��N���[���?܁oi֓�7�9���5�pE����g�>e�/�T�e10���ۍ�J��+
/O�B��Lv�[�\��lԂFu(�)�v�̕���	Gh�r�L�qeq&i_b�ޢ��\�q��!X̖��M��*��B���K)�E�s��i�o��&��9�)�4��Gbو��D�ߏ���Qx�،��څq��q2�Z�����K���2�3r���n%H��o_%��fїN�m�'+�!GFѡK�<��<�c瘧}\�_A��.���3���f�ND�j�iwk��o��ړ����φqw�rKp��^O��*�L1ZG�[V�T�;)�ĊXW9�k3\I�"�w��%8<Z�F�+G� q������13$�lq�Xj���0�U���$����2d�z	QV"@� � 08X.m�V0(u͉��t��JkO�b���HP���V b:��/�a�zR��¿q��Ns.�k����iJ����`���&Br�CNx��X?�����K�r����3�����,I[9%�㹤յ��Z�[�k���1�?vE��hK2�J�s[���Z�� /[Ҕ1�s��|G��]�.C�?�f����Lu���E�%���T� ����O��2���-#�f;U5�s�nd��ąs�a4DۃH��q4.> }oB0��r3[V���AaK�����y�:(��_�����,j w��ko>���/����O{