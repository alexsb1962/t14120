��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����ߑ��#��2
8+������w�k;��B!����DP�zF
�Y	���7�,��$\�%��'j:��FAԧ�VUWk�7�T/<��E)����7�d(s��������1�ж2@�	���͌�s��3��v�C�f�H94q��*�<�a�5���KcV�v�	mpz�&�J|[�Np��i�ֹw)4$�c��1��Jc�	��qxl���`9�����̗�v
�"����/J�
5��-�jQ�osُa
������v���G}EԽ�!�F�.4�L�0��Ft��ˢ<��W�,���me0�� �AO�쒨�<����L��I{Ce9�R�w�;$)�nQ�x����_�Ѳr���M�)��� ��k<����ABS��տi������~�����]��m�k��,������j!�@�F�?N�)��V��j�/6^I��H]�Q]���>ʮ9f�	E�l��k�o�"Ұh�A���7�F�<t�ܔ�9�M�Ld�3�58����r������4U��&��KS��rҴ�k��/���#���8{mQ�3G{c.���y;�l��.�Rҷ9��<|�Aٓz�Tu�i,��`5yR�5�/��C� C���T;�9�*�o�n�Ǉ�#S_ ��T�ė�j�sy�Wa^��^���Em~����h�%�~�W��9,��/�P1��`FH�lvݟB)�ӓ�Un�5���v����E�Bż�z6�l��s&ϊd+�E|Y��g�Ш���v5�T��EC	k�6����Z�v������5�H7G5)��Q�'���B��:�BS֙���'b������a�R�d��zk�Ġ�;�Uٍ�}(q�[�KG���@��<�|C�~J�lqVӔ�.Z�!�3���u��{\�gc���$6YV&�!1��|	��z,�T�9隫ǃm���h�y��D`W�{7UW���U����/�4���q_'�� ��{*z�aM������t���[8<h�ws�S<q�A�9o �9i3�ul|��}Z��4��<8�fr�r��i��OH)��+�G4�I���,W�����;����o��҅�Y�+�cCw��O=K�.A&uJ�n�zh�5.n��O����C_��r�����'�_�fC���BO=��/鉰hq��2�I��gMQ[Av�z� VU7_ ��`�h���gI��I^s�'�T?����`�"6���ON�-�d�Î4H�r~X����O�_J�tߺ�7�\屰�L���B��8�hW�l���Z��|;�PJ=8P��<4��+�9����48�������{����s_$�^D��a�� '����v~iC�9�K���+-OA��Z���dC9��wc��y��֬��۬�G΅0#�3�X�B�L�w�'�VE�������N�|.�篟=_��7��Խ��b<� 2��D��I��|ؖG��,��8��[��ǎ�� J��e��9ՠ�Q��~%���"<dx��z�)�\�.��-_��Osb���p�ԏJ�W��|E���䞽�js����A+39)e��9�z
:B���c���x��V�*~p��E��L�}#s�G��GO�����O����Y9_�׳���II_P���6��
�~�+Q`[�^"���\���q��{��f�K��$Y���Z�ֱ�����*륔77t�����ya�[����M(x����1�q�VKO�k�`PAl��Gj��u�]��9�+AT1%ú�������6��e#�|�4��7�׳�]dh����2@��є�G<�I#&xr�Q�cZ�φ����#;4�c�CP����i���>�O��$5ȉ��`m��ܗ�
^��N��#ݻE��
5�tf��i3:��'%�j��ϗ��LTS�zUD^*���C�=���N8H�rbj2��u�ֱV�õ�ʵBS��=����F1v���h3ו�Z׸�e�=��h��I�H�>�I�8R�U�w���q���֨P�8�\��~��a;�}1�"N�mA�ƥ�熩�d0�l���D�M�W���Io���'[��2j�:i)%A�򓩒�h3����`\��=n�ڥuW��tz�6]w`�!;@�Ly�ac�G��^�l�&Ē�M>o!4��EL��a~�o�,����r�j�u�c��6{�#j��P����,�2�	�
����D/n�a�LQ�&D����@Q��&��Tw�m�@�3�0���?�6��M���]�����ם�Ek<x^r���uP�����l�0��>5r�w4b�T�Tߨ#&]�_�q�K��p+u�m��V�����g.5y+>�!���C�ūX8X��ujs��Or��`:���Y���[��`������~=L�A"��>�8gaeƺ6�Kb3?}���{4��0�K'��MP�y�;)&x����E��l�>K���{�z�n���dݼ�e�{W���.�
�'pvؖy���'�1��6�L��@�B�v�[-O3�X���^y����%zL�Z��_�{j���3���s���ln�PƗQ9M0�-T��m3GD1��g��i�jtw�,{�	�c��ő0ý��-�k���zS{Gչs��]P����g�>�pP�� z�f�A����wd�p��أ�%-�b���B\�+-5�(�j��{Ŭ���	x��8��-6Zf}d9�n��dcr���!�*@f63��(C
�K5�^�翯���lgoظ�Ĝ����IS�/���y�ڨ�V7&sn�G��ɠ��ln!u�a�k�y���w�wV�YJ6�����4
�-�y��KK�$�Ca��N��Q!Ý&'e'0�zQ/��|��g��<=��-��bmf�����N�A��Rq�v��#�E6�f��|Aqr�&�+��e�[B���`h[�i��B���eP��T���l�y�'�2���S?�ύ	�|�*[|Z8Y7�H����Y!/%㿾�Y�;����3|u̡_Xp��3Qx����sEf�l���='�To�g�� �pB=J��q5z㹊�`�x=���T.�	��Ps�H`�iY����,o%n�㧁��IP�҇叨��c�8�s���o��H�(�����W�8?L�������j7�@�P�^��AY�	��m�`�_�����,����m>�����Ƥ�##`���i-7}� ��Jyy���O���=e��&F	)n�P��ڶ�W��w��Үţ�z�H��[���*M\y�.��ۂ���oX}E��0����Bt� (��O���yy�}����Uw����io!�I�d���q�2���u�~K�d�q��.vj]�٥<��S<Vv�I�&�񈧮�&�y����ȓb����_8V�Q려 ��y\)SG��#�"���?s#�b�k��FW2hJ�r	/
&��*ݢy"��B��nS��e����5ˬ]*��U�V��do�g: +`�3 ��]gY��-S��Sd$ZxsMY.��P��^՝�8��C-�FЇ#K=��7��D�b���?�N��ɣb<���H{Qzvr�ըH��p�rzDZ��(�7a@�%8]t�?�v-����/jE���hp�@�Q~����1y���G%3@&�Y�7>�i`�ӣ.��f��o(�g3�14��c��_B�G:�?�A�7D �����J{���#�=�-F�g��Њc��Ŕ�e��d�SW[�F��zSAc�E�"�����RGj�͞�K��M�>��V�N�P�y�2]J'�
)s�e�$�K���',Q��E�T#>��Qb�!$�F��l1X��OF.T�^�	��<�U,�_I�7�R!��b���/��1v[�b [A/?2˰"ݧ#�^��s��Qei��F��y;��H}�V�����jc�h}z��1l[�������Xj2�S� ��*6��뀾|h%�dZ#�'>˙->�+�J�8	C���)Kt�s��9�l��Ǌs�t�{B0>��;�Sm0z 2�� �����;`�#�+����2k��}�0��˛������r��-��<㞳K�|�^2`���?�;��1T������3��u�5Ы+��(ƔL��y�X,B�"��D��R�kg�\)��x�{w�m{i+*S�<��b��҉��g��u�p�>\Ϸ����3�?S���F���T���>i�"�Wv�:6�Z�_�	�/������v�e���l��ʖ��P>I���ԭgN}}K��r*��1/���@���A*ImĽPI*�f[����V�;ֈV�]�u����z�a ?�O���J$�)/ �Ylv�-�����N���u�S�I�[�˗�����Pn_�kQ��b�|��Y'��[�W�%���@�o��W~s���?���� �YRT��g<�/�c$2�P�>]�G�'�V�3`�E�~{��^!Z����Ic�M� �����N���묜�
���!�n�աVN��C�d��I,�Ƚ-�p�'<����4K�E#xZ@QƪY�J] �Qmp%�oq���9nֶ/ߐC,+ ���j����7>����*�13���s�vx���ylhZ�.�I����M!f�XX��We�ᇂ�:�_Ƀ�jP��^�v�;��kv�Z�1+!6�������Y�gdq���s�JV;�i/s����@7��Ȇ���nI�;��2[��<�Qj��s���To�6ӧP���ӧ��X�QN����W񺦼�Yz��!{���ꂓ��/�&hwM#� JWn�Dzg����J<�Dy��	�F�cq���(���T�wBRYW���bG�	?�HP,���'���Z�x:�o�~Ii�e+����am�O�JK�P�d?��Xy�t�j M�bf��6�����|�-��@�Szc),���,X�m�Į�g�S�<���k��6b�Y(�m� �H_ʷh1��-ء�{��v�<�[���ɭ9F�',Ϸ*�Ϋ�8'�2���q�8V�
r�6Zk�}�4��@\��mR����[��c�o_��� ��w�'�!�F�}���0�.g�z�
ן��gS=9�������"I�����r��cs�������<�z�]��F�v����
�ɲ��騞}N螅��ՄND�#�,U�����Y�� A@$_V��wʷdw^x���K��:�u�G6)O��+\b��+�!G]4�.�*d^D{�Ѕj�jN�����k+��[�&���V�������˛��\�b_n=�M*{����|j��q:&�pM2�%�LW['��i�;�����$*!}�w��c�.�qB�����N���~!TÌg�̤�5��0t�9� �>KK'*���6T�Tyߠ̫"����n��J�l�\c��	/�Y0��S�f�%��z�:1�컇���)u4�X�F�w���I���S���3+�\-���No� �q1��s��'П�뻎1�׀4h�f��xU�����e���h� d��hbM������� ���Lbi���	�9[���h����>�k�_kM#�+�y��A�? v�������pT��f���l&�����@&Xi4�	I�{ޘ�P)��ە����/��or���3&4VH��η dy3Fss��`���	��@��T�躳����W��J]�g^�X�2T�Ahr<q-�Ga�����8����|m�z����_%��#�h����YU�dI�+1�t��%�7�~ ��`����v^չ'}=�g�S1�J��<AH8	� �	;��yPg�=z��sb��C;|`�����B���0l�\�Ǡצ5����:uN�ߢ1�v���b������I��1�|�V�kAű���sRyߤ�E���Y#=X�k0�a৳���x[�3Hj
��	1�*3��5v�m,�u1`��؋�XgJd�F��Ç�L����5*�_%�
�t�c̔��9J*�n�)�T|��n�!T�r�'��sPm�es��_�˙��ODܒ���b�虦���ҡ8i��p6�r7�%y������b[����r�>o�O`���I�GZg{�?,f�1S�t��FY|D�i�Xpod���~M�&L������(�qe�D-�*�|	��>��V�� ����I���O ᰥ�zqI��Ms<'��9��\U��cH�͝�$Q�T��'ł+�;��0H��~�:'�9��3x��5�w: ��ch��QE��լ��uCFW�6�~R��)�����j�{I�Vmd����t��o�P�6I`�q6f�[t��ro������m�wX�n�`!��UI�? 1W�j��xK�H�XL�ޖ������D�Æ�0�W��8=�,
������ ��H��M+GkN=����/sH8��l$� ��[�(�#�qk��V��H�-⦛n������JN��b�!b"{�l*�/�r���/��?ڷ{!�P%G��}�K�\��\����xٴg�l�DzC�����e�_?']\*�����Ș��aCf�����D#�Y�P�m� ���&�O E[1m��GQk�7s������K��$%���P�?�4F"Ik�Idҍ	f�{�^���zT�G��k��F�|�=�tb�.��P��(:H���`s$v�YK��R�4Ț��_�m[p��p�L;�[� ґ���,O��1�wzx������F ���1�Z��p{�����KS�>���R���?�R�z���SuՓ�Q'�7y�ޔ���(�ɒ��_���}iQR���C��������t~�Sj�T��{�H��DF|VWf=
K&�t�]AA~��q�<xK���fI_aj/�B��û0���<�x0�ga�Fބ���>y�~ry%c��Fn!S��=�~�C�쐵lh���G��ٟ�@��.N�0n���
`��¼���(��/b �6s=D����z+��6�仜]�v�'w�sr^j��r_Z�eV�A�~������dՓ0�����tG4�ү�g�a_d�Cj��-y��:�N/��
Y�G�� E�xpw@�f���X`��U��O��:<sC�7E�H^��ٳ&��6�k�>����JY�V�\X�l5Q��B�9�(����m�6��(q�a�=G"�v����x~�� Ș�鹧������u��QB��0~=Hš2�gt3f:�Qo�WֿV��QvLZ�A�?COw-��]^�n���F��bVV�9(���s�rt�Jܼ�H���� /��s+���	$Y�Ub	��{=^(�
���������vGe:�js))"���ʆ���<Ay4��ma�0�4BB��sR�,C�<�2�(�C��x$�`] ��z��Ic,a��M���N���E27;Je�Ů��\���l�x��tg�XI����0��E��<�x�61��ȕ�F]�u�~C���VHFn�T*��Q,�A��9�m-=lcz�|1�W�,��r
�J�9r�U��/� �Xl�ke����*K!b�cQp��M�0@3]���[VD4��֢�N��)�v�ٞ�4B��x2�
 �b�\�ĳ\�Cv��mM��Å�r-�C(&�=U�>�6��׵lx�4a�]2p'� w��=�~�U%%T>��-%_��^wmw�FܡcQ�������}�Q$w�x��9>m�Y^S`+*V�Z�ł� ~�A�J���H�OQ�[4��n��g��	�`�F��yK��f���̧��A��7h,����7D�ƕ����^���M�=�����Ǧ)��45r��8=�ZF��^�C8��u&K_�n��-��rG�W��P����oXRYk�&k�vrP�U���g�/�){�5�s<M��T+��֘��^�X����!V��M���R83�Ug"D#.�L���V�է����1x7�|�ز��_�Q/��9�!ڃO`�&��y�ɵ/����Ne=� ��I{_��{o�r�4�A.S3�e�o��Īln�8nBd���3��O���BU P�_����c���,�����W��+nԿ]���Ԣϱ��u��V)�m�5�u�Q�O�H1�Z:��G8 �{�J��N* �Au�_��#@s -x�����+�}�V,úտlr��ܬ/6������vN��`(�
d����3�x)�#~qټ���t�ݹ¦ u�Rg�$iu���PXcm0�r3]�K�0|����]���.Ү��qXU�I2�M3�{��ȇ�D�B3;^|�"����xvŁ���\��7#����#�# �s4>�n��������+G=��#%��T5zE�L���Oc�}���կ~�+���M��󒹖y<u�.:��@��b"����/oʇRA��|�`��Y�X����K�h�/~n�ek�/�8�^z�/>ॆ��rޓ��+�D����'���[/�Ģ�]��?J�E��@*7���YBx���ރP�I�:#�8���G��HZjc��-׭#r��r�e�9��G��3�!K�l�A4&�~��(#���|��韕Wn��3j�v*;1�k����H�n�.�t�2A��r5&c�,�9�ȼ��Ti�v�9�%���G���䘓{w����]�8��5Y��%:�W]�]nɉ�a*���2V�3����j��X$�K|䜚p8f��zܹ��4��Rؽ�!��Jv�_�Y��}�D�?{��K��w�C&�U!��#��5��!�v�}ef�f�|�5mc�F�>��j�~X)�E��l#���ۊТӘ�:?7��͔��E����d��ZD�:��j��f�U���T����xr��ܟ���98��L=�Z�#�v��W:z�M].F|�@e
a������z0�GzH���$���$ju���*	Gb��N�,����"4`�)V� ��fH����������Lc]�X�8wy�+���3V������/��1dݵ��P	rl��r8Y�kˁ��ۆϓC����Y���s)�$kw�~�e�ݷ�w�s�fm�~��.J]Y�\�oZk�Dv�'��RRR?�]�q�.<)��[V����Zzy��7oՔ�/[�P$�w``Y�����mÁ����[4���S������dr��c�D{�

��D�A�1Oi�Ѻ���h�(�2F�>����gh���0����J���e�a��M���"����xn%�+�J�?��H���K%\�OƓv��&�׀��2�|_p�
*.�if.s�x�O#�ɦ�6�ub�ӑ���\������-�G͗G����3���A����^;�#E�����NW�8�x�sxd�V�E�}K�&8���X�|��.�ɮ�lh�Ԝoe��MXB��no�wr��H%$���C�	��Q<�o��'���"u��-����;�j��gPWB-�ݿ	�FdrG����K�;����Qi� ��Ѕ}��'z��@�+Ѻ��M��,V�fQ��ͯ Ɓ43s� F�$�����,[Q?��ܛh|@�m/Vl��x1����{�P+�?�te�:z���;�	���&y1^4`�î���[۳�/��:x��#N�N��'(Y�B��n=lJ���7Х:$�aP< G���Q\ˬK���`�:��:�֟o���uQϋ���>�lY!�Ma��X[����}t��:�f��^�`S�L�|v�z��#�:zM�g��t��5��2*K-�'?�.>�n��%C�T!F�J�H�������"/J�*}èS����D��������Cu�4�&���� J��'����l�\.]�����?0��y���^���qſ0�Ê.�U�X�����;��h��O��U��:jrX�rc�����7ߙ����O�X����&��%�j3�Z/�-6�{�]'EGS5w���*7��k��;[��c��JQ�:Vʇ�>���HPϏ�8�1f�R��?��{�/�8cc=�C2k����Y�s��Of݇3��ٚ/b�y�!2�Mp��PԐYӖ����~���])���6Z���C�G��Ѐ��hnY<7�?������o?�u��n�Vf��ԥ:���.Tdm�iIC��5 ��np��Xr�#�Y?�3�yx���a���kk�fyC� ��K�(Ć�s�_5�S�Å�����Fx�9��HQ�V��)��.���Vj�~[�B�JE)~Ƭ�/0��p��Y澃j��C���s�S/F��I�y����|���-�}��j��G��5E�R�.�|ߩ�,��4�xm�TƑ������:#���te�XB�K0��b~���&���-Ouro����
R��F�VB^�L�iW�Y��`��S-9?6c3TrsK���� �)��q̟֎�}y���!�oAXwH��f�s�ȋ�X<|���TBeLc81���.&��~��z<�]�$"�e�:��v�@�Y��V�;�jA��\�.����&\I8��ps��Xzb��\��+��#��7�]A8�CW��)��k�3�������q�H�B�D�:��ƙϛU���!L��i�A��2�C>S�2�vYL�����'3���Y]�Vа�0��fA
'߳�5����A�´�h�4�SpɝS(g�!��l|.��4�����Ք!e��?���`��SR�:O볇�I�xS��XirG���8�vf���}�"Y��b04�S���[ܡ��lR�y$��Ѕk�9_3��8&S�V��Y�q��H����!_y�V��~�S�S��]TX��P��l����X�N�@���y)�����@���;�9e�q t[R|�O1�o�2C|�g����4C~�+�0����k�ù�� �U����� ?�u��ff�:�O�%`���
!�C�!�L�Pb9GՇmȌujΘn�,�L��I��|Ϳ�B��.��lEC��m
��� v�Y����5>'��&�L����o
�U��
��A���up��c���z��5,�犼A[@��b�2Xti�e�v��N2�QiN�;�dF�O�&h�xZ��s6���D�y�p�������S=M;p���_�\t3���Vt]zlxB�6ss���l���}p���#�>8Ǉ��jv�8ņy�P��%(3A'hho��*��s{�Dw�sl.�1֜Dh$tv�)>�C�ݼ��-˞�w���O�ݿ�CIR����,~���c��(�,��S�"�84�W\��{�~ӱ�������!v��]���IC�6�	)�����Ҡ����q��Zi�|i�J�UrHTM�D\��e`i@&aM�8�����I��U"�@��k��ޥH��uӧ1��s���2��!:�Zu~ݳT]1�˹�w|!�H�I���%�M���c��(�ۄ͝(,�_���|��Г��;�����68~�H�n#�H���i�b����b"�����cwD[3Y�yo�|-��{&m�P�p5��j�u;P��:T0��	w��z�iƇA�3����R�Կ���Up6v��pe��=����Vp켜 -��;0�txi�p�_:�QZר�"�&�`�B��i	��3���f�������I9A�XMy���01~��n;�?�6����~Nq7s�#IhD8��ulXZ��!"Ņ����fnu���|� �A. i��(շ�44Z�{�����gGҮ��Z�`RC}�\O,����MxeX��,Ovc����ħ)C���c"���P��	��L��"����j��I2�Ǳ�~����ES�����F}�*%H��ĵ�=�2��wmg=�[.�B�[�N��-��$�Yn��x[����c�<)�n�)Z�c���p�{�>���CC.P��%<yZ��H��|�"���r���(q��>���R��Zڟ.Ƞ�S�{��e)�r�2��?J�F5"T�X\�!~�±��g0�������t�X��녈�RXإ���C~\�Z��xa�
��ďX��J#>�v�� H����U]�c���Lf�لuS^�O�B��j��f�k���C�Ў��ka�(�nyv�\+X�(��۝+�q�<��s�V����aW������I@(2�ˊƘ�����f�O���l�>&����UUL��;��N���]�:VP韵5~|�=����u9��(�f�*����z��(������x�fh�y�Q���J�z�a72���\W9���7du����%�F��,�>UqP�v��sD}�����V���G~�[�9��c��{Jʈ?��97t.U���7C�l�s��=2
��-$�oi��=����/M>v���,gz�J6C��R,��(r.a��mKߍ{���;�i!�t덪�����dV��#>���x��b��:n������Y��϶�{V��>��ŔQ�<,�
��9#^$��q��/��ĉُ�;��3>O���	_�a��IM+NI�Ɏ�eM���+��?�}��Rgݜ���0�0�@�O}L�J7�v��s�x�(O���i���E�c�Q>�D`�E��R���p����س�����m���D����\��mvo�]iv�."ܣ��+,b��ʎ"&���,ro��m��8�G���႙�q��E[��@�Y�J��0� ���e����'U+ċ�G=��3KT����AYY@af�F �������0�r��oČ���^��9o���9��v?E�þlS��z� ����]�~�����~6#d�� E˕n,Y��y�����?C��C�Wvw�"�krKTQJclY�e����i�#�O�t�0�"k�av��UA�
z.��z�z����n�p��m,c'��%��.�&B���5/��&H_���n�BT��n}��p�[3T�<��Q�j̩wC�4T���#x��Q'5�.�,"��>R��ܴ�t=:���,�����A�{�CR�@���鄰C��B��:��V3y��(�Vd4��3�x�#�cX���Eh�Z� ����fԹg���H�Y����IqS0��U��A��p�}��{R��z)��������
 �]YD��hk�IM�TO:�Q�(�y_yv�c�Z���Y)�H� ���F4&`XԺ���/6@3Z�VQ���Jun�*S��C%H�6+_��?��X�Xbɇ��]�a���U#�FWҎ�����w͍�&[`x�ۿl���E��e9CUG���(r&�)I�
��REjZ{�c#��C�����!#�W����]}}>W!@�>uO=�%�=��?�ӓG���g���)�i4\(����v%�^P��K��#F-N���.��r�`pJ�����NԲ���"=P�����k���������`�b���Gt3=��,��D�v���
U?�� �*�9&b�l\sx�(���,�:IS�)�k��zNi_�?I ��\�<x�V�w���7n�%pI�(�)�ΕF�}�>�`?h���Zx`M���0������/0Q�K��u�K�vŚ'�T�eB�����:N�_�~T0ҤV�S��vH4V�;�ix��}*E(����H���/��P���8�)��2Kg�[�T��4&|���p<��Q��"e�8gEdi7g*e�-[�gqnE���>C��-�{�lΒP��?K~\&5���V�r� ����	-��"�s������,MYyqz��c왥�d�%M2�� �{����%���(w���3UWy(�Y���v�20��z�ǃ�¼ݱ����UF����5��g3�cS[$gi��н>���~�mf�iMB��p��x���mq3A�w�Z���U�H`�jx&߰��<�+����"���B�:?@7��&p���Q:RD�O�<?3$��?�lړ����R���|�+w�eV�|��#��q�lՔ���� �,K5�ɟ�bIa	���F�?�P�Gr�M1wj�$�c���UI���Q��C�p]1Ɛ�)�̰�z�ܫ@��Ay�uk̑]��v��PG�N2�F�̿���9Pp>���	`�8���lW@0>�'��UW�VA''����n	���~�`jS$t9���9`eo+�<���{c�k����V�@��k?�w[ċ1�1}{�����◊��� J���=�sQl�r�l�Zo�4*R⤧I���Mo۶�]�?��X{ocJ�;\��r�{�M�	15iHFtS�[�� 	
��ҺF!�:�����m�[,rK ��e�:�3_izxӬ��B��$<>�z6���F�+^h�K� �VNi�|r6�
]T���xdm��5/2��o��.@�#<
Z�VMs��.bh��G��.i�c���,Ut�񠷱�x7i<o��}��t�U�T7^:�&%�Ў��������~��|�j9V���L)
�h��ϑZŞ}�A�0]���|i4P��i�}ڟ��
:��v��Yr� a�G%���l_н��bӊ���(�Gg�7����[Tvr�n<+��o�9�d��&������]�r� r�˽�jt�q�l��H��D���L���f�U�F��_Na���%�gb56�A�YW��2r-���dP�iؤ�e�� ť�X;��A�h(+�C<�c���K��)}�:�h
W����0�:u��ֶJt�C;S�r�y���a|�3�u8�o:���]�6M��鳹�����	*D��m
����Ǡ��jؓ��V�˧���^���!kj
�k�����T*f��f�L��	�B}�n�-�6�5I�á�	������C�7w��^&6��� l+�z�����,��Vʬ���W�#�����
�D�6�z�T3�9��OҁN�
�g��=}k�w��w��׬�S�,3M���.�O���V\Y���Ew'l�st�B�Z����&e�$�rw�G�����R���g��i߱���.x�-B����R'Y����,z�@�>��/���e*ki|��cG	��(�C!0 �� w�:z�yr�H5��l�Q]��;�5�����?�'�d%�d��1� <��+����
]��0�G���	p�;�m��&�d̍&� ��L��I�fq~i�Ga*d��	�KV�΢��HX~ v��]�-)#`�c��O�À�xcO�]Q�O~biL��Qw����
Z�Ge��T����`%Y,,-
#�J���@��>>-����m��x> ����_�?�-�4�M��*m8a�챋��h�n&��b�S�ʬ��T�>�<�x{[��+U�)+SckG�I�N@�SWXK�!�*PiYdw�Jn<u��še����盓C�����R��Zu��$Q�J�9��e��e4��A�N7��L���'��VP(�,y؝g�i��f!��o�l*H����(�	�z1�²Bŝ�JKeF/��m&�Rc�E�5��'��d	��佖�R�U����q
m��S7ì��z�O��B#�# 4֖���`�{KA!��1q�n�|G��-N�&��/}d>g㾏g���N1�����e�ǠIɆdN � �]�֥� ���m�V��XF.V"J�ӻI|��>��0E[�8�+�>�s�q��o��E9my(消x�9��S����@0���8��Np�������q�ǉN�J�NQן&0#/�}_q<a�bv�mEC�(�=����4Bj�"�N�FT!�=��d�WZ�z;ܜ���52	��g�p#�4&C<�^5�\�f���W���u#f�N�A��Z�d	��bf+@�ͷ��Ҟ |�CC	�Z��WD'���o͌��@uZ�hzΘ�袟Ƃ�?�9��5�Ұ$����:�*O��1�G�Ô�&�?�֍��N��*��=�8��v{S c�>���i�)�9��p�]�")�<��G]�z��L�`*q<of&�aG�=]��e�L��.������q5J��%]U�F$\X�'�H��D D�y�*���8�E�k���J�P����r�.x.�Y2�,ў��k�Z�%�N�E�-,��Ѹ뜍�~K�cN"Q*��C��c8D����4�^s1��F�Z��$�ݺ�Y�]��D���+�h(0\�d�s�}bHO}���yl���E��I-jsG���T����WA/�n#G};�*�V�s5�ǹ�s������.���>E���M�hE�.uH���������\!3 D{��s8x���i9�Q�������6��)��S4�:����/��bR�Z�adH�<l���cϗK[.���ͺ�{c���Z�7����PY���F��V�t���)d��G��ZcČ���s#ΰ���:FW˯B� b6o>�ndm�#Q�}p��4.޼h覼���%�b��iZ{^������x����p^Z���B��6V�n)WT���H
*��ח�U]l�J`:DX
p���D�?��p��g'@s�֣�Jc��;��@�X��#���j]��cv�6}�7u�a�	�q���>��%		� ��f�?qd-��J�#ȳ�w %���{���.�]f�ܲ�6N�@�xR���L�����Dw���~2���'NY�P����@���m�C�џ��7�Y]��j����[���<qj�[���l�?�waD^\?lA��`���3��eP�cC.V����d��er�p���-��~h��:�NZ��=�	S9!N�F�d��%�ণ�w>B���r}���#����Ϭ���~����l��\��<-|����N�%~�rCW�za̟�/5�����>�&*c����ݦ�����b��ԁ*�Zy}�҇����kh�rN�1c5(ϳ��_��$�+�qpi�s����й̤��=�0��yxo�z���5 ��ݨ�r&���$hZ�9������h�
������nh]��I0@��4T��sq��y�hd�eYf;D��ne����רȃW��zW���L��|^|?[��k{\�v��c�X���⹙e���"υ �#��\xH�Ԗ�a�,�ΖT�e�s)8,��jq�2A�AgWѥ_J�� �od�#�eW�;��j�$Zs���_6@X&��sԧ�S$�lm��Jv�%���:��29T�ԑ=�;aND�3U�ZA�����@�d��G)��hBJ�b�>�x�0�0M��c�i����/d5�3�]U�QR
A����MUh���K0 ���Y�X�jgn��t�������K D�-iGid8�elq��?13��Xm���Sd\�g�@2��ͱ�|�J��q����4?�,�D�T"7�X��Y+�H��$U��@Ʌ�
#��p��>o��.AHo-�Di'H��Z��._���m�^ "i�4�����ΜGаͺa2��2CG�Q7}5*���C�Fn�zS�m=�|�	\ը�C'��i򖺌����z���lX�o%^����^�8�u.���kE�7	�(jLD�>���sQ5-=�Hk{/�P�z\:sC�0Q�]Q}e�I�Ge@��IzF���?�>��9�[�>'D7ܳ�u[�J"�[z��ߦ˔��e���(��
bX�o�m8_��}��ȅ��h�*��:�/`/�!ڂ��"��x��p�ԏiv������{��qfO�2]�hA�QYԣC�^)��v�<�~�L� �%��U0����' �Nxǲ!��66B;�'��S����	�C��!��f��ǲ8���׳ ��5�6��>�n|Ĵ�J�7_B���Jm/��@���i�xR�z)/1����J�$����o�k`"�(�R[3*b�0�� i�{��I��I#-l�i�U�`]M�q6� 㛌���1W4����|�9�!k�*���FD�yFZh��!�e���t�s�O�{��]8�t��ǧ�r��k�E~����e]L�7u<�����Wpjlcf��d?XB����8􋄆�y��LY����93�"�|�̱q]��]d�"�����<��k���YϜI�	~A9��l�s�z�)z�Բo\��L����w�?�DL���^a'��[���L�S-5'+z��x��jc� �عF�8n`A��T�n��0QO8������rK�)�'�������c��/�q_m|N������*�Աy�@�E໋��K� 'A����
�������u��;�����ۼ�|�?�kUЩ��l�YKe���3��@�I{�ԧ���{e�E����*�.HB�Z?�����e' c C� 2q�U�x?����7OG�$�O��.Nוx�zՖ�E�M���Y��� -y+�8���� ]$��w�p)�A�5��|��hT<�^koϜ`���wR^���oW*_�2]h�(Λ�`GPn�$�<̹��0Q�cU�f!}%��>��/Xw�_�1���S!�j������juH�PL�� ���x�J��kަZ�n�&�-����A�Y�5�ǁ)� ����beqӐM1_r�oL��HX;]z���xy�a3�`6�>tG�f)\v���o&�/�	�3O%����6��R��y�Z����6��Q+'���P��1���͝���C��]�b�w�#�3�[&7g�c#U� �vZ�.�{�ir�i[��2��c����ؗ��l��	���C��G�U{7�16�s��ΰ��A0xykp����T����D��@�Z�?�Ǝ�nf����iF��B��8�����zS��("�V���I�&�]Tږ�	�'%�CE����-����-�p��Ӹz���� 6w��1/�va�~��#w��7�-J����{�e�L� �fs��W�t�Q�� ��ѭ�ly=8�]�:�I��a�N�W�4������sdJ���{�D�I��1�r�O�q�WAGȔ3_���%]�������1�lg�
	��)���E���1Jp����R��5"(����x�>��$�+�&��Ȩ�7�"�W��=�rUM�d�V�����":�B�\�1�l��ͬ`1���s���^��H]��{�.�����\>�`F�%฽�VР����
�~N��Bn�T��ث%#��N�m�cTX��X��Y�QvF�V����`���G���^R�����T�"N�y<�θb�ݺ�p�(ojW̗?8����[�q�a��5sV��B�����;փg������[=�J�SМ�o�j�99\.u ��ߞ�O5R��şan����X��2�Ns�7/je|��v�)D{��t���a��ڛ]�O3��Oc,�B��͑�J����A�V"<ш�1C\RA�B�O��S�}/\���]��q�Зy`A�-�F+$�§3jC��!+��.LV�?�����gN�gk����������3�mp��*�b���5?�%"U��)����к[�g�y�R֥6��A���;P�R�d�X;U�ay�tud�b�iq	b�FC��U!<��bC
����=��V�����3.uMgBվң�����td��!G9pc��Ī9߅/|ObLk4~��7�y~t��L�h�/U�b�u�$:�q����4��y�Ǽ�e��,��)�P�(�?�4>x��Q`~A���Z�S8q�{s������"�YT��ֳˢ��� ��%��.zJɼH�m|<�o�k�eh��h䱊��I"��&ŖִB>�PV��,g��ka��ւ*�xĊ���0~F��ޯ����;A���[��]G� �Q�,:
��tJe�����y�r�������o���B83Iw�!t߮П\�	���t��\i�q.���3���05�
���ː�螽��TaJ�Z`Z�§��l��uEK���s�H���7��z�$>P��8�4 �\�A�i[��k�{� �U!ԍq�˞4Fn#"5������9�!PB�ݙ�j��A�'v_�Bl
��w�g���;��0���\�)R;ð�'��m��H1ˈ��q�"Wl�iH���Y
5�[�m	T0��º�.�p"��A[�����@�u�P0�5�yg�������ּ����9�2��Ve遈�
+��EՃ��_�-��'�_8ʾ>��L �ZY!?���9-�6���"1ڇ*j�Г1�h�$����z;�̔7��U� c|�)ip�1/��(��Rխ�!YH��i��1;�Y?�o�3�<�BY~��Lk�f<�/�_�+�X]����5�Kc<P�b'�CJ�N��e�W�H�֘$^��A����@%�������H�Uv�~�����/=ha�F���^�]IO�eEa�Kym8e�O��H=.B\�xq����ƠYٴs�̵��.֜��"Ϝ��6�Փ$����O�+���$m%�D�]���܏�R���7:�=a��Ƞ�"��į�,���A]'����X���w݊��q�b# 7���OE�*�0��/��"더e��0����K��{q�Ũ�CQ�������U_���H��$�f���q��_ЦVn[�ͬ�O ʺDܵ�P��j !����ݱ~^�K^��V@LWY5��I҅3 u�|�[��h*�=�hC���HrhG�hTDMt��5���v]r��i��zl��nfQe���DQ�姑��I Y���h��}�ؾ�=��hTWJ��䓋u
Ie����y*���f7�5�����B/H��Z��&�e�����5�J��)&�k�gO}�@<�їa"P�ד~���X���5mH�PP.���8�y����g/D��g'�� 9�9�`E��%�,ޗ?\��fz����Ue���z�c�`�}�4��u�t_T>m��FU�s1$��IK�"���P@�����7%�4n�����c�g�;�d���ch�mZн��u�XA�]~�(v�":M���3����/H{7p�BW<�be�?#gV�t^��oQ?��I&ԬEs�8��U�xToy��xk�ॣcp�f����8�
_�n��Ԟ�c�x�Fy�%ï����a�֠���݃Z(���s2���C�Ɋ�5M ���sV_���>$s��a�X���Q�i������j�
@�ݛ��gz����֏/-�I<O����C��5�3�H%�AgTk�� s7��&# �ї,�;�N��R��U�<ۗ�ߓ�$:���?�890�7Ӵ��?k�RpU�/?1@����#��c�*
�j��e4����� S�	g�'�^�J�+�<�ֺU$2m�ÿ�9��@E<%ڢ��e��\V/>�3���uzR�;V�v���D���E!��J����E�W��Ă.#n�m�E��� ��p=��2?�78S0g��6��i��}����{8���B������+j̶�WO$^�!�{c;`�|�ڔ4�21$���2�n�w��jf�@�Y���f8]��!�DN'��5�<�AR*�c��<��|��r�]zQ���󘶗�+�x�!��L��`�-cX��롕o]�v�5"eF�������N�D�.dǡ:�F�ܥwzQ?:�J��pX�mwVE�>���Ѧ��Y��$}�.�Q�ԼI�i荤a�'=���b���Kô�j�2c�����x�������6fh�#|t�ﬞ�I�d��m(�����&ŷ�|Qr�k�Չ*�%�Ha�ۢ���N/}J��5�v_4�]�
5�82�`���5@�~L�Vz�[L�*�%f��o�K.�s���!���ֻ�q�
ϴ�y�<Eu��xO�Lq(} �A�k��/��VA*����P叇�{��,��k����aj��5M�Ae�Nd�y-�ȭ�ε��)����rgY��+�ػ�X���\/n��%�U�eϲ1}�E���?ݏ�
H���f~w\�,9�}���qk�����Ŗm�x��_��<��dl�^�k�cи�09��^W� �._5��-԰w�#���G0Gy��]&�g�pk#��a�����|g����>c����i�y@o9��VER��tR��O7B�c�?+,�$��A��σ���,�Y����?*<|2[(?$>�+!�z�E�6P�Ւ��ĳIU|��0~�c�u�觎P"�2��_�hs!f3�Td6����v�J�==-R�I���L��D��іӌ�r��`�CWn���4�T��zK)�k�<����m,51KJ'�yrRE��<۵�����k��-��9\�6+z�$"�.��Yh��Y���s�OO�j=o_MO�㖾��+
%�6ֆ�m�_��TA1dU_,��Y;Q�5�_��E|Nvbl[!��L�q�� '7��!�4�z�ǚ�)��]��ׇ ��A+����Θ�3�/��,��+�ڴ�3��P�+o�p��)�-�D4������㓮`qh�EӉ,-t�� ��V�jư��e�9V��Dҩri�W�mᮆsήE)������������k�ݘU�F:��o���������+���9���Lx
]k!!L�Q�C�������V;��D�Ћ�r��%B��*�3,�oq� ����F���*qn@�\��m���������	S�{�p��(,���瓌�����{�S�c�\�G�ӡ���6�&�O�1�����˗Ʌ���q�\��X"%9 |����"uד�C�;w@���|�W�d@�ܝ6Ŧ�!h�4���z��A(qE3�k��Ե��Eb�7�1�� �-�~3�]�Jq7��F��$��"eglK�|�Y�$(�A:���!P�a��$�I�t&i��r/>P'�������0���+p�D8tj�- �\b1���"�]|��~��]��ʤ�5i4�on�i$�3�,�}ǒ���͆6P�+�@�&\���'t�8���{�gHg]\�<�xu�ͤ���s�[kT�i��K�V�1���cߡl$���:�Wi�2¢�%�Di\��q5S�B��&N��oS'�k��9���[�<���׶�Y<�B�@g��}kC!ݧ���#�Ԍ)���uZZ��r��(�}�VR�~�~SIL.�"6hO#�)&;�%cG&�1o�I�d�4X��d��@�gл�>�T-�_��=5�c%�K��v���+���(Z�,�Y�%?%�]aKe����q���½���������S-�g�u�Zg��F`�Om�<F�~&�g�W�4�rںN�"8J�D�F#h-jr�����N�.�^��<��V�4����˙3�_��f.e�S�"x���%�z΀��7�\��ZG�?���$Aǈ�8k%��7�c@ߌ��3$�{��d��P�M,l�B
��7�z��a�m9>>ݠ�љ��i��4�X�9�w�
�x��̝C�jW��v�F�c�b�h1/��8{H5���H�/DװS$�\1��'�a
8l�g��R�������a���~q�Bغ�����_��nؔz6#(���	�)r�{��J�p�O.�M�C	g+�.=�1\
m�C�)�z��cf�U�<����3�u&�k��{҂5ϟ��9ؖ�����Ca�O�o$����&*��~�J�wq��S4)���j��������\�FOuDwv���j�t>lq�����x������: �sR�ts7�)�~ 8y�*I��>�����M�Օ者aO�O:�k%�q*���Z��M:�y�E�ѯp��k*
���S�r�d ���fb��Ke����ֱ��qQ���]��t�{=��T���g��A��^&���XH��z�{�ɩ��.�;���k.BY�_���}���7ّ�h4в��#k�����}�j�H~Z��-�����`�Z�~�6�#]�A��]����/�����Q�MDb�	�$#��d&�P,�8P���R���v�H�˜N�<�� �%k
�>f��q�W>�cI�rg!�Q�S�t%J=<��yGŠ�}��_�BdDC@��{eet1����cfM���*�n>�>��/�}�?�����;��{�	���
wAnN�d�m�-����<٫�զ�u��*R]$�_�4}$��
���:
�㊢WE�G�GjJE�gkp��ҨXx��g"��d���=�FeDk�y⷇С�W�f�].Ö4w��[<�N܂�:"ha��*�6�lL3wf1����"�#��!�f�~�f�z��Vc��S ��W{1�8IW� $˘�t^{y����*�Wr�a�'������+�>hS����D����܆
;IrVڶ��{�X�K�W��<�t.q3԰�����"7ZT3�y@E�"�k5�r��$��r�?���f�C%�y6�PSi�1Q�'UeX\�oQ���?�z�Cuz+��H؆Dz�%Lt�%9�� 	%�5_M�ַ#�����_����Ɲ�1V��]h�t&�QH�v��_���l:�"N^̜��Q%7s�`��5N8?�-�'�
p�"`:2� ��I^�D�/崃���%B��*8$�`�!�?66�2	h��nn�t�vƞV�m��ܕ\�c��1[	HD��������xv�TVбk�&(j8|r��bc�������o�\�+u�z���`�*��l3r�Ú���TB�^�k���y�7�d�m&0�Q}����Q�Ƃr�%S޺�D
��gN���G`t�d��`�S ]��b���l���!0�,a>G�)�q�d 9Qv�!eXՃ�S6�?1����ZT�Y{�2S�^qZ'bF���7�#�v$��S8�Fia�ɔD�Ég���D��-qu��4��*��Tcᇞ��$����$��<S"���M����~"����[V�Fa3W)��W��M����c�u�N����5�
p�i>$ĥ�ѓ�"� T1����Rb��[So��8�1jǑ���׼H����t[�y�� rUo��ع������d�m5g,1�ӵ_!	����r?�T����+0D��t����.�w�H����-����!=V�r���o�d���������7���xe7�U;��5���
a�CȖ�����4,7m��F+\(����x6��&�e���C�#�f�=�rQ�P�cs ��6���ӡ?q��Vi<EFDRZ��n�F���ǖ���vI��+L��F�2ߘ�q�#j�������Trb Yqt�C�?_MV�o�p��Ag�jcI~vQe��T
cBwE�ay�/n�ZE��S������?�;.˒�7���o��r��cX�ՙنߔ�u���0C�j����YJ���$>,�;i���i��D��G,�ZBVÑ�Y�0�.�<"���6"�w%�«%��W��_ek$]�GX��*%�Dx��7��G���H��I{�c�I�%n|t������t&K�����5N�g�K�`�f�;M�?H����I{��O���@����|9;ց�7�8��gr��p����m]
�D��};�M��΄�삅�;���u[b��?���D�mƃn�Sڋ�0]c�8����8Ϲ��V��d.Z�Ҩ��TF1n���.�+Cw�9��.P�z�wOZZ����w��{V� �I�R�������n6����BJe���CDyC��)�ݬrs��r���>�QH*Q��<�Ā���4���o;U��6 �q�i�<�G��x�\����Xz�����m@���ĵ�	���L�ca_�	�?�Bm��q�{��������*�/XӢUS�v�β|����#ps���;�O
��!.@N�4Z��BUb�����<ꃉGZD�P����v	��m!
@�׎)�舋�xSU*"~l� >v�i�~3K5�l̄4d�8c��x��0O�0�1P��d�y���=K��wU��k7�Z����j�?���H���Γgґ�����L_V�Zf���O� ���_)�5��(	����9��?8��E����Tl�X	���HH���͵\k�������+�2�TX��S��i�X�0x�_5�sJ-J�as�uu變WG�|
,{�o�>Tdz��&g�C�5+Wo��"�^��t�$V�o��z���s�e{�[E�Y3�<7�8Y��s��)ވܐhu{��`�P��?����]WaI���&�_+�������X�{�u����h�"�� ]�*�QB�p�8rm�6�w��=GK�e҉Wjo"�X�p����5��ZRt�y����ןMK]��K���2�	�B�Nl�jX�J���0���-T� ~��"�>z��,�,�:�ݑC�y<�݃X�v-l Fj�H��ĩy˷�mʃ�i���w�B2��@@�f���u.��e�4����Q��'h(�u(zY�O��q]��̎��Ic�-�ԑa���8�@����4�r�4ǳ�E��^�?擫sr�zm'�)�ٚ������� 
\���G<ƓW���e^V2 �~]]ԯ��l����Nζ["|��H5l��A���#����B������4*�Co@�M�u�$|jذ��>%�A�|�xC����H�,�LaXv�(ɹ <�V�U��\;����D3�v�Q�~����Z.{e5��|�ڼ1�ض�Z��������9�C)��)l0&:ѳ�Ԉד�L.����!��Ⱥ�wAߑ����4�Uo�+�^o?
!$4Kսو�mtwZ��k����sGܧ]4�3q� IO|����GJ�4u��ã�9b�Ĝ��8����P�??�{JluN����|������>��� �Z�m,%{�?�z�o�h$e�����9u��W17�y\H��:Lӗa�UWjjޚ��P�ĶH����V3_�)[?���&VB
_�E)�����E;f����}V�6��t�;��e�sp�h��Te��4e
uH�~C�R>���i��q]nJ®��X���s]���~é�3X�h�������mޙ�������'��O���6�`�sd��2�w��߿d��+�����I���l����G��ao�b��N3����ι���!������i�%�:8�j��Ѧ��� .�瀭VC-Aa�����K��3D"H=ɞ��TYM����,��R����,���m��j����Z�d�r����(���
��'���k*�L�͙����Ky�t��0��L"e_x��A�<Δ~߈��� J�5���կo�a���d?x%�zbо��\�k��V�� '��uH�0m簅d�2�m��]��L��d$�x<�
g�l�ʬ�n��/�^Ͼ�'W$r�>h��ia�w��2<��	���0�L��8G��Ύ
�������z���J:Q}<8X\�n�rb�Y{A�s�j�l�^G�����d�8y8�}�J]��4�v�p+R�㤕Jjwjjv�"#�d��zmQ-zB�K�wO����O=�b4��W�D3�lhǮ�] 5أ��D��%�W���⊡Ǟ/_h*���:b�߯���i�6�l�	s�F���d�v�p���>qJd����)w�rJa-Q|.���w��u�fyE驢����N�TH%o	��٩P��ZD(<�]���vK�x�D���J7n�u=�B�o&�$��m�����%��H��
VktC��d&bjR��wC�?���c�$D��@@��� Ȑ��_�f�����T9օa�s2��Q�*��m҂�~�%�N˖�����B��V�W0��O�"0O��sĐ�0�Y �f��؍~��q՞V[����1�Gm���a��jӹ�H��J&��BJ�YN-���b���p��R��W�y$���+c�7'E�be��쭭�H���&;>,P�c��4Ci����ǰ��gW2>G�;z�Ǹ�殺¯E�;I �����y��s�eA�����p����M�:�aGg�Љ�2�O����-�7�a�_g���V)��P܏�h0�g~s���Q�C���\�%��A�z.����G���Y%' ��ѽX4���K��[DGa��sg�4���9�d*Z��<��0�KQ ��뽞,��x���r��dH;G>�}�9r�s|ѕnUm�_�8qEV��"��[p!+�����hEF�)wGlL���&�(�,c*,��1��b j������Η�A���M������p+��'�������f��桯k���"\�I2M
���ӥ��l8=��gΜ��ٙ��1�<b�q��XX[��0���`����j�}���#'�c�/�i�y�j �g
&�(�`P�gl81�=�9@>���h�8�/�4��������(�'ìE?)��|���|�G~[	 v�k���>�/V2��t/)�����V(=FJ�4g󩈛���}��2�S	���)=gOh���_�O��J�.ӗ���*�`?�F�7�%���������u�����E �!)FQ��S������xbaGp���b$ƭ펙Ȱl���`����ͷa�����2���[r^����Ĵ���Xc���	�X+P7>�D�/Q=;a6����iB�!qA@_�O�&�94$@��zNG_���H&��O�'�_�rw7�=sCi�qC�A
>Ǵ�O�:g�'
�5��-���r�5�*��	��Ϡ[%���)w��\u�P,��;1r1�)�^|g��}�/7�oQC~��7h����[!-Z�O8� ���}y�n�=!���e�5ӛI�"��87D3KN�A��;��܁���A��D�n�fn����&����U{��"��t0���o���=�ك�ch�?�/�H)������+(o�k�_����k;h���W٬,`u�D���/��u�ݟ��6�U��Y��)=�+��kM���qk^Ma6*�ξFO��[5 �B���sLw�f�����X1`}��N�� ��b��f�+GL><�kO(%Z�;t�nވ	�Lg�բ���ߨk�*<�u���A ��A��3��8Z��fRC�n��iUJ�L(٤��(�5�'J����jy�KH;ބB�2�� )�L~�,aѾ=b>���e,+S�������j��Ü&L�_9��}'Q�/�>^n-������e)�&_�����ݮ��ί>���O�6�,����?�,b���_����A��p������y�.�[��ٵK
3�Wz�8�(Ǭ����{g�D<Z�I:x� [~����yr`����Oo�Zi�m�ՐC����0��$���D�5�(XB�h ���xn�����V]�}Shq  ��6���t0�Ω�(����V�%Lw�'��� �_ZWb�F�#��֏-�&�쯎E5���RP�H�"Q���#����E�a�"���ͯU�b��	�k1Ȕ~�`�U�p|�-/Qz=[�ؓ@U������̳�b�	L�kN�U��@i���i�<1�n}��-	�<��F�E���d�F�Cvp�*r)��\�!�x�>�Q�;^m���p^���d&�|++{QP�
�l<�<7���{ ��)�GD+��5o�mE(�2��e.����{3U�h�K'!��m�:���[�\���� X8NB���U�*�eh82���2	qB\��)Qd�ó�C�� �Zw�QV�a�y�y��:�=ܢ���%�_�����F�??�}�5���q���eı-T��1��Ͳ�>�&�u'�RQ.��r���G� ���P���4ĨS���m==��˃�ck�}���@�g����"�&�u
IYf�=u`~��^;���9fGE��}<�D��$tA�q�f�{qI&�>���x2�]�rK�|u��6ޯ}a���iuG�}�#��`�#^)�&}���4l��kDC�ܥPó�<�n}�o�6c\�k�Ȝ���]��go����� 3�bM�C��AzE��c�R���B��}|>=��� [��`�ZG}~<���n�m���ڀA�!!i�k<�b"��L�+�fk�)'G�`-6��X�&�e!�&[~�mzN�y�$�RE�!H�d�\0Rs&�,x�Mr�2��P��,'	����������QU�}*�f0{){��-�~�ӫԃ.9*mo�|1	T/�mQbȨ"{߼kT2$��{��b�7�?XQ���%#L��+K��m��!p��%ݘ L��Ǽt"<j:�S�f�������P*/��f�X��2uL�u��E�6K�L����>׽�𐕗���+��E�Al!]�==a1;[��F@f���]�Xq?欺V�t_�g��':D8���u'4�M�k�-����	
*9�	��\B������ڗ��k*d��{�j�%��7H�A���B[7�Э�3���'aqݚrG�%1u�]�^½�csԫDԨ�ɀ.�����f	BC��@=�NFd�ۤ^���ϥ̲�l�z�R��]�7�eg�ʦ�r�(�2`|u�s#f��SX�l6A}nO��A�(,Zc7�+ �#��h�P�I�/�2c�� )FI~9�=�0	Q|�2^� �CӹM�������du	fD�&P��>4F�ɂ*�8����=e�bp�K�'\�v�!��4��L�?��f7��H�=bk,��v��{~�2z`�-d�L����+�8& /�o:H1(d�O}��Ұ$���#,/����Q��d��x'��>�{X����"@���$��bR�-8����Gs<�^��J�1P�k�/�c쫋����j_;�����gU ��|��2�Ç��������X�8�FL��>����u8���D����a���_0�%%�A57'��0h��3a<9�>�,�m!����m!�T_�k���t�5��z��E,�3c+�����Nq�鹲�M�kڞFfF꜏�K��5x�?C��)V7O&��F�^!���dI���9�o(�ڍ�ʣ^Q�L�ӡ-c;)��p��'	�"�kN;��ʙo�3ވy���"�)*jg�r����@{�ܵ@�r9	�_o�Fɐ��L�m13t9��K�#��@]*:]l�7Uw��1	����.����N��f[9���O{5�E)�	�L�]|�}˱TX'}�$�v��2��}(fyW���2����o&Be
Z�W��.r�9�d�r�t j��8'��.	+�o�,S�;vF8�0�. ����
��o>��6{m�O��`�U�m���ܤ��~��i�D����rf���E&{����7�^v
������	/K;:{�� 4�f!�T���[;T�*)۹
�� ��W��5c�|F5rK�<�g )T���g�X�"N=u2��CX�
�I�o��|���9Zd��1�"���Deǰ�dkD���fѭ�`������#�.�mŖ�rx��?a���'�R�� E��	���o�wp̨�k\p>]��7C�'�%2Ψz�1��?�Z�Aw��G.��5&�HO�Cř	1��<5��Ցm0�z)���YmZ�k
wFb�҆4��r���*-X���ԙI, *%H3(��=� ��1�6��5I�Q�#�e��?���'N
;�B��d�P�n[��A��%����n�g$=T�{e˛�@��f`j*J�Ief��� �?h0!xT(0�D����M�{}"Sh[њc4�V��j���������S@6^� ϖ}�y��ӝ����l���p��H�՜���WL���&�v���溞��-
�L����:���3Eէ�}p>�no�.QmY�|.�L��j<�x�����?즫e����G��7x����������'��f��:�0���f���x�G��=Prc\G��"}�>o��,�tUW�`m֜����5!�[S���6:z�FmY6+�0�����dg^� ��0�'�c}:��������#��yH���$��d�]��������6���$���O'�A$#	�`J��Y0����S`���#s�M�����鏸V�?�_a��ݙ�b3}DGN
F�0�fwE��ʛ�|(�zV�J��?k��:�k�B[򴂰��j�t����o.L��i�8vN� }'k�Y�/ճ��>4���g�?㯨[�m�9�Cʬ�wI�P�,jB ܶ�`�Ƅ� ������7N���^��ß?f֑�ChE� 9�f�&����K��T�u2�&�F�LbZ;��@�}�ҿs�?Om-.s�i�BHR���f��|�z%�i��-���=��H�H�z9R=mt	~O�*�K��2oꁮ�M�'o�"�Ds��8r=�s9�^�\t	��m؋��)��P���f�S�L���P�L���Z%'���1�yF��ɴ��"9�@6��mq��V�����Ҥ�??����&�0��N�yd�j�ߋƱX��i
8!<J�bY�Z6�h��)m��3�)��bbB�-i�-��*K��	����I��͙ge@׊���_u��æ��1���E��� ꮘ��W���<����9�+�C��0�ÆY
G"LG�#�}�]��U#�$@��=kxVe��)%�a�|%���a���Ԙi���I��׃.n),�E~�x�9�:j>�n��8�������I�|@L"��������>\#��4��̩��-�-:��{��\�7d'�g�tV�nd�17Y:��Y�B�������h��ZW���7D�F�e�˓Xz����@�@�B��e]�o`
�\'o`A<�e�v�S��ͩ�0L����}.�ϗu̿����%��ME����>��x�bp%<���A��L<gx��륯�I�P#�ZZ?��#��}An�T<��w�؝~�k�[���w�ͺ�WH��ǬU�gV-ˤ�N���W�PLAɘ�x�P����
��A�d�e���P��݄M�&�0�ɬ0��L[�+&�F	���i���y�*������D�F<�9��|ݿL���+�圻�
@�Cԑ���ۗ��2���(�&~�f�+�	�HH��V8z���l;@x�6��xF��b�u�~�ɨ���z;���$�j��`���l�x)/+��pbȭ�(�$n�p��$ky.�?�B��#��m�S	B=�a�n�ڷ�q��m)&�_qg^�`oUݮ+�g���>($�T�ݾ`���]�n�/BZ��J����0�8d��e�Q]��B�G�K��(p��VA�q\���f���8�	�V7���3ȁ�g���NQS� �P�ʬ�&sq��'��#%#�9�����I���$.0|�@�G�m���+0*�l��tzz}4?͛ŊDS,��e������Z�a�	hf}©��GޘM���\_4��(�z;�Q��M�1�f{�]\+� ؏��Vt �B����P��Ĥ��\i�� p�DS1w���g�r8VE/���V�8���;��	S[��x��GBx��O��5�zg��U@Z�;A��Oq+��}�8�2,��L���N�Y�O��m����}ZMrpa�_��l������T�q��477���ٸ�8h���^��L���>����^Z����m
i!�1W2/�89:�[�b�;��;��Z,��s���� g�Q�B�Rm�r��h�d[>�)Ё����jfj��s	hc�R^L���Z��8�#'�ܐ��J�g*�-�k����MmZ�C����3߲&��J-$"ȹ3E�"��������!�JC�dKJ+N�	��K����\u>!;�u'�����i�U��>�C /��6Y�4.��_�t��u�sǘ���b��i!:�GXOy>�F�.ՃP� �|��Q�C�u��:y^�@
��'=~kO��E˥m�Œ��O�s7�^��=�+��<��M�"���o����M=�x���ˠM��Z�HB������C�����# �M9����9���'��U�m�V%�RK�HZ����U��g���@�C~E�����[;��fy3X�s<6|�g:��ۨ�#` ���41?���8\�۬:K��u.+I-�z�w����z���0��,rny:��=�^�ޫ�`H[OE��Q ��J~ș��޿�ͭ�	Kn$���؎%;;�z�ݱB�����[�3��4R,��]ɣ̏rF���<����P��]���s1���KݓO;�J�|k��lq�H�M��e��5$Õ��;H��F��r-�Wi�`�u�D�w[ĺ�r1������a���|�cc�l��!P����$�Q�8�g��ˊ�I|�����f�(%ؐ�S�@Q�����z)��r��L���}ß�mK;;+a�:�&��r+����x7=Į�&`c�9ʞ��6t�8�cd ���$dS:�9�k�������@�u�l�Y(�xz�Xf�Q_pM���S��>�TV\s�d����-��5��=x���dӀs�X:˻��2pY�Xy�m����]�������6�w�9T!�F��=�DK��Y�:�|�C\S�L,_���U�z��&�����r��gG͠���������5{��\��PO�0n$m˙Q���|Sz�_�Q�Y�t�s�,�����Aݼ,}�&':j��,��S���>���#��,��!z ܦ��"���M�#U��Kקb��/�Y�a��,5��<5 ���(�$���\L�[��5���c+r�(�(+|����y�Z��%�I���z'AC�v�iuҨ.o�P���i?��go
��W2�W0�i&תF�V� �Ϻ����A���s(ɛ66E&��Z�LӺ:�E�"P�&R����vK�`��B�X�Ǻ�U�e]9�dthn��u��	�S��va�AW��)��޻�"<jk��-�
 :�����.��+<��N��n��]��nY�¦�p��4�?=41L$Xެ3���R�Vv�Y')q�k�~�0����c�����5��J/Z%�ʏj�1���Qa:`����%Z2�u���Bx�_�͂�K��i�j#=៲ߒ��X��oW�{�[~����|_�I�b�3nm1�c�׊���-�]\3T���C�����S#�h1�A��$]�"l�+Łl�I��I����G��/ҎXa9�*&x_�r� g �KD14c'��/�b효9'�����>�G�K�v]É�н���(:�C8{�+�뎚j�0\��dje��k�Z��x�W��	X�� qHM��,q����|����D�����Qwɣu�+s��De�bっ)���?8���ՙϟ+ef�������[#V@jt�� g��,��:�3��;J;�2��<�a����2c�L�A�:cJ\zB4����Cm����*�7!+�ڥ�>m�D���!}'���FnoP�i�u
���jF�d�V$ULJX��%��DM����N��0� ��ר��i��&��8�\��,�2iN@�f'w�A]�������*M��!0Ӕ��H+d�u�ɚ���©�7�K`����[Gu��������ud�����ܵ�<5!�%�]SiF��%@w�-*p�I���}�򱧖��'��Ea�?�nBjJ�.B"*̫���1J�B��;x�%�:[���w���@�MLn�q��oÔآ�qo<��L��U��ƾ�]5�@/
�'mU.�u7��8!��-e��ݜ�������me��j�k�	#�W0K�1=�-��=�]S�&ר���(a��'�Dvz���`��,�r�2��ُ-���N�c�R'}"R8�M�l�̆�eҍ�n��q� Ng��f�8�c�c=�d��Ԙ�x���/!/Z�r߁4s�u��5��8��	��G	�ٱ�UW�G\�a�R)���N�eX`��>��%�P��7����Ц!k,��Z�7kKs^�x?�!�<0�$��w.[CP�^�3�����8�yܑ�*�D�g�=zi���r�m�%��������*�t7�9"K.5�.��Sû�x� ɎǇ�~���NAQ�M�� 0m:��f��:�*�\L����m���<�>P�Ц��n�KC�*���0U��W�Iq0:��[z,���"��	Z"j��nw�vY
N۰޸�&�/_���#d1@��B~� 8~_��i��w���,B���g? ���=84�z����#t�~���S=H �A��,!�����/�xեL�DS/�M߯�М̂Ч����n���C��q���5R� 5j��Ip%�S-d�y MO��_Ǿ��{�����/�����!EH}��*ꘪ�-u�����21Ȗ�i��jT�Qa/�#��^t�D}�ڤ6y[j��W��H�7��i�i���O�R,�4r !%��.��}�Y����-V38 L֌�j�tiFj�����P���+�[�<�9z��2/c"���zI�ˀdF��b����|�<���""@i���y֔.�Q=x��<vH�K�9o;㬩+"l��_3��rj�����t��!��X/�+�nAOC`y�&(�����<���U�JL)m�3�тS�߽�Q�\r�����ɿ��v?�l'��p�9{"�9��ae�rp��Zg���Tz��Њ��:B�j=ڝ'�*�M���8���9zB�N�!�8Sa��2���C >K-p4�
��TZ�O��?�fxg]" `�_�:��^K.�f����(��<�㎔� ���L��\^*%t���]N�]H��M{�q�\z˟{��o��u �v�ȸ���t���W	 ���������0r�h�6���S�q>GL�P�9��Rs������Y�uz%V(�&��h'h���zf�d}
�e�t�E6�R��2aP��>!J���1#�祮c �x�~��{�E7�}@��r�nؓcoSxc|���EDG50�Y�N�WΆҊ����j�B���.`�!�\��S��k��5���,r{�L�-*c~a��c���r����+�&K���!F��D�\��y�{��' 1H1��3� ����}|4�3�)�E�3cW�������}��ǋ������]�l��<�}|�K,�s�[{���e���:����.a�A����#u�Ћ��lD��'�H�X��;�X�Z/[���`�Pd��$�Ȕ���%H:=�o��@)6S��1�t�����/�Dvlq�p�D��G�p�A��}��7p���'A{jY.���5>�xT���f&X)8�̈���Eyb�YJ�'�h���-!�$8���vv��)7�%���{B@��ŏ�|�5���N��9���U).���1Π}*���\�ܤ�f��7R���@�jhjw(��J�n�Y97ˠ �sĢ�:��xH� ������Z�8�k�$�Gl�OZX �]���?yn���kq�5�R��ѿ��a���j�V9�f�� ?�L�.z߽� ?��/���@s����F�o���� s�Ҥټ �M�w|r�Z��W�q��..��,/hlb�O��?ySSr��)����>A)tG򖰂F�cؤ��q�o&.D(�=
�����_�I����h�ץ��.���?���T�c8�S�+�YП�[��X��W|eɢ�oy,��'�V�9��	.N*��C����џ����%[c����G�Ci`�[��;��a���v(ǙT���T�>r<2�;t*x0��F?��k�A.?ޛ���9~#�D"uI�I�8�����0�"sK�:'	b�ym0e���S�}�0:�.��2���"��ہq�T���몞���!\¦T8���,�[�-5���W�$�: q=>�u.B$�}I��[:N�5B�'�p�Co��d��Y��5*Q�ԩ2���(����#~���q��IM� �N;@��KKa�mq��B�����6�i7, ��
Oa�C�$RB��Z�S��!C_���9r�"O�ɪ��-�m%�!s�6.�h�[Z�����w��gD��s&IO��IxW���.���\~��?:���5�z���Y:�7�,����q;ULk9�3��/H�S4��m'�d,��I�aY�s���� T�6�Q��z��GL{%��l}�q'T��K$�;1^2@���[�Y]=q�Q�z�lX��r?�i��!�uq[M����{� ��kj	��l�oQ���J�����^���ht���}���:���.�wZc�Q=BC�i�&�,έl����6-��T�%D��~S�@�	*o�j�h��~'���*�'�]l��Dtŧ+{tpu���c�$���h:K�RH	��5�8SD8�$���k�U� ��3�l���B/J��k��C�z,�^�9}D���L�%�!ڜ땁 �Ͽ�ٖ~���7:���|��^�����kn��% ��~�9+ӌ�M�2#NS8�~Y�b�d�5>X�q����^,�jt�{�҃��>m��\F��#�T$��B�S���h����t<C	�=�%~����k����t�������B#L���^�y���KG��Ű��LE�� ��/��+��e�ѽ��GJ�Z"���@���q���7Ȑ��k{��y��i�nf��j���Ͻ)�u�g�����C|X�b������O��kŲ�a�&
@���L8go��9�I��\��U�nD�cJ���k�!���֯�S�s1k�g�o`�^Ȟr���`W���B*��v;((�-��{�l�+3k�<�o��چT�˕ni(0)\똁��s{AӦC��_{��=[�QSzW�k�#�r��4��K�Q�{-t�b���B#�w��Vo�M7)cR'��Y^�A9�<�w�*����e��rpO���D�T�)k&a�%lE�	���Hۑ6o|# ���E��m7�'%|���iW{� ����$���Y�ҥs��l~�j`Z���%z1�����V�Eީ�}S��E���s��3)5b*(���%��W�)Eڊ"���@7��#��~* 7�0r.�>G0��Z� ���$%1(���	�Y{��د����s8_� �y�g:���/gG]�ę#�I�x���DS�@�ӽ��oX�}n�K!����<�� I�4�uR�^����S($T��R� ���M�W#���J��wu��
�a�J��>*J��9�"\�"��'����41T�L��m�7de��q��^р<�c����ms�e�ͩ�p��Etû[��N"�i�{n��ye;=��^D9p8�F��h��z�{7»�>hD��|F�Re¤��ְp��#⛟@E��ma�L�g�آ_:��u�|��9k���s���S^=�P�7�G&1� �,��x#f��������1,������c�ȏN&U��`�H���\���Y͏�3i�`R�f��:�����������;���SC:ŇE5��ߴ���#"b`q�sAD��0RD[�g��=�o�]���pT��p��CЮ6޳���ikp'.Y�������ȟ��.���R�+m�?6ܷ��]!��x��&�嶵sr�)��G{m����pǍ��Ň'6���d����,�ڏ�9�8�LxZ��d�b�!�.&�#���QD�ά�����./���Z;x.�%,���)��QoqR9g`��˼�w���aq���1�F��D�����TK�=!Qz��p��"G3�w�ov�wx�S�/���q<6�1��3_P����7	dRs�Z}\Q�h�SbQAQ/��������H-+�Qt$,_t�k�;�,�1���փ�Q\6)�|�~^�Ӥ%mx���0B\��EՃԉ3�-�{���|k�;/d�aH��*j+��h�����F%��M�z��to��3ږ��W������4� �OQiP�1luM�ʰ�o�������},~@ۿu�>��x������k9�Ô��� �9{Ӟ񋋏�����r3=W�!{A�9�ZVF�W�J�Ë��e�gc�ұ�$�;�Ϛ;����������!g��w3�~1K�i��M�y�
��z5~A{[�gC%�����M&���ڽ:�_���7,B�'��hf�(��{}�;Ds����з��8��f���)0�i8�ٚJw)5��TÍ�s���	�ts�>q/}�^�^k�g1 ��jqJ��k���q���l:~���z���:�y��lW֏	�V�l����ӻ)�4�P�J�(��m��/+J��:�&�i�/�T�!�3�A�{����'������ٕ��H7*�f��.o1m� \�Qk�г0�Q��o3����W�(P�Sg�Ί{fgu��V&1���Q�\ �6�����ټ&/�D�q������T1d2np{v��d6b�E��w�87p�l
["}6��)��L)�j��5�Hr��uW�a-��CN��C6��s�	��vCu2DC~�AlS��_��I��Qk��w�Z���!�Γ�nF±��T ���ͭ��� H��S)0��&�(o�I��sI��G�q�vͯ��ŧ��*W̗�[��J,UIU�g�N���cn���)`<
����_�3T�Kj�.��U�Kaz���E���,�����-���:����o�aKVRE��Qz�篭���8*c��i(Zѧ���*��y߭�}�+��9�l�+j�
�3iy#�lśg�-�MG�UO��cT� ��W	�~���>�Dav�Z��њEN��e�FԕК2��#D�+���aF�+h���梷����2��k�ІXP�te�s�h�;y4ƫ/=���U��c�3��n�[{@���� X�ʽU�@�~�V��W���#O%������K���%L�p�Vi�v~��$o�73���%�b�W˶�`���6��c�J�
Ļ��+���\�x�@�&��i��s��{'v�	������"���š�W�V>R9?%�]>�d#��ߗ�"����}�<[��r"d��'mC���l�C	V���
���,T�?p �щ���Y�	��	`�r�δ��'�Oapw�� 8�6����'�G��d�8��/��w�9�Y�[l[�^T�g�X49̆���
�g��ixJ�cv۠2IYd�Ԅ������+��"�ܼ�Q5�����g�ԡM�o��5�h��aQ/E�	h�Y٘��9q�ܿ$�dJI6Ú���~X�v��~3keW�ͻ�G7�"�R�vL[7r�o<��H)��O��\��-7��@�X�A$�2\H��:�Z�> ��e�R���������:�k���񗺢��l� u��'��-C5�e*L1�)_��s{M
P�$�? �k7k����㙗��]^��nV�N�L�qY������1��C�}��}q�_�v�@]e{�T�I!K>+��Y��S��J/>m?���⊿���a����=��;-@��GD���0��W��-(�����-"R�����۳�{��>Ă`a��0��*�Q�m"v�up"�&�Z�!�7�|w�kp���\8Î�}���Ӯ4��ޕ!E=aY1����U�4M���ꋜ���Yݛ1��$���	�y�i\��[��ٕ�R��������&C�9I*^%��oD��E�{t�
Ը�A��i\�|bZ+�Ŵ�:���^N{���ֱZ�YV��Ɓ����`�g�%��w�N�lGq}��cB�˕H�5l���fzS�@��s@��v�/v,�)A�/�u���zhiq���������ιV�	 -"
�����!�Rae�k���g�w�<A��Lg�?�a
� ��nH�i���j`Ū�7y�%��[�?��"�=�]��s�k�Gzi�W�B[�����#Sr��˿1�bx�.0��ϛdABh*_=0\r���Jr�����U��{� h����!�f�G�>�!�	_Z&�6�h)�jN�� /����"��߿:9BQ6�YD ��'E����FH��k�J�)Q�@�5�������� m>�@T��[ �\�����R���pV��U8�9���B���;O�"�vۈp�`��\�B��!�_�BT�j^(� t�e�i4�]&�u>S��j8�t��TWlW~�υ�ݠS�7�d����T E{��;�/`NV������v�[�]���*j5�������7ɮ��� ��S��@�>G|�^����5���O�E0��K��q߭��bp>����*�ma@Q6m
���^��at��/^a�a��m��@gE�l�����J�N���S�6�Q��ũ����˖�3Ң�������S�=�ğ��ӛ�����b�
f0L�u��b�< m��eL�uY9����a�8�/�J�*�1��E�s�;�����P�k,�D��#����S´,�{��z��W�Z�Ƣ�vW��{~r�W�3M��a0��B�m�*�P�2S�rЬn���� j�?;�x�m�c�\�����`o�<���뺳C�7i�A�IQX[���W�ԟ
�zH�б\Y��©\tֆ��Y!�֪�h�@�"_��g`���O���F�"��P���T�t�̖2�9�q�~L:�Ll������lWVK8-|h�+��sC%�ɺ��pW5������=N�2������S��/�2�'r�M��tׯ����oľ3W��;H�K��yx慼pTڽ�޿@ߢ�E���5�e�X˛���˃t�o�<uZL�{T���c�g���k ��j�oV��+B�{�#V��y��RzIs���<~+D/�����o-�h����,�O%K6qee��Β�T�3�s�j1��f9���J�GS*�/^�d)D��4���fUy�[2��^��x�S�!|��9�)���P�P���IVjE/})��G�6�M��7<=|��l�u]d�߲<.0�$����������$ q�.���UA�Y�_��q.�OX5�R�x>D^�'=��ӶFR,~bc�:�E��~G)�1�~ ��J�� ]��P=ը��V����p�N�Z`�U�'r�i�Q�C�gصid����2|��v�'�+U���Aw����`�),��T��hm�TT�]�윣;����9z��^(��p��]>��Ia������ڔ�%-��Z�&`��ft�^B<�O���S����XU�fqK܏�4�CH~#�!-�P��:}�@Р��Eo�{\�G�S<;mB����5����MS��҂���ڀҹ�H�l�r���r8�.�K�;a�m4&xu(� W:�\rG���OA��e�x��x�֍U�<�9H��u8�=T	6�C|<�[�V���B���ZJ�y�DɭG�X�yCO"�!�7X;����E�r���?Y�us�p�I1�:^��J��Xn�@��U!!�H�}��]�Ъf"0���g��ZPmTa�eX�@tU�y�u6� q�t��/.�[`Wօ�چ��5��9�_�[����"��H@z*�hn�(]���,V�~<�V�V�T�Iw�1�j�;��ȁS�o��}�q �c�&ˇ�c�|���.�ɳ-�H�Oc��!$tQ# $k�{�M���� �Ѿ�λ20�H�Vj�����
���f��	�a�%��F�" (j֢��7��/:�&G۪6��2HjT`A��o	IL���3e�R�Gj�V�'Eƭ��ϲcE�&*���/�x�����À����0���7�dʅ$a.��򺆢�M��Zg��5�!a���U�垛��y�H*i�Mz|��QT��W�#^�*�]egѰ���'�n��2�'��u�!$�3��I�"�����0_�k�! C�l8�#:�T�o�
//�3`-�5�v@�`��n��V�|����S-���`"���e���7�V��.mZ"�����!kI%��M1r��k���G��+ǩD�Z�U�Oև��gf���l;}����>��s�L���I�W��&� �l ��M�eh��Y� ]�#U�H����y%˷k�'ã%+�'���z֯��z�v�b��N�� 5i�N�x��M����~~S��
 ��,�k�żT�����b��������j�|=KԶ)Gt+u3oXV�cɱ�[_�L-*�X�����`��}�̛e��1��En����$q"�:��3s3�?S`+4��]�	�d���v��(*@�קe�[�h�x4����i��x�͡�����U_d��mA����|�g��۶P��)�)�D �	r��{�:R�k�k�5ٻ�W�u?$<����2)����9)8�^��C#M�ż8�e�#��/��(�*�H��/J�p,����ްf�����,�o���C|I��'��ߎ�i��*���2��6��+ATٗ5[�.Kr����x�?��=��=�q�s	�?a�~?2��0d@��Kܐö���t�B���H�T�U7��j`�3$��@s�6nZL�h}]�2�.���ǌ��o���H>���Z9����V�gN�C�x����T�D4D�+���N�]�)����n2
��[mj�FG�DS���"z?��-]U�(1�g�+T�a8��TMb�9^��{&N)pM\Zޖ�]z�Œ����~4��|A��\}����IF���P�����j���>���k��c	��p��/ŉ.��󊝔}Mͫ�)�4����q���hO�y�c'�>%��k}4��.Xif��Ck�bi��Em_���8��h(� ڣ*�bjO���$y��F����U��������*`��Np�9d�7�1��C�0�O j�K�0����u��Ɲ�3�-�Z�d�X���kT� �Lz�/ҜBpZ�m�
R+ɚ`P(�܈��n^R�U
G����Oӏ�]��{rX���f|G�og��鱗�[p�= ��3�ѨV^�����ҿ�T��-V^�����gٻ�*�R�o�{�h0{[:C;2/�PAP�W��>�Q��%������vڷ�Rz�) �#Iy~y�_+nY5%	���s�Ί�w�
q��$�VTz��C��W�t_�M��zN{Ƌ�ʡ���]��D�G$��tŰ��+ކ�nh`��exZ%||�����L��+�1��ݯ��������2����vB'���n��ʹ@6/ik&+���wb ��A��Ǘ�R#�y��xI�Yi�=C�MB �I�}��b��obٮ�ݕ�����w)ۑ�PcI$�VXnTZ��*�~�s\�k��2�2�ƮAf�+U�H�=��d���k��T����� �_�'^G���!e�}[H+&:n99-�/YK�a�J��`a�GM�֪yf!a~�ʇ[NmB��oy.>|�^0�{D�p�С��k<�)#�ֱdk_՞����;��aGK�4�޵>y�Ao�8��[Q��g�Èe$��s_�d��vJ�=����w+,��I����hO�e�0����6� =����e��'|��`�����kS�/��~@x$�[��j�~�l����;�{��3���B�]bJ~�̜Ư����!���>���UGS,c�r6m�xt��y�Z^<^�Lh�G)��]8o�k�W���ȕ�`�JΞRS�-���p��yK���j�r+'hJ=<�4��5�
�:d���,��1ɩC�\z#ȝ�q	$���Zi,w�����0��t%�8+��<Xp���_L�F��v�8���*��q� �c�IԾ�D��SPf+E��+ޕ�{�������ew�BƸ3���ؙ39�3�<��t�b�3���'�@G�K��W�Բ+�Wt!e�9�F �8J$9��R��u6P�R������r�2
i�2��w�#Y����)��=|R�n�q���n)�+��.p�$������(��u��w»uCH��*E*�N{�C\fM�;����n�� �2M�ZS=~��������:��i}�:8R����2%�|�>���٥v:yMmgX�^m2����m�H!���z[Awڹ>�Op�)�堥�ֲ�YO�'���I���AD ��#��~��T�	�@�|L�%��G�er)�j���Z�����䨊���Tt����83/�8H��Gj�^�\���R�=�zy������8�㚷��n�S�P�iKT��d50f��-����������M��R�Y�ۣ��V��i��B��i��n�W�u�x2G8������T��L��~ap�P/���A�v)� 7AY���D �Kپ须��AT|�}�D��F$�篞9�C�+TE�[��IV������y�U�#s]���b���boXt����ఘ,̌���t6>�(+���j(��h�غ*|uT�޼��r�5��3��GyNr��gQ�AKbkv�J���B��`l��Sן�7�$��Sh��lC:Ԃ%?�7�(�v��Q~���IYy�M����9X>]��dЏL>έ��8uO�S���G�&�zP/�L�q@=�'!;ː�uM
rP��-:v��'(��ks���*�lѥ��_g�UZ�gj@����5HB�>h�l�;����{�`$��X�LO
uUJ+�����#A��~,rs��j|�%K �.MGXE�a�
Vp=G�TU�l��yP��BU�3�K��h�r���ki��5v y0�ڏ�Vh\?Uc�6Z2٭]�a �q�p�h�6�'��"�|1�)!�����?*�sI��pV���\��P�bh�.4��S�V\��6��	̇��1O�z�(<�o%�����X`g��<nAG��~����f֪�j��Uq��*����H����z*.����(ڹ�6%�[���ᄴ�I0n��]d��<mԱK�����m�x4+[�J�0���2p���x1=@�2��aq{S�?H��
��<ɕ��T�1!�Ϋ���S_�l�:_�V�
��D8ҡ��Ox���r&�y� `���f�?��A��^$V�6�Y8?����j�;~�#������H�� �,(P�����d M0��.���.y͗P��d��XW{��G|��˥�MI�ÿ��9!�53�y���	m���
�Q��S�X����{GR����'Hs)���r9���(�8�� ֍�rz˝
�/i^��Ӄ0�DnCV��@�V}�O�)���Z-Q��!^"V�Ī/: g�6�å���*bVm�!� ���dɟ�ַ]4�}^_TtG��x�c�M��cP��IaH���qw�Նy�W�b>0�N�b3^�&�b����
���7��*A�jIF��"��;(i�?����!���
%iˑ)���c2��vɌ�"$����W{�^Q�Ӝ�@j�ui�C��exJ��lN�LT{�n��L-�M D[z<�T��eM���^p����J�+��*�8�rTiE�c�]g�so���,a?E/r�`��%ࠁ���T.��_�.��8r������`�&V ���137��4*��<�̼��8[�^lM=�Z�Y�;ï�8���+ qQH���˿"�A�>����פ�Җ=J\~��с��(qDsOՒ}f�>��ԍv8>�B�2Qܮ|+ "���Y�����B��'�Z����.F���dj��㦫�"dLν��b��~л:z^cv��P�N��e�~�%|�Jy��?��6B�[����
�&�z8������U�X�Hkq�p������+!C�@�
��3�T��g�Qp�N�?t��i��m��){��
�%��4���K���SP��!������EAè� f{`9	pN$�E/��Ȏ36}���Q�L�Q�s�M�)�#�姠lrA�o���M�=M@�4�!5���Y��+�<Hװ���i��$l$хln��f/���[��ь*�h<Y������"=S�?��
A��T�N�DjC�/���"��m%+O�;CDsºŔ� ��V�۹��O����>����w�=�8�w+AAFΒ=G�7e}`J5:4��W��ݥ?~��c�\6��L��z�����>߷����2�e*/��u��S7�O�
+�P+Ya�Z4��!�x�WY\&����^W�$��b.!�Y�UC����]�S�G)�� V�����!��3���1���c�Y�#����C��sM�W�
[���{q Ҋ�6�*X�W� }�\����KZD��<��!�]�.}d�F:B�F��d������m[c"���"�M3,�F��t�il&�Q7��|�Tª�;,� ��X>g@�9��� m,�i�jy�peW����ge�A�Nz-���}�}(3�� �=V�>�i�jjwq:��m;���z��U�UAcm=f�Λp#Q��?&(k�XJ��+�_m&74��d���KH��%>|�OG���a
˭Y���vEQI"�K��
��-/��+�~�f6�n	��:���J��5 :����w��s�vk� s(ILS��fQ�t��+m�wzgε-,S45��n?����mR����nZ��t�>��b�F�U֢ BG&��G�n�����Du"���1#jJ-]NLO�P��)�m��}Ge&'��ƈ�-��M��Ј�K5�Ű�~��$v�A��,�mq��*t�8A�B���`o�t%:Y4t�z�'�;�J%M+?�O����u6o3''ݣ�����2��g��.�Wv��L���������҈��]3~���*� �U/� ����[U��z>{�ォ��O6[^Be�<�����9	�guV�v�h���ha��;"�Go�H�_nލ��ԯ�;�c� ��q�d/v�UҜ6��d�/�{2�%)�-l"�,u�T�÷��w�Ey`�K|�4����ns߿�I���_��䶿��	|��:kH~�Bؤz��uD^����Ǐ�0��Y+�ý�SG�w����4�&7���}���ɂ��0$��R�PW��P3gV��ƿ�t�8�h+�P*�s�� qWo0���/cI���`ȋ?ڌ6z�6T]��<�B?H�n���Hv6v!GN��3+�wa��<I��6*r[���pl8%����W�*�v�)���E�`��P��|m�)���u��������.��#�b�y'���B��m��jh��(~?����r�����]�uҝ�beV�<驿� +m�j����`�_�m\��,;Z��T�i�>��ϐׇ��l��fc����&b�T&oNwnH�_�͉�h5~���%�Q��	կ���g3p����[�Sp��d^<R\X��5��m�	Z[���-SC��i����P�O�5[G��_����A�F�_*�;E:��w'�G������B�Zbc�O�"jS�}��4����@�e��9re��v�:�?�`v��jb�q��d���C��m��t�T��P!Ou8�T���.���9p-=����y��.Dy}ԒU�_6i(xzR��"T��ʹosW�C�E�AK$=TOoPs���e"ڇ\Ń� ~��yX�8��[�_�h��͞�AVV��u�1@||{y�d2�dc5>�5U�5�|��Q�k��G�'\��"ìqfö��Nz�Q\�����l��@�A���� �����F�3��҂r�0���ߎ�j+$1�^�B�@�G�'I6�I�ݍ0 �1��-�P6]^���R'�c�V[��{:oK��R%�QQR�t�M�y��]K�u��F�����a��(�G� �/ng%98!�>�kl�u���j���scMO+TJ��g<�����H>\^�S��}�U�b�9�wh�N�>x�m�2���˫4��b�Jt����aoii�!��OSX';.n>\�H����q���QV����^H�o5Z��%ur�¨�C�mh��L��ň��7����W��
/S��Z���>T2�ü*+��{z'�����$E�F�$�yF,�|�C�?�Ԛu�c2�*tn-_���9������׫*V�=1����}�4��Ow<"�,�8xI��G��+�>b�U,�����h�ߩ�1uo""�i�s2�5��*Ƒ�:����Cg�rf��.���-�R=lOg�kI������@�1S:��.�0��i3��^\��<6-J�i���n�����1��~27Չ9���'�s	����)�p��-|_YP�%.�2V�����y=��N��`��d� �a�]�������3h�n��>��(k�����ӂ�}�	���l2y"?��!�5���B�'���U��>[E3����%,�TN?�0.���Ey2��D��{�������\)�S�$Ïۭ��\��z�py��u�o�} s�Q%�NN�"�5�#�#��I�Cl^@AFK;WLS�%�1}1�@Ց��,�w���]M�į��W�h#,��b�����v������y{��sZ帍dC��w��Ic27]�\���$Zh����K�W�$��2颐O�b�f��˸��y�go�Q�۾X1��F=<�A9k5(����n���i���v,�wo��+[�+�;}��e�S�Zt�㎹7u/_+���lJ���}��>��)���=
��4jY�z�,�$�d�!'�D�KS�<G�XI�ؿI���[b�?�lwۉN<�|^����ٺ�xsw"?j�J���c��Z��Ł�tJ_��"��̼�9��$l�\\:h�aǗ���LZCq>����)�g����G۫�$��/O���j������c'br��'�M���3���{f�rGyo4=�D�"nۨ70������|��{E�`�b�ł8,���}�LN%(��Z�ҁԝ�o��v#L�['�#�#���R�^*����s	d���(��f�E4�zq3g$cG�,��I#��<���T�%�?��Be�� ��,����_L�ҺUUa��co����X0aی���W/�w�.�������`��@��Tu��l��q����I���kd��#Qq<Y����-R�1���`�#�JpaIҩ���ƁO�v*)��{�Y�w�QS ������2Ň�m���Ȕ#8?�s<����V�$�(���ũB1Cu�Z���,zAf�:�.gt� H(ֳ�5ԃR=�>�V����c�d�[*lӶ��N�$��9��w���w�����R�%�=����W��![�5�����?Z\Ź��5�ʙ�w��Y�S�ӳ�u��,",��{\����k��e�rg��I�v��ޝ�bↁ����o��R�!+!�Mk2Pp0�Y�X�|��NH7�-� ���i��|{�_���G�b����o�_}J�P�����ΟHr�t�Z[6�K�z��_�RY��x�||`��Fd2��M�L���Z㟁T��4,v��
����[7K���Y.k/���¸ �L��,�g�8,��*��ZM��x��)�R���Z�qٚ�<�^��Q��v�4I��©��P��* �؜pV����
�Rǝ@�	��s �X�9-{�ΦûP�v^a�@3�݇ɩpU��a��nL2�9�2%��}�	H�&n
#�ō�L�P�ֆ�G�W��q���R��j%r�O�g�s�>�>3�G�9�t��vgQT����}���s"[�D���֛3zB��rr�&ˁ_*Z�j��s׫�K$���7��S4l�yql7eQ�m���Q��x�Q��u�K�8�N����fi�+x@T/�ݥzA�'#�5M���A���x��{*%8�D��5B�Rs<e���u�͌I�g�q�y�D��(�;&KX�V"�n�L{ΐ����v�)����G��ٗ^�;)���� �8gl�"��e`��U�g�偑ۜg��Rt�Ss%S�+QZAf�gx_iP�1��)�#P�+�75����`�؂Fwx��YCz8������W�'߷#����=���%Lw�Ҝb]�(��0�n^���/��@[�ܛGx�~�'��Y����	��7.�����Wju���=9ٖ��F$��ڳjTj=��J���ߕa{�wmF�R�Q�͹V��d���ħ5�;GQ8�o�iDC�+������짞��:}5�S�z(�bPZ~/`���]X�0���r
r�&��h��7#:啝���iw�b8?~�˙�@�w��s��e8V�lK��ǯOH%�#�����d{�m�?�`u8~{6]�}��̟I�������w�r��2\[Y�{���a��V��Uڪj�I02D����f@sͺ�
�pLV������&�B����J�]U����z|���x.FE�v~ ��*�5� ��j��>#\5?�ƌ�l�u8^�������Nob��1/"S��/�}[VE�k_�t>��m��xta8q4�q���ϫ�_Lv���FV0��E]{�[Z�>ʶM��քӞyc-�u�A�8E�v���u���b]A�k��W㥯�|�n���@s��0��50�R]c�J�ظ�_����i6���'3e��c]XO~���wv��2�j�USn#*�D����'��o�|xdu�=��i���hPF�Z�c����Cby1h�86 ����ܱ�n��So�P�,���D�tH4�
�4yƲ�%���lTIQ�v�Õ+"6ϲ������ dt�'̾��������5:t�W���=�w��� ��/�	��ۑ�XS����Hֈ�ܾ�ܓwo:��GԻ�&i���Q��{��k~�j���X��㈏���?��SWr����<.A�:��u/Fue��~�詯���')x?TU��ҝ�OH���M�E �B����#s7��Ȯ��v��w�������a�2�"E�k*��n-�r�=��utS�ۤO��	'5��y	a�'�9Ai��8��hM�p��?�OP�$�;Zo�c��}��߾\�ϼ>��O�^���� ��w�n�B�Ӹ�NbQתHe���G�����1=�U�+wN��M��#�Tq�q:_�q����ܾқ�P2��	���)7�-�V+�\��q!󾘚JՄ�3�`B�,�p�
�mrAB%g�M+1%�����u�ˠ���S	��ؓ��~b1w�ę.&{��<��I��"3{+7B������I�1�ˤ�P��M#f&���'.��.��OƦ��9[Y��%۴Ќ�ű�K����-�lŊūV�|I9VHNd��7�'�cE�����{�'�.���_�{�6wT���L�`d9�\��J"�*�XЋ$��$J���C�0)N~�X�{�0<��Y��Y<��m��k�k�w:j�yI�\q~���_�/�Ӓ5��UJ�@�̏�Bm�a����^�gC�+B4gs!ĳ}X���P[ 5�����!���20f?Ĝ��On:V��9��(Dԇ��`�?l(��G�j��D�^�#!Q����oy���� �+e	?����I%d�q!-��{.��Bs ��{�f��b�e�k.��Az3��ב3���d\�����?����[i\"N��E;`��ߟfQ鎬����$pS�	�+�Z����8��_z�E|5)�.F|�F���`5*��H$�����p��b}�u?��t���S��c��6~r�r�!�ۀ��!@�x��	�A��-�'~*��azWC�)�|>6������	�R����Q���$��DV���`ȱ���w$O8���Lb�K���x�8�������p��
Hۺ�:byș�Ӓ���{ҽp��Q��Of;�&�T��v8͕w�[� �X��9���;�O}��g_�D���ׇs!F-5X��?����6b>�K��妘CX����� 4-�&T�ਹ?h'�X�08wDA�$X�3��+a�s%k��Z�@ଝ��>!o�5�1�46O�
���FuR�����,B�@UHc�1�r0�(��Y"øuP/.����>��Q�S��r��8y���{�]t?��v-��g<�	���[���w��?���<�y�Q}�Zׁ:�%}��?���3j�8���]h��7i�SFX�&?g�GEs�����ֺ���{�!���L�Jo�2V�3]Ik���2���IN��	8���:]>8�q�1a�pua�$��"*Mr��r��Ls��[���?u��(��-��u�$ި���d�M��N�DY+��A���4ōC�z����X+]�*���o��b�]�:\T�e7��"_����̖j��@m/w@��д�G~q9��A�C�1����敎EwJ�l����	I@T����G���p�\�U�y���V9�8�W��,�?�~n�QA����t���3�W���ۇ�ZJ�k5�YL������=�(���cL��`�TxX�����w�nG�~��:�>��سb�[��;�7����_��<E�yں��t}x"�x;ؙ>N3u�n����s?]�0F��L�ʢ��4 �:����ɏN����i8
�v�Μ3C8�۪�(lA1��Fi�F6�Ϳ�q�p���lf)S�Bk�l�:����� ���WT����v���;� GHl�K�7����Yq|���/Ӱٍ|����X�:���b:��!�Υx�6Y��c@�%4����,)b�=T�*$�.�D�Y��h{L��yW���׃�*��]����&���F"K6C�[������A�i��8H#�ן�O�����,�&ߺ�'�����J�
Ի�l�ΖvO]L��܉6���!8��u,��z$���JX��;�J�uA����І챖B���*�c��S���?��v4�M_mŮr��KB{�|X��I_j��9U�p=zZ�j"��=�n!��qlf�w�~���l'�H�XXۿ�����ぇ�>�k.��X&�Ιa
Tu�csr'��p =���#�g�{X�o���rڎ#�י�������]O| �!1�@D�LR9���-��e��0��ict<�]7��H���H�O���������)Q��~�$���?J��#��5��E�����]�q(Eވq��d�2���[�h�@�9oS"�<=���f�(/��Q#�Vܓ�J~�t>�Sn�-��L�!X� ��(c~������jHbGe�����v԰��cc�^"��g�r���K�Ɇ�D���Ѓ�JyA�ri�C�C<.���B�$��nRȪf�%Q�f��S,Ƭ��j��3"�51��z9��_;m*~HQ��n���CV����C���jǝt�w�D$w��9�T��y�}y�@g�T�<���չk1"M�/����\�`�8Q��~t8��S6
�/�Jn)2���x&6�I���`?G�S� +�g`*��_�{п�"�տ��y���n|˶-"�g���#��0<�������Mp9#V2(ջ�;d�K��TU��x���-W6���}��={}��� �q��zr��OM7,������\f-��.�P��E9��uxI�x�Jy��Bz�U���_� �;s���e	�:�����L��o4��`�B�������[(�@(7�����ȰnE�n�۩p�J[Kg�:T���Z�%5�K۷w�|���8}�a�9�����#QΙ�1��fqۺ���9�������͜�j�����伓�g�5�-�U�1�H���;I��	���y-ɝ���cΈ��{(|�a�n:3�s5�M9���v�V�����t�R&��%rT�C��!�٭X����Q$)^��j�w٬�\��"U�F1�����1N%�o�����epN+v��\(�L�:_A���&�AG^n���[�g��_F:���B_3�A��G���.�1��Q�`氿)z��ij4��.&���鄋ː(�!?L�T�&�Q��X
��:{��ڧ��C�P_���������5���q�����'^�F��x[w��H�Q�-��J���s�ns�8�O��\y����mu��=�3��r��Ū��e#-.���i����D#(E��-J��X�g�1�L��sע��/&�0�2��o��-{��FPF�#XU�NV8�9م�&!��u��a!�y�+�����h�k^�q���y�_�F��q�lQvW{�Ҙ[>���"����n��l��~	�����YB������|���>����=����Ԯ>� )�P݃@@�mO�Cx��H��y�n
��5��,�(M�뎽n!4!U��=��$]�P����R��F�)�/-U"��R�k��S|���HZ��_E��ȝGI�Źꋘ�;\�l�Y��Aܯ<+�u��@�9�x�*�d��k�/��:<���<��v��	ww�Mb#wv��hNq&�#�uڮ�#å2.���M�`�E��پ_���� u6n����8�^/_lݱ�U[�i��}��P2qi�����6����U�?���Q�B]A\��LM���=��O��ݷ�U1��A��v�.��+�	��-���p�ȸ(�;��ɰ��6-�T�����M��;�5&����z�$��2�װ�2�������p�2�(�QRn��,F7�UÍ�fm����hϩRs����Jy���� ��^��������-p�
�bS��H鴐2r�����Q����T�=��J,4�H=�tJ�ߚo�d%��;�-����U��ï��=�� 4	 �Ϲ} W\R-���+B8�)��׷$��[�5Q������)�{&���������*̝\���ɘ����L}��^%v���+W%&4�m��+�$����~�'_D�����Ǫؑ�pJ��zЮ/կ�mðq�Y�]�p;~�a�!��B8��hu�!����0�jWcS e�{�����a!�/��^\�6�4}EXP�ߒ+�W'��ƪ��mOt�F�4�Y�������/���g�!Z��tPu�3�/�kv���
r�b���- \�� (7s<�֘嗎[�����������)Uo]�	�D�������Q��]HuT���"0���4j��?I�%�QN�6pZ��ϵ7(�(��7D��g�<1a]E	3��M�������:�\��y�|?��3�]�rA�7L,P��L��Y�FC8����/?|��+�N_Bd��ayZ�W�B���b0;GVPtY�v��f�i�w���9پ��O�Ja��`�~Xjt�\C�}�qY@7�0i��>�̒μ�}�F�h��6o�6�ʺ���)��v�@����s>�t���t�0�g�6�N�Vb�9�e�������AΟ]E��Z�΢.��9���)�Z���ѿ��u����l������:L���g�l�V'\vCv������D!.��$#��KRX� lo��M�q&����`���6s]G_M5;le�~�w��E'��� �E�@�V��r���Ge����e�B��P�+�L"-���:��(��I8�k���Yj�m����"�%WSt�]ޏ����n�6��A����"g��Ĥ�����B�G�D;>�9�*ܓmR�ѪW�;��
�L���H��}+�蜅�e�S�����>�2��V��"/��J?zI|�~�֝FD�ݏ�crK��RBb���2ɥ���:WP/,Mډ ���F2�=a4z�*g�U:4u4�.	X���~�$YV�Ù�5��]�A|�f�e��{9d�?�-����/���QA�t�u���@��F�8�+�>��䀏�Jx���D8��|��t�	[���H���P�V�Va�f�Ll�u��,���P9�+n�����f�3�k����k4���;'.���҉a �L��3��U��J��h�'�����l�^�P>�է��Ӥ`� 0�����ΛN
f m��<���Y��ױ:P�S��ୂ_��b �+�Cz#e�3�l(���WM���X�8"^��h��<� �lc��=���o�f=�) %�5�2{�K�9��-*���r2wJ�s�7��ڮ�i-�L}x�� L������>Y��G����٢3=>.{Ȓ�N����f��ay��$�k�����2a�$ٍ0dA5���t����.Iq��,R=Oؕ���}�Qt R�x[�Pd�FTc@5��X�!-u1n�:���}�`�jT�
� ��f@9�����NHX��Dh���a�<C�x���4	��J��ء���u��˰�d�F�����q�f�^�"�ϢU�k��?W�@뿤1ρ�AL�<�i�P�iS�:vM(�j�������;^��B� �Cc ��&�, ��h̚,���ȝ�`�5��A΃���^�G6��� �.�ߡJ ��ۃ�0��2��ވ��VF�޷�n[~OX,+(b�pF���ʕ6a��u��p�,�ː���IC�Slw�d�� x�a'(=�A*��1�"/1/2��.ż3�s��6����#�;��Z�m����[�E����	�m��N�җ,/��i)�7���K@��j@�9r�x�+	����+��4{$rH�BNe��^���
 ��aZ���S6L�պ��(�F�v�p�����S4��f�JK��Be�M�5���-t��x}x���O����X`�6��!z|$�YÛZғ�J�/���cC�.U�e��4g�DFJ�z���>�A�)P����[(s$a������q��ɔ�X�/>�$�`7������ݤ�WiϡB|ՁL|XE�蓉�S��՘_[��Dg����H�E�['	8�RB|N�Ω�m�F�Y	[4����X�磂�{�E�����)�[G�;3�#�fn0��>f_ě������{�i���̝� �o�ƺ�1�S�>�"��0]�ı�.�%g������:O]>�d�!T�:͈Y�Z��@
C��u����y\��?�d䦴Λf��J�O.ݖ@�/W�i���a���.�O�D�I��I�v)Vi"�����Kkg�;�����1���G&���R�[���?h���)�Ò����C�:��~-`o�^�9��?G�|5'3׊���04�a���C� ϫ�FS�\���ί�@�� ǘ���+�3���[	�͜�%���
��3Ԕ� ��iPU�'Ǯɨ�a�c"����ir�!���m��pc������2�^y��6��[~]���F�2h��58!�|�3� A�������$��̼o[݉��4���_2ViZ���t�`�Up��1:u`0 �ʿ��x��W���KGB�(����%n��)��нQ*ǫ�����>)��Fk<_�(6��ϡ2��xD��]���8�D��Ti��͉���3DQ�>��]?��Dz��&��6�{�C�G�8�����[ k���l_����*�@�����0$��!m�:'F�}ۈ�x�#�ʇӖ�	'�	��rg!���[;i��(~��;�EI�Plx������rU�����p|�/l�����f7����s���R�2`�F���_���h?%Ǚ1g��e�0d�P���s�[#O��e�� ��X����L��cr��:p��O���T�>��Q�*��zq �a`��u�����ů�p�?�x�5����"�v\�6͠�N��y��eX��^_7N��#�\.C1��H�?�;���)Ҳu[x,GJ$H�>��&�g�r>�f$�%y���`�8�K��~��j;9K�b܄�ۇe�TgE3ھ�H�<kߋ����Tqc7k�%�$��E��C�OH���ڊ�<'�K�'�ȕ�i�|;e�wB��'�r�6x?Wè��I�z_8�a�η�-SuO���M�7��Vŕg��LrR��~P������-�9ث�n�}mt�ȇ�#ڄ���L������BW碗��;���� U�$�9!�&=�~����� �wc$7��"�M��8oM"�#ւ�*�ϛ�� ��؝� WnE�jK��=�����I�Ļ�F�����S����Oe�-ˢ��B�Y�n�1���]EK˵���0	�e�$��@��.#+���7mT�^�iZS���C�1^��}�|$�%sV���ؕf��-$��7��3&@Ui8�ƾ�j/V���������7����~-���zm��Y���n���p�n�m�y|p?w��''����F�G�������wH�	�W���}b'�>;���{t��5���2V=6.~t�I���/�M��QK�,�N)����/�0��Nۼ�������u�B.H	�6}���^X���~/v�$'x�T�������to�k�#�^������7�2Q���/9�����\y~)D�欦���*�Wa����3��xj�YE�Ut)�w��R����8T$6���0�"3B������浇��[���-��'���)����!��y1����r6$�n�ֆ��y���S��Q�3E�R��[!8ƥ>�/��3N8�p�ؘc@bJ��r��	=F�+��}����12�"z���X�4��i!i@����0�	�B?�1-�F����dt���:d�m��IE�zb.y�P��}��^��8?q|N�(?�җ,M��p\�
�AOw�X$T�.���	�A;.�������yd��2#�07-uF L$������BI"���e<����<`���SPLl��qX!.8a�Y&M�o��.p0H�6kz�L�|�}����Jyek>�����'�F�Cٞ���r^xC�RJ��RӁ�~ v�ܮ㉰f!�zH�����W�@N[�;c�-T��Y>ѿ���G�Dߙ�I�_O��)�����H=���I�|+��)q�cn�<���Y���j�E#f�fف�,���F+�=F(t�~W��IKQ�CO�^K��Z�0����ߍ$��H��O�i
Ё���/m �6Z�:��`�OI�o:1*�El N��@�d!��3������z��ܼ�%*�+��(<j��jE�B��OH�e�y�x��]��վw��$Tz�UΎ&�]��<&��P�"ow�%�+>n��O
��Ϗ�1�B�x$w���E�4��eO��j+q�����ok���yg~>Ep�'�x�0�B��8�V�֊u?."��9�ܑwO��0ʼ���G�<*��=�~��Z�~;�6����[���rf_�S�
3��R.������M���"���d�0����R��[�Լ��� �r0���~���E_���K�NQ���&�������O�Rqy��O��7��Є��|(V�Q�L�2y�Ns�e�&K��\������sL��=�_�3Ԕ��o�x��]D����9K��Q7�(�=Tc1�'4�zZ:�B�hג5��R�X�C1�Li���	|���og~�5�	�/V����n�������c��W�z������x��K��U�i���c������;	N0�� ��_���̧���n�U7�#���n7p�{����b��y$ʵPfuw�.
�)�
ODaY��/���C��Z;�#wS��cj]/=�E�A��M����t��T;�P&�4P�כ��|8��� ����5[[���	װ#���ɔ �o�#�a���O	� tz��:~,�y��Q�	�H�'�be���y�4���Ph�NѥR9	+� �����pڄ١X�n����g����+�U�������Gah{���dB� <�3�ZM��)÷���#Y3{sB
�����k��p�}�Ŋ�y�6y/��\%�Y#�
ť���.��A�(0����� �% /؏�o�C��h����ǌ���6����&M4��m����Z��Gۈ�3����!b��Z���u+t�3<����|��sG*5�~K����<��ʭfs�I�)eU�[�UK�T�B���${t�㏱��c�T�F���1��PZ����ڕ����E��ԗU��Zad_�w��.�I�> z+p!'V��{�OA{�=;��v��$%��X�Vw��{3���R���2�� ��c��q��5O�6����(�����y���݋�Uc�\V0��� �V)#�_z+���'�T}}���X���!��O������zU���֧-�UhO6ō[���A
��|���Pndd#Ǝ��k8�}�V����z9O%^�NmU�;х�ŇN�C�2Ձ7�����d���1)#�Ȼk��ͩ/"sCC�2,�2��E���}@7��Mې�(�h0� ��o�]\ů�r��g|MN�SP���/�۲����A��r�@�I�_1"9��{)�g�l'mč�3K�Ic�
�6�s(
���a���˿��Y홎?��G\Z��P��^ܣ��%�jk0�&,!�A+n��ٟ�(�����=�-�żS-��x��X��1d�~j5�=�Zĝ�� E�e�^�{��ty�JPUz,����|�N$m�W��:_*�	f��w-DB-�}�l<{尻�<�3z>�˥S%/!�k����<�Y_�1WUʋ�ͨh�8쑽*�;G�[SZ�.����>f�?jD�N�m�k�5��,F���?ە�����۽g���C�3�wN]�Y$���bPOY��n�qڪ���4�/��1ـe\L��Jl�]���#�I��'t��؏&ki��Uw�R��)�����E}%��QG��Sp4��M|�&w��[ͳ9+_A������j�eڽ2�E�q��L-�l���&�eBU �#w�Ϊ"�Zo_{�Ck:^yNXU��kg��@U��pp�w���dnr����K�M��e{��l��i�e�狛��c�2,�b��w���d�(vQ/Ȭ�
��ƫ�@y�{�^Wp��}8q7{��!<����.�g��
�K7|dH����*̸^���\,��UC��q���P>Al�nڪ��o��[o]�k�äH����2<�:��RC<~
u�YRIeY�C�B\z#����1���1YW��ǡ�(�����١}.�"RW��I��%3'���w�I�J�Gs�SQ� ,�a�ɢ �������S�^��N@��_�o�C�H��K	�!p����s�1�}��]<߯�5R5Q�Q��	�a%!"��ϫ��Y�4����$�R<�z�[V4N<h=5;v�St��߷��͇���<Sj5��փ�ެ�ߛ� ?�e����8>PCݕ�c�jkU� +���*V7h�_A��G�}j>�j��mA�YF��&L9� �b�n�A��h_����r�D����囈鯊��1]�״�s��o���Ƙ�!=L��_�Ү���5�^v� w����f}�(��z��Ş����E}5��&۩#�lC���M^9�`S� �ZE�9c�J�s#��s����)�[��1��`�,�5�n|�N/ -�$Qו�5�,����J͒}��BN�B������#*{�yO��2\:���ˎ,#�d�6Un1�?ߦr�����"K�j�	�~���b���i�9бdHe����a��$��ґ��D*W�	s�a��@�o�V)���I@C(\cb� ���$�i:s�����採������ [O_9Z���g=bg+�|G=Qs�~��!�@$�3�!)7 ���i�o>%��j�I8.`�d�5ㅚ_r�ʾ�_؂�:��qW�����[�_Ǯ��V�������ҧ&��j���c6g�{cSfܸ��;����;	u%hZ��h��V�]�s���¡���Y�T��2�gQ�w
/����Fed�2XJ;��Nh���N
���.�I�T��$���p��E8�P�@����sy��<fUC�ۉ>	5�m��������H����.t������d/�����ÉG��(Ћs��9���,-��Uݹ<n�_��wS�9�L������NO���Z��u�� [���p���ą���`>��Օ�����z��a����K�6��nq	�8��7�+3z4 ��1
���0��C P��z~�]�|��i.�ww �����3��� ��)�$����ը��n�?��SR*7��y�E{@;T3�v3�;i�m��*���_��J���Pl9N�{��{ʬ���8�wd�'����>�Mh(o'H3 i �L�q,�_��4��#�k���X7�2��d�UqE�~dY������ϣC���1��oYK~��{� d@$7Ъ{��� �]��3Uc�w&/yك)�Ýla�����O�����P彐7t:1@�/xz��?�s�3O.�"�@İ�VJ�r�Z{���)U�G���O3�#����Ϋ�	��h�JDc(lkt9Ey#R|��3lƄS�型9�Z��G]�?�S&R~M�O�K�I��y�Ғ�v� �+k�L]G����!X�V~^�E���"6чo5i����d`a���y�h=�E��1[ҭ�$C�N�}.��OZؙ�8?��-M���U0�vJi����/�Q�l}M������\9B�ۮ��b�/�s��վ�aq��Я���Nxt*S�X,��"�}ྴ2���>�D��nd��u�oh{�h K��Vi�][��e��W�ɍ(�E�.��,;Ɓ�g���>?�4Y���2��ݗ�o%7�95�0l�����P��=��!�`!�l��P���¸�X�^LX2��j��9R%N���I$z�W��qF�8��U�0#�z����(;�h6޶��n�IM[������C��)�>:G!7m��Hd~^�uu]74���BP��0� m�)��L���%��Vu�x��?;b60�(�h�񶤝Q��	������_Dji|����e����D�B����W��9f��=f�ΦYF2>�����/�/��@<w��3�������k�p%I��4�L$�tr|��I�C�^��H#4i�iv�:4�g�o��)���P�ʓ�f���R�<����Z��Nv�A��&͊z�8epP�x-8�ё0���j]�l�s���?y�������I�R�R�Z\K���bХN��*��*�q�z�4tC����]{�-�SZzp�+x�-�g.�Ӌ�gF{�3���	>��~[����nF�����A����&��
�����Xi��5�)��]ƊI��EJ_�h�8�*_[��港B���,���M@d"���>ԯ��XDJ�����障=f�zBw���O��Ea4<Ȁ\喾>/��I�rj\�i��6u�����pu�:���FŒ�S-u0�kW1�{>��8>w���񄷆j�p�r�ja�Ok�<��ćO��no��`?`�H�ǐg�E�筠���E�B*��*��᧰5~G��/�ߑ�z8S���g���PI,��,Åa���H{}y��1z��Pf����{�q�.Ҕ���uD�nHځ��Ni�.㜢��ҩ{���$�����Ni H#U� �����`��6NY�U��3���m��c�ws׹-���������~�M7����\������ ö�֚�'�S���g�,�k��o�+��ύK���(y�����S���vt�93C�b���7�4�*�)��+��ߓ��5�Ж,�'�-`q��o�,u������.�����}��	R㤈�F;��Be���mK'��Sͅ�� xY���T����㊂�¡�_ħ��;E .��1c��m'?�@95V=	A������K�<^J�Z���kC�c�7]�s։D�;�{�[������c�� ��-X��H���p�$�u)H7�+P��?��^@��0����ދ�j�C����Ҋz/�/�n����D��'�,���8��)��N�]b���Хo���{tmo�OaG����Gŷ��Qe��җSΓ/�r|S�?|��
dقo D'9�	n oN�q���_��@�t��=��ыq��+�
:�\IQS�r�ۘ��`�#���Z��!���9�Cr�?��!&x�ؚ�?��"�=������I�"�r�s�� ��o�!�p��t͇t�Xr���.ԕO):@#D����Y)6q/ο-�PU�w��AxH�����5���"vQ����;y��̥'�b#�7���|=[ۮ��Gm^s���^��
�5��I��Ru*�"�'A??w.v��pn����+!��o�y��@��j�b��u��ڜ:��Ҙ�zbDJ�򼿛/��/��*E*i&l��r
����hS<��o`�QĤ˰��׉i��)ҭ��bŀjߑ�s�#"�$�lw����gS4�x������UyEhvA�Ϧg��xn�1��mҰ�=�Y�V��LTǀ|BNͳ��V��c������V�835��]��ܮ��Z�����l����u���S6��<Z&7��b6G'R)$��yr��"��o�͚������)���Wr�+�>Ms�	uX�[��W�l���+X���ӈ��T7%�V�u�m�B�0} ��Y�r�<���,�a��Ŗ1��~\1���R��"��+c=���Q����m��שo�3:(c�y��C������ֵ��	H��~5�#G��VM��t�J��/8[(7us�j�.++�f�����O�%GB�:ұ�z���&�e��h��@�%��ó\,eD
��[��(���]F��I���nx�䢴16�`1ٗm�>���[�UHÝ��oH��7�"ί�d�ä:g�Ȁ�ص罊������Q��ߋ�����8�B�ݘ��ɰ&�lD�s���i50�%�c��Z�q��B����k�5�ҽ���%6���V���	SI��㛸1�qh��^�:L�r���˖S^�w\Hz����^�K�M>a��s��iŷ']�b!�P��1zJ|l��W���4ʭ��^S�"�����6ɂ7����0���A�0�%N�gT����,T|�MMHN��w����rH��boTW�b0�bC�����b�Z�yɬ<(�L��u�s%A��>M^Qh�@:��$�Y�f{����u��/nN�����%�>&�:����`<a����l��n~Ӿái$k(�0gol3��&��lʅ�>R������8=_��4<��aD��nLSeO����QG�/��m?��9"�.�8�Y
�WO��sL��*,����� ����B�f���|3�|����a�2�ۓ%��q�ik���Â��*�{X��h����8��&�ц�N�s>*	��;�֦Omh�u|�Hp�QFUˑ�毻�t��e������Ӫ�'�vuՙL�f��>1";Y项u1ާ��kD�򌶱��lܙe?�`�|@�9�W�Je ����;Q
x���ɽ����'W�O��a��A�ލҍC�:s�Zw��W��zV��C����F(4�JV�'D�U���|H�fí�҉�X5Ȍ�נ����#/B1�I�U�]�dR�}}�[�H�zSk���c��br&o�Ɔ�d �8��/^������޺w�© `*h���=��0G�n%P�X��C���Vhw�8#ҫ��2��{�Z����/��- .�g�Q��܁����H�&Y4���Us?!%���Z��!��1`�/�	|�T�0E�'�	?k�-�y���(����!'�B[�Ʀ�n���b��?U�N��h$�����n]"�<wR޲��
A��{�^��1N�佒�\���km��g�%�����-�Ac�Յ��6	�����U:�$���B�K�����꩹��wڡ��X���c����̽5��r��!����u�ą�,��޳oo��<�x�T�!�@WM�*/���l;���,�a��0����p��U�+�4/�3���;ݨ��@�f�%׻$���#ы_ �Q���?�V�?��* ��Uis�G���|r;����q,�M��O��އ��J��͚�Q"���F�[�* ����\�i�Z�t��_0�B�b�����z�% K>��f����Bp�
��q��C��l�ŮY�]nAj���	�=W_�O�1��ˑ=<��V�gY�*�L
q�����̷Ҝ��T�x�����ٿ�l,Z1WZKO��H���!���3\�f�vf�^�'�sP�����f�+M��g15�GK���|ش�r(	��N*�_՝��XCY�bb<�v=�a%B