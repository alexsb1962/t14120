��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������U�#R���6k��ME�,��,5K�7Ey�S��K�s�p){�N�ǍB����dq���࠙F����gI���Lk\[%�D�8�I��M�!�/�OWb����-r1'�j�4]O�#�8k��Y��Z����Čt�#N���Vખ�ԛ1������
�hlp�l]j�Z*%����+:��������:Rzz-�cg�����sԺ�h5}�XE)�Z�cI_t�q��$��Aܸ���L�:��O|��<3q�.�nH
��LW�����J����[#����:I�}��\8ΨxY@�LtL���^�f���X����v�4=��"�.�'Oˍ`2�����[`Qe�$�z���.}fd�-��kKmǪ����N���\�;4'��]|Biq�����ϑ�n�|jqm#/�вYm��>���ޠ���M�+'��*�W��i�e ��!�V�6�ad	[��K���6@�ni��'�+�[�q;wo!����Sա�$���� E+��-�tQ��Z�5B	;�T ܁�s:x,�����D���`e�N�g ��
�@Zq���Ň��>��-6ݑ-`����F#��W��5���Z�b`<���ӭe������H�\�j���{�'���S`���B
dpYD�u��S�χ�m:V��w��0 �`4Lpv(�Of^y���o@t��6Wb�]�?��!���K������y��������������We8���M�#�z��˔���*�
.�F\9[����i���!:�Z��R�@=�>�O�Wi�E��b:d�pZ�W퍣 ���b}Ӓ��[�ZD�'���ɇ�&��;�,4R6��,��ͧ!MOm��j��|V��K���d��[:y�H߃��o���I�ԛ��y'�VS�b{���V;�����y�o�:X�$<���qŜ�6>��o���Dr�%'y�	�h�jy�=�]�ze�W�*(�4�q���A��l�&$��l~�O.�r0Sk�����Eml�SΥ��}���gH�5 �&�V�o����>{���vk��sg~�M˅���L�R�v��X\�~t�@u@4��Y4?����
�A��d>D�
Z�p������7������E������}@��+�}X��2���3�[��"�q�J�9\�C{yV�b2�J0���#F��N` Z�?����lZ�5 �.@�l�aPn+�d�����U�	���ea7ܵ3v�N\RQ3�
"�:%bC)�o]V7�M�?���e6w��]���fgj0�e9����*i#�tUf����:�=a1�x�A.k�<pC�@B|ْ���+�N�^���e�eB��3�Q�@���1�p����HU��d�14O4��qD�$\�K*L���W	_�緬��[U_�1��4�lU~Vh�M�L�t�}N\�Y���A��+~�G�׷�I��	ʠ�������5��'���-�4^6{.1^�CѕkSIM.�G��H���5�q���"G�[� ]e��är���ԬO
�le����FL���i�Y&t/*y��Et��d'�QygL�f}�s��W����)eN$H��R�p[���R3�,$��eݪt��/�_4��@9�e����\b���
��KϾ�����o�4�>�l�AaK���oD���3I�;l��[cՕCu�guDp�J��=3M�9G���0\(Ұ��D�"����}f\pQuO]���$�ǡZ��-�p�1[�����PA��* w��c�;Gu��.��C
�6��s��s�����o푈7Dug�n�X4&U�5W�������-+-�����,sK��`�`�j7�y8����ʔ�E���|�p�1Yt�i��\ua]%E��)�jg}�ڼ^pY��}��=0��1�o��h[��F����6C��Q���3XOٟ{�5��'}�א��e��ȯ~�m$.���\�_���$,�l	S^�Orwe $�>iQ>x7�ӳ&���ɻb�[}��:�nj���1,���Z��4U���2 紬�K�'MTv@*�����Q=��*5��>>���NlQF�����s�"%9��r�����Z����܂�^L7��l �n��yx3d����h�k$��B"�sOK���M�%�H^���y̲�R!(�Ҳ��`�Ј�]|� �f�wi�<�-��b~:����<w����g�.ͭ���~Kp�͠��f0W_?Q�ckL$����m�|��>�@Q�Uh1��F��T��ւ��k�0��ٽ�Jw��W���#�1y�HK��NAb2f��.��D�����M�-Iz.6q����3�I딡�����++�hB�B����@a�e�Ky���KZ�EA�`2c��핺��e<�x�y�g��L���4��e��^�� eߜ��̈[�!$$~bн�V+瓿a[�0-����>A��&OoD� F�
@.�s"r�l�L�. @ͻN��!��`kH���j�?L'+���ph��jC�������XY��v�0{�#�H��#�Y��1K�bd�_����[?��Y�7v��S���{�8��H��^N6��9/��T�1�����&)������k�9��F|��L瘇�K�ނ4��N/z�Ε�}&_~=�֒ײ]������Jf��7:Nk��)�ؓ��,�!71_�� 2�99
[��7\��X��N�lB8B�"ޫ�g����7Ǟ%���C������$��_F��}�yX���ǵ�u���*�+�7� \�?!-
�5�)��ί��\@^���H&1M��⾎5UA�W)��}����2	�0�$ vzE`N��O�hX����OŶ���O-5�/�)zV-��G����n�����hX��9��q��:Z_�z��/چ�;��:����d@rl�� � �"u��)�R����%���Z����}q7�HZ(M�EA�#	4�B�z��O>��U'�s�nns����!�+��^M��Ms �V��ڐͥ���=sc�SY�DWf0{'��Fu�A��u�8��u�������.ҹC��h��J��b��t.)�%h�Ft��~�k(����D��J�y�����V�k��!$J�غd���m�KhV�x:yz0�ȭ�}��<�S9�7�'��]�j�)ϓq��m@�mZ	�q
c}K�DC���+ځ�S���]���x%�ߩU���N�:������_Ü�g=;��UآzF�T�l�.!DrxI+��Z��Ƭ��ܦ�j���8S �k��d�BI��K�":C�q.sS�r-�Tt���d���?��,!M'�/��b9OL�s�T�oϾ���}���[�R��\i�	��/� i�|�?6)1l�"��י���X��k*���1����M�M�Nmc�5m9	�}i)ۺr��6��kul�N�g�o��ET��o�HZ$��B��\ h�}/�7{�5�t���N�����&|����������Ri�nۦ�{��	Kc+3��nz����u�p���4�s�D$�EQWO���u����8JV�m	�__W8�l��ȝ	v,���<��5���&�0=;�w��~O�=��T���*)7J�4����%��/+m�z2(�
���Ɏ�^�L	���'��#\)!>u����a�����AF�`�=3�0�]�����6�S��Љ��q� ��%/��*h�����x�.u[�s�#B�]��e��h�k.���V^g@8�
�L:�<���o�܅�\�8��j���,��`���ѱN�#�p��'v�jq\~�/�H�6��k-S,*!oY�Ͼ�e���6�]~�ݘ]���C�����w��[��n����z�U������=�I�Ў8���MKwSD��V�Ո�^ՑQ�v��T�w6�r���4�Sq��Ď�N�%7!�"A�������������aOA+Pa�|��@t�ّ>דDU�ò���U�aѫY�Tl͕��:.wu텫v��TŢY�Ɣ�K�.��kV ٴ�uT�I�k/ RƞC*U�/�>K�NR6!�Va�j)���鱏�&�ʒTÿ��[uK�`�o��N/�6��\6�o�7��:�T�'��j>s��C�����
��[mkt#k���|>eY�}�%.@�T(tb�4�8]�W�s�`,0sf���U}T��'"���h�.Ûe�ǐا�y�`a��t*�P�<�F���c��a�;	�1�a������Ѹ�5\j'^ Vc�*��=�O���p�m3���:�4q�����lS��C�\& �c�W�۸��~�S�<�Չ�h��6]o��3���E�
ωT�^�;pG�����m�l��hځ�:������A���ç�'?�bM,4%�6���8�o�W���%��ؽ0	覂&xQ[*�ҋC/��
]��e��7�M�8�&��h#����n����q2cOp���	^2H� $S�)�y��c>�0�������9)�����C~�y"^U����3�82Sq�f��]W�(�&5xh����:f���n��i-5�:9�U���Ěn������W�Ӆ��D��nI�xd��ha��w��c��\kI���O�pǶB��"Ch�����c@�j���U#V�P#h��~9RYj@tR��D���D��ͫ�O����2;MKq�6�� k��ͦ�T��p����7�ւ���~��xx<��yv��;��_Lj{�q���Y���6G�*x{�IY��8߭�ݑn)�ϻx6:r1 �6,��a��cwF��Uh�$��.������J�?4�����3�&XeK{�b������$��KfCk��S��8���������7���>O
ȓs��_�$��/�x��W�^����s�&^+sC�%w��U��Kي�
q�}kuz�޷"���qh1�**f�XGn���Y�V�P1��S�_����{;@�뛱���a���q��Հ}��8��L;1B���U�)����,��>1�������\�I��cd�PHs�WX��OsK8
|�!�b7ڧ��sȵ������w�����i�a9� ����PV4w�RYR.�J��Ο�};�r�e���Š�����ozD����٤��>ĩ�	Z5�vy��X��r7q����ʝ��I[LX�Jg@b:�
�W^Iԍ TH���Z�8&��O�X8��C7���Ģe��\m.�w�v~̈�8Pc���T_0��čH�F�A]Pj(PH�"���09;{�����E��[���>DΌH,&��cS���:ܵ�� OC�&qq�HZ\�/�nL�J[��Ҳ�4�3�O��ꩁe�r7�IP�"p�y�vy�ĵ��,��� S��%�_�3����ރ&�yM�<w�
����v	���}MЎ��G�6s��3��X��N�$�&7���B뗋@��㰛�+�O�C�n[J͛��q4��o���A�	�O�
���C�#BТt�3�8�1���٣9�~��K�m�:���C"q�FvZF���¡��竰��0�'���6�]��Ċg�N yW��9,�8��?�Bjv8�G�ڳ���EI;7�4&
˕��a�~���9�8y�۵�J�ɗ]F��FAR?%��B����:�ccyj���v�QJ=�F���.�jb\r0�|��D��>m.�$�o��I�\�܀�h��$��Y@i��VA�-ô�
�� u=!��a��Z7�^�U�H��MD�;u�4\�ڙΊ�ڰF`'-�v�����|��6�x)�|x���85b�oHb,2����&O�I�	�}��!R\&v��ʊ���'�*-�ڔ�S4�xR�l���cl�v�E�6��Oંf�M6�*�b����[l{���&oxS@�§��8���T(�[e1�b`�0'<@�G�H�ǘ���4���}�ٮ�k�m�}2�t\�m4�)w=2:�B� _;�uc��;Of,������<X� �|�@e�;Dh�!� �EEӜ�[1�KTh�7e:�8���m�1du�U�^�Z�:�+|��B���Y=�oHLj|�����;�`H�ˆ2	�!I�o nNb��O�FIn��U���!
��p����m�_�Kl�5�;���K�%^R\�Iu]�U��E[��d��(�|�-'�� ���H�~���c�����f&�Gv����������y�C�N�E�b��,�U�ƊSN�
�����
��wi@F���D9x��9^:�_D_rk�Ưn�~+30�ފ��Y�ÿ��E���1u�t�c�怴����t��xo��3Û`?g[f�G�$d��B�~�����G4i��D<��\e�(П(^�a|�:����b�@���I���+�6<U2C�n�W�S����I▟gq��DO���<t�����G�L��lw1�]�^���Vɲ*�3~��X���omP;�(�I�uK���Y7����ɰ<E�ϴ�C֔��4Ʊ(G�����N�^`b���.�y:PS��|����Ȃ�KQ�:��k�9�݉���~vBb���I��</g޷�BU��VA/�Y�z��ZUcƯ*��?�bD��\�'-y[jkE�0�o�t_�����S�L2����ç7%۸��h�/����oM���8	�L���C��g���歴�Iҗ`?"}/SJY����1i����Vc����>=����Ԙӥ��'��xRk꩑+FOw%�S����Yϐz�h�gǿ���0VJW��8����P�;ݦ��@��t������)����W�3}�����F�P�<��x�[�3w(~��hC�K;�pXF�HOi-�[�_L�O�������Yv�,���~
�x)�]>��l�����*�����g�D��B����.����������:�}���Z���S�/�Gw���?�=���ܪ�Yz�T����Nl�������S+�,�Ez]���>`F��8�E��W�źم�u��A
�gw����
tU���Ϊ�V���׀�����ն�>���7.P~H����Q����%��Bh�{�yZ`��������kaɺP�������}���S	#��,A��E=l!���(hXE@S<W��8���'�-�o�e�&s�տ�>�7a�ĉ�l���J�<	�H�?�k��#YvJ�&��7^f������GI���=�d7�7Ŭ�f���#�(�G�ƛ)d� �J��~�;��.D�@�dt��&ߧ������W�\�cd�."���fc%�,�쑐sY�P�_���b`ui}~�U��4"�xkJ8|1�(�M��֘@s{Y�	��=�vFǪ��o�^$���9^B(!�,9�7q��[2צ�1,.�U9��S��9�|�3NέQ	�'~T�\FJnR�!kH���q���c��C�rC�贶ԑR�X��T�k�E�H�gGd�o1��ϐ"�� h��7�x뀪��#	��Ƭ�I����?`���u�CMY4�����AM�x���\d��;�s(.V�w{�{L#�9B�Q&��v���'����@�����ky��x���f�pp��C�ԝ� ���$�x���٧�S��>����<=����G/X�xLO�.��(��QN��kd� ���aI�f�/�ӳ@�>�����>}ܜYi�P�q�4��d��!�Q0�M0���D,��L�2�ʊ��i
=Bve||�OYK@B��e���z�G�R'qJ"��A�ˡ1`;WZH��r� A��px>��tt��h0:�'��ԁ�&|��b�z�Oױ"%אR7ր��>܍�o�~~���JH��t�̄����D����?
�BK妑��4o䉼��<8[I�ËB1���p��l3�MbXϟ����f-}��,���.u����@���`�V�Ӕ�Ȃ'�&��?D\n�%|�'e ��#��|r�]<�lކ����U�?ܹ��nLd�C�p�NO�=�J H � �0���GVʙvc�޸�6/�p�s�������]'$��r��T��� �cx����b4�Ŏ;�;e��<JT(%h�I�r�z�T�/�џ٧�"Z��0��Ld���_���O
8��JE�p��o/}axL��V3D=������M#�fz�/�SqA�9أ�,L~���c17�ډ��`��̵�?m'ȓ�0E�#u1����#���|��O_i^,7�y�'�����E�GQ�h;zd�B �@g4�u9?+�ٶ3�Ua<�?�������ˣU�;~�:���_f�����6��l0-�U`��%�UTb
%D�ڢ����Z\��" ^���>BZ��L�AX��ߺ�Aw��i�L���7�_�P+��߫Q�� ��\pb@�A��k��ֶ+��H��i����LLj@���v#�csC�o�%��?,�N΢����F��QJ�����ˠ�fJE{
�[�E$���F
&�N'kN���㮓����ڡ�^�_�wǅ�+�"��Ry���>�����W�E7�E���6�Ur����<��Zؙ�>�d�VB�ʨ�ј1
�Y��qو��!�˩kxFsi���3
рd&����[�����|{��]_��X5�ȿ0�ō�)O#wiz3��>�v��@�3�Ƌ�����x�v~��RTi�rs��@������O����?k�̛�*� 6u���}��%I	fP�J݅ġ���Z����,}L�,��N�*��J�I���B�~%ѹ�R����./zeV���y
�D ���ׂ֬��L���M�u%��~CH^�M�-A�E �G���Y��