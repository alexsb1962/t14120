��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~��_&kQs�\�K�v-�h�$�'R��$m�J�ث+M	d�/ᘲ�r�6 �.�w7aᆺ�b����E^|)/J�IG�>�\�|͋Iѡں���~%����d��zj�b�Z��>)ax�6ia�Gi|Gq�-�B:��0_���/��`�w!�2k&/o-]�c�|.>��^ǔu�_��[�X��r=ad}��\�����~�.�򬡚�/,�|!b���,����%QF9������a�nH%�k�?��PxGYī�\��bd+�|ϗ87�����}�llo� |�x,�X䕄r��)������]*��z��7x����%؎�٫�Xc���L?�y�H�:��E)ݻ�Z�l;Mv3�0)�)�c���&L�L���F,ZZX�8�W����?&ks�4�
)�02���,�u�����Q�C��B��̤�Vx$�&�8�P�N�-����h$*�/;J� {����g����6g�	�������f# q��6+��Z�S�w;�Z#�Vi���=��H�)z:���NL��RLۀI�#�P��h�Q����ĥz-�Pj��"�/�B;����AT�v��A���������Hoc$'s;�5d��2����	���u_�X^�+NR�,VK�e0U"y�g���]S#��.J��7O�)�>t�r��x��%��Iӷ/S�F]���id�h�L@O�8N�~z�'��B?l�;qK�[>���)�&2#���+,�L���{>)C���Zȓ�;�d�sq0	c�	�/����,a�\Ĕw��̵���K%E@OM�Ȗ�����EɱT�L���S�	�S�Tp)C+}Z�R�����$�ֳ)X~/��΁3�jH��C����B-��,
�ű5�R�#�BV$���W���N���c�5Lw�pu�`�8���wUHM���Jo E�_��i%5��\�d����	4a
�u
��Y{J��'˛�{�.�%�)h=ﲻ�a�ڏ`�8�\��Z�����qb4�b0`����-Q1�0�V0QI�U�%s�b�ظ�U�%��U]��~��- ��~U�/X��9���Y�c��p�ȓA�&�*c��~̏F"���jJwJ5�]�$�u<6N�p�����x�4�yrK�=����S�D�,~A���Op���&E�`�7��d;Z?��f�g�ȡ�v���T̬��L�j�p3+G�1shB bI�?�����G��D���}��+4zI���5��`�^���thj^�C�^�oy����=�W"�Ɖ��Hʦc�N�H&��WZQR$}Y�p�D�U��/?�&�#x��b4X�n�u�����;bY�Ih�3ӑVuP��%�P2�}�<8�gTR���%$��B�'q9i� d=��M##*إ�R��E�O[S�,a� �Z�V�ʘ�H�^�*����#�̓�{\��n+���:�ė�?6�Z1~E�.�,gmx�j��S�G.���AH���)�p��o� D`�v��6�{Zu�����tQl��`�r��)2��Ԓ��$$w��y�ڛ*����@������6$�1(�`���O���V�K;��ة)	;}h�\~ �'uL�7��2ά�[q�k��������nz�Q��T�U�Kh�82�4�i�����@˪5?m�1�"ʨ�{'��0b� )g�S��qd�)�ɺ��Fђp}g��Um����=ak4���D4�S_����+ �L�Ԡw/^��Y�:/�bi)n	�Bd	�Ɏ���N�8w++��\u�ҽC�UԂn=�����h��̦�?)R�1���n~-�����)���~�1W�	ԇ��/�"�*10�� .R{�(=A�o��_x���gvh�_����?0���7�'I���9C
�Hs�d���c�G@�Ĥ��8���#I�<2r]rv��`���H��3�r.�����vl��'��@�fP��j�$������*�;:�sE��
Uv�*XA$CY�btx�-��ie��gw�Y���"|WlޖmF���OU��>����Y"2�'�L&�19r�0.�v�r��ŷˌ$W�F��h��38kUwC� �8�K�y���Dh;���0��Ŷ����r�X�I�	�g���2R.�4g��+�2;N�f��6=�b=H�S!�!�=�9�~�n�N���i~T}�+'��{��GSꝢ�q��Xs�(��� �Δ,%�6�������`����wY��&��i��;h�#�^���{���p԰�C���:��Z!�J��.��ZA�_���dq�وl�j�ˣ�#N�F%��LEt��V��e�r�(jm4ԵHAAy�){��_�ՙ%����j�$E�e�31BBD:S�����T/l>�!��m��[\b�������N��c+��x�����JI���#Gd����_e41����x�N�V�4�b8ʢ�\ y9[I��V<~�gF�&!��qO�G?ێK�_FҺ;����h�B�ܞ$�`]3ձSG3&p��rFvP�LX�LA-2qʬTeCM� q>���ѧ^ᵬ#'����!WZ�i�aT�̈́95�Il.�dbw�D����(��O=��J�zܟ��	�.��+*�������P�P��ܾx����*T�Jda����1�e]��(Y�Ј�a�Ѱz�f$l�p7��(h�����]diۄ����*)_H����_A�5�|����q��:�wEט?V�dvP�q��'ze�Ʊ�x�頞
�+�z��	�x_����&��7��1��B��U?K�'`���a��mX��ok����3Q%����y*�ק����c�T��M�+�`��[�K�s��Qt	��K��̾��!�=�l�Wꃴ+�L]KFLx�n�XZ��/Ʉ�?�w���]7���=�v2Wh�.���&&6y���O fx�ý.�������H ���n0��#c�1ZTe"5�S[�UE`���;��}�=^����f���!"i=?�W$2����=��2Zb�����|-W�ӮYb���Ȃ�ϩ��D)�K����*~��8�Y��q{�-�2�&t)�Nz�]�{H�\���ui;ƨ�;��^％H��Og��?��% f?�>>�I���#;��J6����;�opH������ŝ&�p�����g<H� 5���$K�<D�2��\��ޭI�E�HXq��\�����lab�r>j^u�[8O�kZ@��Hu)!�NW�tExI~ch��ུxʆ��z���rw�I����5z.����ل�-I3̑�V����{`�-Eض}X�6� u�Y��8!D�y������\������<�Yh^�����?\OpV�"�NQ�a+�]O�������3�/7���my|<�V��|�?x�����e	�k���->0�
b뇭���DE��Gz%h��U��Q��h ��S�4d��N̆���k~�Y�E,KScO������X��w�ޏ�{����Mz;��qM��*tW�wې���Y'�J�-�qat��-@���<��;zrЋ{G&�(�x��y=��$�b�{�x�z{�u���W�D���C����W-�R ���L��J,[����̋�����Șs	��z��;@(7�6n����G��-�ϙ>��]�c��f����w$T�5Vϭ�BS�EFJg�;9�mB��]��`s֔q���BVp ZP��N�E]�h��pɦ�iˆ����oG%[�f(�	�Í�u,���Q�2ʣ�, �e���u���N�Μ�U�r +Y�}�[��f6D�4�����8�T�n�K��*\�V���G��X�i��k �}��������z�D�Jic���PR�H��`)x�5	��SY j��=��n�x�%�UG�2F�2������p6��z+~i�t��meO9�~�c?���L^�OK��/��FFLar�a��et�J��O6����)�����wV��.Yߦc�_�G@��kwF+�wR�k����X֎�G��Y�a��?li@��am�1��8�74����̯�wMr�r������$h�ld����""o/� 6ױ�(|�'*�m�g�mz:� �*Xr_"@X�qRf�����a=�g����6�>�U���>�B��ݧ+��R�!�>�8?�90`��w��f���*��ŷ����O<�Vvo�S��t�/��1�̯�?M�r�j��g0O֬������<x��<=єo���L�ǝɡ�`�M**�n��.�R��7`���M��uu���0]�!���W^̗�Ty�����BB�|�5�_@�h%S��i	�T�:�)`�л�eN�`���uwq���%Y�7� �rO�t��1�`���E_	gG��Ct�ug��8P>ȴ��7fW�-5�̯]��hȳ���V����$
Y�t��i�d/ؘkA�s���d�F���;C����yL���X<���];$_1�|�#x~����DK��y������Fp������b��e_���AH.ԆxX�����r�Y�3<�8�;�T��5;��$-
G�J��0���`��]|��=oB�2��Ng�f2~�f���$��Am���Ғ�)l�x����.0=� /��4堤s�G1	g�<���J�ݚ��9j��o��*b'V��;j��W�sQE̳���H�E�� k��;(ށ6����<�آ��K=���Ath�~�=}N�0���m��&έs|�q�W�y0��S)���H�� �k�z���oi~���Ejm�u-x��m��ǆ^A�ml�ѕ��=��|x�O�|g^a f��ց+󯇩 g����A�vÕ�>9��"%_��Hh� ��҂���v���a]�A��Ҕ�L��4(`Æ��tRȶ_I4lS؜��;�ڐ����}��ICazoL�N@�P�U�#�"\�pi��dSn����ӨW�{��cE��@����NmUk�y��5��/
.'G7`�%r,�7Q�U��e�BҶD{����p!�y�h$������9m+M��|/z顋���[���7��'�[^�_��R	�wl���@5fPWC��_Ͼ���a��^���g�M�'�M�%��B����w����I"�)-q�y���`�h�:2�Ġ%[U��ǿ�갞Y�z��*{�y��.`�3�W���,IM5d1�V&^��p�4U8w��B��ZA�B��>W���LuQE�Ik,�&5���)L#LR���jz��q�8���*V��E��_%]����SA�z�oeD�hs�OZOȨ�J��ѱDY�c�K^ Ƣ����)^����JwA�q�������g��~�bG%r�/\�ʌ��O�YJ����*���!���n�w���E-4�ak�H��qF���g^y�<��p�Т���2ǭ#:��D�@��>œ�{�0s�]��3GG$��x�2�Z�FLH.w��#B�1$e�I�2Rj���<}]:�m:\�Qi�|2�L"{�߃� ��!��_zI��ۨ�BE]��^ռܔA�R�є��	!��\^��§GV�P
�0��əd���?�i�0�������`�+���M���5C�M�%����O�Ѷ-��x�ĒXv�4䢰�o�b�i>�b��C�J-�x��xB�>-|�:#uO��u}����ݏ=S�>��Ӯ��f!��<Pa�iNX�����T��M.���Z.����N��)N(Y}�L/,��X3zX�>��u!)'@i[l��ϟ��ƇȲM����}�T����p�I�M\
¢�߮�p~.9�e���?B:��{ǧ����yH�6|%�VY�$�I��B��:2A֦��g�a͐��<�2�幎Up\25��q�B0�]3Ԧ��M�e~K�{Z$�8����\��2��l�#0GR�ⶊ4����y��\�;c�+���;���WXbF)_�^x�4����O�K�3.Q�=���0%�%��W�Q�W:��%��J�i�����*G���A0���|�����CA*@�d�[VtjGǄ���{1��|M|���yp��C"��oͅ���4f�ùR�y���Z��yџ�������6�ZL�[K̜��)#�A���9.��e��ľZ��U����Y�(�V�+���WTCGk������{��;�t?��ￊ|d&�VWם~]g������;6e�]�����K�����ء�pb��!U�-a�fwD�?Y�v�;��ٕ�3�^�/�r�#H�3ĜȚ�	����HF<�0Pհa3@�#4�(��y��D.��:�-��������k 6�6�U�`����$L�?'����pA��|堋
�����q��۽[=	?p|��B����R�+��ג �Jop��U��m�|�dBp8�rRh�)�asld�4���$������Cy�uT|���N/�G�{F~�Q
r:�"�9�;�uI��Jz*쾙�<_L��sѤ�/!���h�D���Y�Q=[�ٓ���@B�2����Ԭ�ށq�)�r�[�WE`�K�T���`O_*��*0@I��30���]�g��*���9EН-�E�|M)Mwmsp$�$�u�:y�%��X�>�鶓��|p�t%�>����T�'b�_�޷�����ߡ��(CAx$�	��n��){�@�wQp�Z�ex��w��H��:A���!L�����D�A ��*	�$+�d�4�V<{K����eapO
��k3�Ƌ�2���K���V��Xw�<�����"��B�w�o2��GycPq�v������^:���@�2w�R�����Qn~�����e�O� ��N�ڴ��kYXp�p�֥BYX��4�C�����(�MS1� _�8G���(5�ɤ/B|��}�q�y�h&��0��ϗ�H����!�|e[]������uv�xe_�h��eoW`�'ڮ�ֿ�HOC�Ws+�\�m2��Z=�f��*�~���F/�*6�RI]=���2�����%��O.��+�Qz��Ⱥ+�
=�i�]����ʨ�ZC{����Pۘ�6hX)�r6C�lz�@��(���>}�.C���:����sӰ�S��"-|Џ�|l͈+X�-Ӻٳyat%dP(W4�IȔ�k8"�I�;K�&N,�cϫ��pV�s��Ȁ��{�ǉJ�m� ��k|� c�U<F^m�1���<�)���C4x\�f��|^�θ�~v�Yq����=>�����Z7A�gކ�j�W-|eMY�9�A�;G�J�ÿ��e5%ݑ	9!��Ch=T �{߽M%澎s�+�c��� �}�{��ߖ9��8&O9�*���Wb[��c��0�l�}
J����������K$R�ʮ���Y�xS����;.u|0�������U�ʄJ����6;/%�j�#֗�r/-�6L#�H�b�k�`�0P��U��ARz�]��Zؔ�c�0�ӋzO�>���'T� ���ͪ5���ف</Sx��L�>��E�o��q�QY��uS:��/,��S���iyBM�2Qd��h�c���+�H�����J�:D�5�B��ª�F=��u*I����0����t``̹��0xK9�#��x>$=��M+�2- pc�,����5��
*��%���[��������������"L�TZB
�[	��P(2��P��aA6��(-�����ܺ�	�Kٟ O����Y���OA���G��}�(d���,���1R�02q�Py�2��;W��S%�_�67��� �-3pHo|L�i�ɝ�m@��܂lW���5Hxg�V�n�Ľ���|����T.�����Ŷ>���R2�n�4]B������3��w��m�x��u(M� �E)�K��!`nS�]����n�Ƕ#�T���2�;���>��[�븷�\5�.h�V�ʶߓՕ�X����YC����g!��5��Ip��
�vz4{|"����s�!�rh`��/�RU�v�X�̾���+8ɻ8��s����K�K�|�� ٚHY�͗����Eۃx&�1���+z���L2F��u#���/m��|<_j��x�A�\�I݋vզ�*?����W�,�����eӾ�Z��}=y�⺾I���q��v�Q����q��PDT�~\250�f��?e����p[~��C���P��I5th�l��T���ow{�)*^
��O:��ju�NL@�K�"^�F�e�:�O f��'|���XYU8�>����@��J�~gT�=������!f��8�yԸ��䋏	�늦U��_y���'�VI>��BL����r�m�3�G4���=�a���� m�4���d}�#95��&ݯ���L�޸R�2Jh��L�V��X�_��u��|����/H�e�ټ�"��2��vmk8���T������l�v4s���IV��xcP���rN�!=����7��F��mqn�[�j3�94�NNVr�$��iNp<�4#/f���R�@���+6TL�����%E�	O9��/�#��<7�}����i��`�4�� �SI�#�Ot��PHn���P�����`ơ-���貽Қ�{]�J_��