��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~Q����<.x�ʁ��s���f6�eK?\e��۫6<uݫ��bYe���{�#���C��U+������0 �YP�~�/��x����-�H��$(�i��� ��=;W���sY^��Ǽ!�k���}��BӬ�o����5�����rBFk�ȣ��u?|UUC}����V"e�[�m�7�I�Pn)�D/B�̋j68@�	��7��<]W�c�o���J5���ۼ9A��V��n�H!C��k���+������=600���vR�@9�7�>��i��������r��r�6-�_^\Z�{���ե cִ�]P����(���s1��u�ٙb���H�����y�%�(10��^7Y겻`1%�����\w�n���*;�u17�1�N�/,+;2�cYO'e�µ�8	����#�����B�?ϾO05�gM�ѭhY���9	S͊�C�
�=W)e��>$���0nt8�R��ȴ�!;�I}���*EA%!���)n����+I�n�@k�����g<�n�8�TL�F:bT|����ĵ�����0d�9���F<ߨ%s�x�4��.��-�x�;��r��7��n���(���tZ]Gl�/�M2eT�.��p�%K��:���Y�ȭݩ<<�<����qn:�O\0"�j�<j/�@&�ͽr�G�y�;�h|	�1��o�\-�漫��\y�7��=1hG���9�W2�ܕ����[w�K.�oM���71��F|��L�I�����#Sq�@
D�r/Qu3��m��9���T��.��b�:�p_�8�"A@��k�გ���rV��mJ���v��bIņ�O�ڤ]Q�F���-(���7|��A&��o�9u�0t��K�X�q��^�Y69�]�Utf�<]n�0��q��{��n5���z���;�׭�Hz|���IN�����������;�rO�߁c���k����q.��ZFhFXYc�V�����mڟ�����~�a��դ��Q�L�󁾰u`��*�'ǘ�~?�
;�L�t�҅�H��ܶ����E���G_�|�6��eP=��[�o1P�S����B�=Ry6=	;�en��>�o���_��M���������}g�?�B�t�K�e��+��څ������H�����!B���X��`�����S=k� �N��E��	aᨙ�n�4�('e��?>��m	��:��6n�o��������³�����?Y�@uҢ������x�WZ�L\~������QMC���͠$�k��}�G�=����Í�u]������f
.	�T�j�fdW��%����VJ��J�V���e�z|�u��]��SVǊ���:5�8�J%��EYx���K��p(6FI`�k5rx���1m?�Ϟ%uDŨ1;�.�6���tf,��1~��.Xu��� a3�%�� ��&x�-��>��A�����>1��,��w�숖��H�7�yQn�����T��v����t����<���x35���/�aCŦk9��Zğ-a~!�82������]m�V������\������\]$�+�I�)��cS�����y��J�o��io`����F��5(U��a�Q\�u���t����aW�Vp5C�2`<�z���4Hq�2�B�k=�ȕ�ś��s��,!�B�{��r�B[x�q4y��?�G��u(�%.з��u�yЙyj(-�钤�2C�*���c^E��?���W��_Q��ވ���e�55�;|�#,G�T��D6]2J�J�23�/�gv'�tZ�9�pIQ� U3:{���[��5��k�K1p�8��0�N�Xv�۔Q{d�K�����G������J �6�9�VBO�ILV��4�t�^� �\��s�{����n��DP�����soF�eo�!��1D;�C�,:8
��,��.%��k��,P�ץ	�� ��e�ī"n�lK_P��WV���8��U��T��n����O���XY�5����ޖ��S���0	��������+�w@E_q�Uk��cf���ŽU�j�V�v�
�{��ݐTi�N�!�᫸w7�*���ۊ� 2{��L��S@�B���X�nE���А�I#�{U!U���`_�w-�BM6N����!�6�Q�;��U-�,�,!�3|�<s�+�e^>{�kh*�����.vd��FU�[g �ŕ8��-;��~��\{���Y��K(�7���8��H��;���&��tys��v�2ɕYR��@��e{QqZ�5f`ѯ�Z����*=!��� `N��@6�4ᵃ�2�,�{/�]RS�h�;56ꮐ���!�|��f����W&�A{	�3�Ǡ���y�����'���B�m�^�J&A�1�Z����+[4E��RSt��,�(x`�WD������bJ�%��3�E;w��Bf`���"l�9�z&
�k�U�� S�g�Lg��~s5Z	��8*U3r�-�%��;�˻B�谐��5;��4��uӞY�&����O�ͧ��h�W��v:ʵɵ�.� -|ұ*��LJ��f��׿��;���I���M�m�7���Bk���D���q֡�nP��ƙh��fs��ݜyș�)|�F�+��u�ph��f�A�ۭ�
RJ	W.J������ S��V�#K�뚢}7�3s�Me�/�@o������S��C-V��6�Rs��Z=vŞX��SA�*��&�$	q������l�m���s/g7k��5m�MZ,��lJׂ��0����Ֆ��ΈFNt�?������\G~c-1`����v}������
*����
��J��|���7Z���g��[���UђP�k~F��Q����&�If��6_x��^����Rt[Ug�u�����k�����O��:9/t͝5�$r�U�G�6��]��
�	t`-J�0k��:X��?��.�*���B���a\y����C�`�w4��@��� 8ݛ$y�D1��Vh2M�1_`�w�7su_��Ԟ��ӊ�]��<��l�q������KL�#Y�0���ʜѬ׽�/Ib[$o��y�Y��>D�6G������Q)�S�*MT�/@r*ߢ�Қu�XX�3�@����ܬ �;�رh��}�6��9���no0��jLz�S��4燗Ҭ��}��3G�U�B����$J��u_���/�v��/�)����]��
pX���g��`=�-���uS;���H�	^R��pﮂ�d<|j�W���g�=��<@ۮ^龿@��9��.ؕ��l`U�Q��k�x���p0�"�cW?�t�ᛤ=x~4�e��1���:zHѰ�;b_6�ͭ�U_U4��_j_6��l�*��^4��㟛�ԛgvʻ�Yn�b��R[۰�B�p�2��]ڕuʅ�U*w�a�EX��yy9���JɯC)�M����4��=�ӘC�Әyw���&�e�'j}B�� L�%`����~�զb��9�m����0���\I�e�R0��9|�NQ����y�a�ލ��)1�`]�K[�M��@b>�@�&�q������b����3M����i�4n��ЯQm[��b� �aW҆�V�����Ma0��r6��^�P@�U�c��ݐ�hܶ&���Vh'8�i�?2���܈b))��9�v4$�PS�a�ۍ��xR1ȼۙOL���N�;�
�ҹ�@U���i\�� ,�̀����o��+�y!Ƒ�1>mt�t�E�c��� ��z5�$F@�΀M�TO ����^����U�\nYՊ���X>i�/6���dE;�n׷�&��%	F��3�v آ7g��\n�8~=:{��~�,�y},6�e8H�����"O�t}�@��C@�� ���~fS;e�,>�q�3D�))(�1���#�	��7��0��\��[�B�ԧe6kQjfK�Re�qƚ��L�^w�>�����ĹH��!�MZj٥��4�g3��S���^�U]n-��W&��1T����1,�&���B7�Ѻ��ՠ�u�3j��b����P���J0~<��Tw���z,���ݒ\�����Z@��k�P�_�E)�3A��斥[��ʣe�	����F:����މ��S� !�W�P]���b�5CE
x�6����X�vV��OIU�ɶ?L@W���YFvJ��D;�]P�IcV����z�0G^4N��-�	BKs<<���H3 �O�l��sN[_W�uV��*F�nJ�j�l�8�o|�_�\��"Z���X|��ɈB�LG�씏�Sd��$�
i��o�ʕ�y��;ZٞL9O4�z��
5ziPa�i�$[{R)�o�]��}��8�?Q�U��X�2�R<�����V��t���e��Bʻ6��;�ɜ�u��2� �T���|�J0{�Ϙ��Veu,��	��/�v*SK��t�)cr)P����l�E9wD��k|";U��Ad�����쀧5��z�����	�Ά�T�c�md����P̈́iu#Nݨy��ȟ�*���R�m�/��T^Y��(h�q9]9�W�{��\�ٶNC�M)SI���c��k��>�<u�iYC�-�����ENW�������s}S8OXN�db����C��<�4��8���S���yt\ܞ����� ||�`�w%lb�/h���fQD|�r�H@��X�䀳T���p#�|N@��{}f�}���p��B��r���)tV�ƈ���`�&��8xIj)��^�Q�Z��~�u��vF�v!q�4����œ��'M��p�:d3������	7[�w"�ލ22J�Ѐ6����:������:)ט°�gE�%7}:l�'�L.Mג��x�
����^��Z�j�������B������%��MGm��L���m|�´��-�$�=��X{���b� 6HOZ��T���e��S_џ�P���m͆ӍK��,��.P�$�u7;��I��Q�9d�?I�0��O�I vc�l��;|�\|2�s����UM��������q�&�P�8+��!9p.�U��?�EU���ب�[\Bm5xF��pLk�	g�xt�ws,�����њ �4a\�{��)?aj��#?�:���OvO
�]@��s�q���ٻ�4ڙ(�<���;��J\3�OU�I۝{5��$2ǆ�G���?͜VL��� 8�~Q��[Z��0�V�ǚ��N�R+XV��S$*�����N���)l��c���|���S%���'����>�i��d��q���7	�c�-�X5��d�3�վ�ߢI�A(a8���1���v>���̊��j.={�?��k<��GY�y�<���� ��V󕕉\�C�Fw=�20w���(i�����&�6��i�r����4��P�Q����B�����G9��'�z��,�̙Yrn����C�o~U��/!;Jb�	����Nf�V�z;H.8���&r��eܒI���qV]��@�fp�⅝ty[��A�㸯]&D���Y�`�j��!F̵����Zc�����3�a�)�r�:K����N��3�i7Ě>"�PacE��
�-�Hbm��e!��&Cy�,���x-�,�������vo��`��
4ѤQ0ؠļ#`��vƑ�n�߃��)-X|�h a�n��ȠѲGs�W@B4�朞� �X��f�Ҏrv�ڢsH�����S?-��}t�'>%�PD�H�;}�7�ru�߭���hh�l6H�����0s�i�dJA�F�8��O���}��������!�}������}�ZS!�P�p�.��C�D'=����C���:v�;7�A��1��6���G�a��֨Rl��	����o��C��y�&O�$�!9m�@���z�T������lOZ��*��C$�u�P�q����T��ڧ=mE�q���%u m�G��l2���)e���A�zJ�ey��z�9Ij��`!�_�-�_Uy�����������pq$�p�%J����C���8d�x�.�d��m�����^�����B��y��]��!��Tv��7m|63��j!gm��{{�1V������
D�#W8���8!+x$���a�s����;Q�����S��nm!�q	'Z�8&1.L�: �����!gu���'�ڈT��2q}I��&4��5"0���J�~���㒍�x�QCB[������l"d,&�O��6�#C"SS�_2i{I���%��n�[�oNZ�K��4�A�-��?)�y3���p���d�R�k</�S����q��ٜ!�
�`L9# �X�Q�i+���3α�3���y�����(C���k{���Y)��`��x�ˑ$��-S�/g���tZ�����W��QP�Dw\���e3O)(��~�6S�9�W�*�\n쭒|qs?ߝ\-���w��Ud�W����m%��$��I�3ӌ�q�*i����ֹA��\N��U��꼡N{��e�"�|Ə���v*H��1�y��9iƁ��ʶ�RF�aLr|��<>���p�i�_�c�
��ژ�����ڊo�W��(V��1�A�#���6_�tƏ�K;+�H�M0ͩ�ip%NA� �Y`����JU��uL&�E��8��Ց�.�]	�@�
è�W��*��$j0�L�י��5"Ѽ>�r͇b���;�GY�R�#�-\�_�w��呝�,T��&%'�֓���P�e�y�v�}"o�,��n\����y�޴�O�����*����i^�����B{:�.�Y��P*�l�ׯՖ�t��lk/��FQ�ל˹ݵuC V"��{��R�������H@���a�.�;���/��-�D̎�)���S3� ��Ե
��(����*��^�C%\d�of=߷�\l�_N�8���~��F#��
����hI��EU�D��nh�AL܊W¦�\�5	K�/���^��`��7��T5k�]$߅�����v��$�����d��b���s�n�����;��kU P���%D8�0�!�E@Y��ԯ�.�AsQm��p�};�=����o�3�NA鈛���I���(������K��.1�o�FUh�g��ل~�.wX�+¼?���k6������\]���Ù@I(���mI0�q�҆ԇL�*a�"4Z |6��.��@�p��d��evY(T�B��mg��P��{!��t]?I`9�����\�[��C�̅�mֻͪ�L�Oح M��/2�����b��zi��E��2õ^�^���A<G�J�[ ��9\?��s�h��AMH"���ƴ���o��}<�%�+���;�Jx����)����5��||~���p5���߷r9 >�Ԏ�P�]&�s��|	N����eu�D2��|�|��"�i���������.(�S�OXVh�Ѳf=�t��JX͙� n@B�I6���	�T�b��m?���b�HC����V#��+Ig��+�J��+�)�8Vd�A��й�$n@?�*�D馔�����}��)��zc�s��c�h^����βq3sR?VB�7�P/B����RV(�&�9��d�4r�e�w��ta�VeuZD5oR��m�Ȥq_�^7�^fQ6:`D\B����3�cC��'���.��f�sM�;]��_3��,�R��ҶH�=�=���2c�"�k\���۩A �f��"n0]��:o2m�2��
S]�QҴ��#�`�;~r��*Z)���sJ7,�%d��]�J��A���q��K6��ma^�6�X�@��T$�����?I�`��;q��n�͂%���P]�m@=��.��"�_d'B�IYv<�O���#\k��7�]��Ҁ¯�r��9����@7Ч�V_l
������L��G��e�/.K�q��$V�H��w=�F��\����q�켍8H��1D`�/�K�BB��<:)�v���'��=�&��amƗ�g*�_�$Uv���e�"?��U�08�_��(M�	c��9x�����Fݙ:�O^���7ݙ�ܼ����Rs�R*	zh��N�q認:p��dQ�1;�k�R�֞�K��?�� M���|�*d0����S&�;��;�wW�a��_L��3�R��`|i@�����l�v�Sb�-Ӫ�x��+�[����4�Dy��E�<�����*�v(�k��ߦw�d�{A��:�h��q���@Ι�Da&\3�wd�O*����S��3�\���8�d��l�u�����Sk�P�>��ֳ���}�9���S��y�=H�ɇ�����pB��|%�0&B����!��1&��;~c9[P+����N�����!�"p	���h��R��G�Zj��&�+][�F�^��V��>�nG�7b�Z��O�ů�l��%�EG%��
�S6;�p�{$L��E˿H�?#.��ܻ�<�����A \�h�6I�.ҝFh�_��|vy��C�݅:�H�=�V}9d�w���X�ȏ����R�(��.Z[9�]$DX�N��t���ŉ\�$LXg�Z�Ϻa��K��q0��'��;�a��t쨰���e������{��99)�fJ�k=�32����̱��^*+�*��K��e���!2c�t����/@��D�/X�<7�=��u�\]0pD&�n���� J9��`���������q��d��}�Q޷�
u�����t�]�u�d�GԼ�!������h��%x`&K�孼V>�����u��:��U���)��ѿG��ٔ(��8�0`:�$6n0K�jB�f�.l�|�S��#�?5yE�E��/2y���Hc� �Y?׭��VaG�����>�9.��~�5SA-�*�iF�y?�qU��B����l&��Ny닢~t6��np�>r�+�zo����p���F��]ET�{�O�R�� =�ۂֻ���}�@&�C���Dޭ��w 6���]�z��5�(_I@��Nr衯��e�3�9�$n��9�f_JRo����K�,�Z�!\�癋z1W�.��6盫*����gPW6�%�ܷ����HLj��H��	�W�_b}��-�>|�l�}��_�/����
�朜�J��>�� <�zݝYn�:� ݑi<�FVuq�=y�b^�$|�u�H���H�%4��G�Zzd�F�A�k샱p�.��0'-<����_������|W����_��"J��SeΊ�:5]P�?�K5���S��f'�J�|��c^��aog��8��%��T����	V�Y�����3cb��d�U.K��`
��Z�r�xLP�����B��ч���iN��L*&����-8��dD��k�g,�Vm�,6��o�ʷH�5�V�%-�<2�UW�NM��{ ]�rmhL)lJU�f�X�V�/�a����! �wZ����&��2�T��m���$�@�%��vU�#�(��|l2� ��1���kt���B����CS�==C�`���AEϷy�q��F�ۈ��^��/v�z!���rP[=)��YP�>��{��v\�e�;dH���}2�t�<�Ne���$�o��K��sJf��H/b�B�	�B�]��2�ԢUD�0�r�rH���s����:.3v�N� ����-�j9<?&�waE�R.�v_�8��I�j�������m|ꁁ`15���D�Π��,�e���t:�S�1k"�;!uu"<m��)EҲ�������W����t
F�=L�����8�u��?�@VVxz�)��t>o1� EYA�U��y���h�,H�R++z	ki�&~�)�����q��	�㬚�n�q�ShF9�<��*��CƓ���D5&)��5y�,�[x�
�m2-��<W��u��V�f�_���x��wxz���E�qS�7���d��T�������7W1Vܹ��4¢�8�څ�j՝�#~D �����I���H������S$�i� a��o�R�{��r1&f%ܸ2xD����,#\�,趥�{\��97�]ӿPm�G�v��'dU����C������cFy�0p��6>�?6k�4^���#�e2=��sE�L��I�1��v��s/[�iH�r1h4&c�:=����[�,�����TX�Jz����X�l}��[I#9���'�/t�u��g��DV���T#��N����y��g�-��#9J�Y]vq�]@��#w�;�qz�7,!��2�����7�ԛ�|:�o���G���a��/�/Q��9��D���J�n(�]�ĭ�E6@A�I~�Y��[�3��FM&3O��������Wr�r�x}�X�vip�c:x�]/�W]�sͼWV �Їwu|N�����@'�|�{��s�dJ]c	l&����Y= ��)��Ze&�듢�)��r$B��'�Y'���,�����A��v��vl���sޮ��t�p��?�I��`��Ѕ�A��,LÒ�8�ғZ�w�փ����,Mtd�gӀ��;�fv� ���*��*��>� }�Գ$�p�ޓ���V�y�|�GG�ǋp7�T�D͎s}� ���B�C�L���! �:�I��q�Л�\����R��>���Kv3�'˛�������d^:\�˷|-�8�JcE�!�U+@��0J%��/�2c��P��Y�R��iJ��g���|�ɬ"%��Z��<�4�5��#��&�n�9�@���/�$��(ۧ���!ւ�S�2���eӰVo�6M�9�q���w���aJ���Yc�19��շ&�oV��Dk�$�S77��Nrj�p5��Yz�]d�0,V�`��%�'�_�_,�b�N�b$69�rQ�Z~A֛m�r�d���k��];,z��x�����gIԕ[D>��\C���A7n|(C��&��vɈ�����O��~���]�����g�G�.d(�,�1�حߌ�5J)���>_+����d#�
�9|���N�lG�&_��%|�*=0�``�O�*�_�cf=A����Y���s��c�,?^~t�e��T zWZ�&�&ǔ~*�p`�q���:�X,�ŗ���!Q�Tc$�b.��L�fX[n�6�X����V=R�#�����N`\�r*���W�'�Ej���S��`Kűs�f\wP�0|�_�������ly#6�h}����1�l�AׂM����a�{�3B��GJ�{K	�%&����a6���%{M�BG��%��HJ��z��������uθ�(FW�K�j�l�8BՔImc�'M�	��S����k����~��`�.5IU���,#9�E�Joѐ�M���{AD!$D��|��N�Ud�'��t��bVnX��� ���1dS��xQ��mWb����I2�c���q:�e�5��c�X��n=
�L��a�X�W/z`��Fv^�?�������'���p� &�J�jBy%���/*gCl~ӥ�?�$�GH�]�s��5�;ĨưA�H�x�H���Q��U��e�X�[D��׎�� �yU�#�[����(JH谲N�~=�9�
�#�p)�Rr��$BE�iBT�pv�C�����K&���R�e��WU?^xAO����'��qP�XjvR��HU��+�N���C�Θp�7��Ʉ��冺|��+��������n.>Ty3�^��a����D_ρ��Ť/^��>����L��";���B��ЈW����@�^RO����Lվ�J�O*�)�Vg��9�����F��[�9C���y��KXO����D�s�%����ld8��ae�O�	�,K����٧����!7Hl��
�|B���L��@�ԣ�����+H�՛�PG`/�=e���`V��Řcgz��^G�m͸�Z%� D��^|����?�5�o��%��ND�6?��8�Swr�����XX��(�:�B\}��j\�!�[�o�nT�G~��d�-IW߾H:�u8��*F��2Z*����d�\xk�!Fw$cm�䔷�&I���Φ��}6�0�ԒG�4)t�1�.���f��2b��~�傑l��E=��U�k���M����_�Q�9�A�4A=�?����G�E�Z�P�G*
�H��;y#�*�tHF����N&5n!�s��ϧ��Z:Ѽ+��eo���@pQ���_[O�r̚g��t�z않9�bH_����nJʨ1B:���CG����b��`��87�Kǅ�W�S�}�uc�Qi�=���\�)�R�Y�$�M��wd�:j���h�g�{�51N>�'�P<&{av��9�Z�~#�/cVJ��9�c�Ӳ�W���p��QI]*%g�n�^��{]��������6�}zd0��,Lpz�0X��l	��֕�P��4ΨeM�B	��MN���lUҸ� �e)���ց���|\�>ʇ���U�A�}~�����h���
�M+�)~���_�P�#��%��Z"�BS���P��{hP`�ʅ���ZU`����{���B�ō�3l	��tibi��硿�V������uԨ�@��1�����k�!&�B˹��1�Xs
�b?f"��G��
mfI�ӀT��Er#DֵK���!o���,���G��$�x7R!�L��Ǚ��D�:'��׳�C�����=U�=
{��0XWH��=^��YϤ�2�Ϳʽ���_<��E���f�ׇ�1�A�/����	���h �?��E|��$�|�m,�b��[��?�
����8�Ƽz�CKqk s2n^���kIr�IbZ'n7��U˝�e��'Z�-ã�
��+�ܗ��m]����C�8cGk&��ҷ�bp�0x
�g<JAa�$�����p�j.���KsBݮ6U5���/�A�3J�Ym,�a�(���n�U�iǲ[���ڔcR��Zgx ���,9��"�U� 	H!ٔ4B�i��GR���t�>җk}�9�<�g1�YMH��Wǫ���3Ң8��1��}�dLW;�E�~y�!Ĝ$�@7�ŭ�:1�bB&.4�9�yE��`���ѓl	�Lqz㉻Z�G<�aB�o_EK3/8�
�{����9 �K�
�\S5Z1���D�+s)L�q��L�o��d�������L�ǒQ.sDڲ���C�.�pU	�pP���&��ݝ��Y���/#�"B��tN��X9_O8��^*<����"�UJ��G*�
�Xq�Ɓ��lյ���P64����g숉'�\N��=�-+�q[�:(3�>M���� e��J�`LVT5�2::4i/;�JEY��"	�a�L뵢��S��3���E��`}�z�A�h����jCK���7e�2�@�(�Y!�l}���ȩ��4�	�3�[&'(��?���y0L"�,A����+�s�4�l^Q�.ЪK<[B�HPV�%BJU[���=��|��`fiԈB� �Oo�*���	��B¿�C1�����9��&.�v ���-�+����:�+&��'8��9-��8o�4e�8�R���i ��_7��W�1
�'&,5�X-�[�Fم�Y!�QΔ9��r�	��vN��� 8��М� ����ZAE6|�ym�qum� �\�L>Bfg�(u��ޠY�4F+r���<tP��pQ�gɨ��Qy��iYU�k�\��L㸬y���exHu'�/Ͼ��˼�Y�J�<S6˔�,}mW����<	�O�V����ٙ�7�xk�����8ר��X����i�v�Q�X��:h<.c�S�4��3��h�(��m�J��C@-��}�R ]m��z]��C���+Y�����ٟ&���/��<���fY:*�Ӻڝ��[[V�LE]�2i/��>P\��r�u�n��rRw|{Sd��(L(p�
y@P�U/�]���s����BE���R�Y�C,A���B�	�Z����?w�tj!�=�L�gr�S֙b�R����t��L;rR��YNw�y�3v�VL�n����'E��g��_��<g����q�.F٥߮}��>MTg�������;��C|ɮW�j�{���*���}l#|�n��`��"Z��ς�a��Z����^��/���ʖw�T-y<S�W�s�*�4>SF�4��^?�gj�O�$���GL�i��k�%��p��Ȳ" V�eƕ�QK�-ݻuQ���ERo����_'�a'��gT���#OA���M���s�#Nߤ�W�&�c|b��1b���u^�
Oz���5,*�<�_�k��Ln�RN�|�D-�f\K}����� �#%�`>�Ҿ�&50]��ӏ���R�������p���&6�}?�e���D5dl8h
-��Z�>,�{���A�=.L�ig���X2����<xڒJ�<����R���ff�������3%Y" ����ҹ�q3�d����SG/z̳��f�l�sG�p]�C�`���S�^ҳ��;=�w �� t+�3���5׃�4\h9��ɣ��y:������O��Q��Ǡ�i1(��(V(�ӌ�c���Hޖ��m���H����(ǣ۹S�#lOZ}�de��;U�U�c�:MÐ��@�.�	���hj�[�e'�D���[�`���Vw/�����7y+G'�.�H���]����-�)��lO���\�"l[�p�>?8{�VHR�,R�؅�$��Ik���>U�?�VT�F���*���a;��M��o�pA���"`�[��%��+п0b{Φl\ˎC Qs1D�@5��m���,������	��-79tt�+p+�O��_ٜN�`���*����I4�}����� ���ж����z �4~u��^�6�GZ:$+,cw�'���:��e�翛@H��)�ٷ�����J�y~���+&�PO�a�E'f��\�kð�d����AÍau�Aŀ��~��*���l�/���;�hK] ��ZW�fͿ����R˂����Ԯ���X�?.�JN��9܄�ن�� i�D&Ǔ%Z��яԋM�:\�. <xWJTr�!����<q����e7\�c}�
��w��>��������%��Θ�x�.�����/U@pը�^6 Z	����o��$^�@S�YeWk�d��g��֒����iR<Ϭ��\��������U�&/�i�"���X+u�9R�� ���B�7~�Wn!�jN;`Q#no���|�Wk*#T��.*	��@�F]�E,�qa�o�~D�!�G\|"�5_��Ձ'E��e:�4�_݆����z�"���d��_��ix}5�v �����k�-�|Q�aP*���҅i�]�\�t��겋�4xuc0���8�L*�?v�F@��g�?��{�\^�F�Z�����|%���r.�0k<�+�A��Te����b�be����˭� Kz6�rMm!�����0�f�D#GN&�8��-W[Hf��$��u�I��5�F���^v�:��ŉ/���-�#8���V� r�X��$9�u׵r�����8���!2��z����*B�m2��id4dl!���c]�S�|�)Xnj
V��j�ڪM�/A��]�_��(�H�1��	f�����|~K+q巚;s���u��z�D�̌U�3�}�1S�'�gx�U;)���6{���o�o�@Q�t�=UO��}I�;��(�?�~�ݚrMb�T�4�9@�iT�&u��f�H�Ӭ9LՔЏ�P�n�����3�gF��I4|��#,�\�.{Q>e%���d����V��#��n=�X�*p��M�ѠBd��T�F������h|c�ݻ�Ե>1QF�����%M��x�73�Oы2��O�6+������ �e��5&�F"�+/��'H�emZH ���̳QEͨ�``�-2͗T-Hb�>��D[�8��d3:�;i�푋4Q�9�� �q��\,�G�Dz3��������i&x�\ �g=��J{�?��'hi	�Q&>C=Uj�~�qDRg~e���dЧgh�cDx=r�S�Oi�à�L� ��Z<x O�Sup&g���AGH�"�X�@�@�h����@w��d�@�� sψ]u�Y�}�Bu����{�~kJ�ע���.O�K����n]�K�\�S��MW�t� ��"�1o��'���7DI��!�$�l}��Hh�L���b�k@�8��w�Vm��>�Sӂ����ґ���8�g*��׸�:�ĺe,�(r��K9(�����Y���:(Xhg��Uk>9D�F��5��;��D���Y8�Pv�q��bG��?�(�!=e��l���֬M��i~Cmt|[�rS�]�eh���Q��iM.$�p�,?��&Xk������s�j�B�a��V����0�ٷR���m_�����췑��]e>���_�I�A�7�t�R<��&�ps��#s4���+��/�U���C�H��С<�(bO]f`�m�K!m�gM\u}�,܉7Hn����|/��ԅ�y�x�-(��"�>ȫ`��7n�5_�1ؠ4%y|�K�N��.+`��K|(��<td�=�Y�񛝢@I�yQ����L)�t�	��J_�?SpQ4��w��v�}6���[���ܦ��ՅmC0��̈7�Wj�0E!ż�*�����0ڪ��+�%[?�n�!ښVQYΩ�)�OB�);�� 9�ꛒ/S$wW�?�2�o��Tl���~Yt1���ue=Y~�d�	�a�޵���6���g��6����P��gڬy�1՞8Ɓw������]��W!�
�V|�4����G�l/S�##���]�%	;[z%_E������f����]�z�u�ٕ#���I���K��QIF������
��T�x ��n�تgg�$/��,?q��Z�6�'�����#(�-YjL暶UP�A-4�4�G��+�6��8f�#�Z[Lf���ᢦH���%����ID{SK�7B��<���M�����+�IS�א=���.��5Pc����{8&s_��脁4�w�Է�<E�7��C�]<sZ�[!���}��^�܊�o�fL��zH	���"7��'p�x*��i˔�ً��#,��:z�Elb�&�%¯�L$�q��,�,�Bb8���p[��oCl���Ė�:����s ��n&�S	� X�bJ�SULT��1˟�	ɳ�^m'���zf��B����_�ѥ�k�T��k���]ǁdܿ�*WD���9��U�)J���NP��\,��'�f�G2]����I�_/�с�'p.�0O2�<�����*���E�XGAL�5S}��[4���(�H���O�8$|+h��1YM
������%U"1=��U^���T���P"]�mF#�x༫~n�hw�� �
%Ffrnc�B h�8�O3��������|��W��H�����y}�c����1� ��]�*g����(C�#��SN��qv )�+ܧϸޟIx���++�Pb�fz���U\�v[����L=�	ͥ�E#� �y�`3�p:s����|����i�*B��u�MUrG�^�Ԧ���6A��H�@'o��Jq|�x�%3$��}n��R
1sL��/��� \g�>'{�ܻO����L>� ��il�������K���S��`��ݴ�2ab,!.��駕�!�B�i�J<��9��}�؄��M�"�PI�ZoC#}�'X����|�/��XZ�hZE9p4|s*�q�pH:i1�t\mqicl��IR��;�Η�< ��K^�zv���K�Ԥ�8�z%�7�.��c�R��8���^f�|�d��W�`B,l
����䨥�@�5��R:,AK��rƈ�V�/�"Kd�!�ބ�Wg����
L��ic��&�o/<lٲIb���o�b�d���]��S��(�
Q�[��UD���4�;�M}��>в>K�F�/=�v#��'�S<���t4��zhh�I�Ɩe2�J���W3:������_EN�k,5De߯(C�%_�4\eu�W5 +��[vi��q�Ҋ���ߏ�n�RxQ�U�6�e����h�JA�
x7e������p��SP)���~���~Z�R铸�~�p��4�%RpF~�Y�;|�|�p�-U	o"���T����rcɒ���YRhSE}�]�	3�p-���6��W��ߋ� OO*b�囹�Hg�ʭ���qZv@	���ky���7�ۈ.�s��Y>ړ�4Vx�q˧�s��V��S�n����3Z��٭p�5ݽ_ʦ���b|:�v.n0w����!Y���R_Uk�>���������'��@o�I9��e�o�+:�s|d��*���7TT���@���/W�|�����t��䟜yͧ(exfpf8��U&�.G^YLRU B��ai1�hD��`�M$��;��l��bHU5��R%Gv�,�����1��I6�`�a5��gk��&�P�#�����sSFHW���vYZ}X)槫�V�Z=O�q��=�	��#;�s#je@�RK&��J<��;��x�Zs�v���$FN�+]E\VrBς����(r��[.
�2��!~Hv��h{�;�FVv*L�X���ݲtl+�_?G�W/EJ� �µ��fU�S��|�2?�D(��}�fw @#�^�vG��%HY/%�ۆ��M�Ѳ��.�i����x��(��!XW`0ˉ����+k!GT�9���������������\�]8�]�Ʃ_Yj!�_���@�����}`�p�V9��eؾ�Of�5`�7
b�
]ƦO94�q�t�9d����M����)m�<�M�	��Ͻ�����u��4$Md7��YNM��y�6��C�pA���a��t[������#  $���,��{�.[�k�VP��GnȞ��x��y<euB"ueR=�$�����2�9ǌB�,39�t7_T�
�T���>S�\���5U]\�
^ț�-��	=�4S��f��H��#eӢ���O\z���"`��~Oy������W�� m���q�ٵ��s����K��ΔV�̦����	�z��)'\Їc�d�>���-�q�������e�B�1`3�Y�rD�-f������	�`���r���TB�~�Ȕke$�K0�3�|؏�8�o���d`:�]F�c�QYLq����`(lOB��3���#m*ҧʺ
0�U2H"+n�	��Y�Az�Y,段�
 �ۆ����E҄��Wh��6A�_�`'"O��BVS��~���"���pF�x#]s��j���	��4xɅ�^�\�@�7���v�B������ot~�*�g��ށOC&󝃴^h�ī!�| f���(�Y˻(k����+v�ǾƸn�7�jhe��j�b
�}��Px
~�-#Z����*�D�N3	��IߐZĶ�/Q�����:�Eض1���N�9ބ�������r˩VD�
�d�oJ����$kڱ�+C����,y:���������DogA��Uw��)p��l�T���n�5E���kH�-Մ�!��2�.`�7�ۻ;�.��
~�����l[�	6yJUd�)��b_��blQ����5{T��N��	s.���=���!@�ɖIu$�Cd�x��I�ޕ,1wC4{e����G�o�*Y8��*>0+%��|�c�[eY�����5U��S]�UA�g��V�k�+���b�!8d'́�{��=��h��=���R�9�4��E��oՂڞ�y�H|��u���`]6N4�#
S����\�U��,���l���
][���Jp��w}�S;{Թ��,u��r
�BA�~o�(�ɭ��ɓ�f�)j��������.N?�W?J���;Cp\���6��˶n������,<Hq3l´�����D��Hlm�%Lu �-���ݶᯓ����l��TmG������دmij|f�EF�.�]���6�O,.@��\��ё���r4��/��*w�%i����J���*hx�66��#��ٿ�*$Y��	�	̖���{����� <�Gl��*�Yf�s�z����ck윘ҙ�2i9�o�Z��o\�߉m�6��<��G��k��>m�8S��4��K�?3g	�i,qC(�)l���ž�A��7�E%m�)��釳U���������gz�*�M�Z�E��d�%��GLZPA����yD�d�#��Ïk�i��� d�b���h�)_U�rKv�+�GLE)��4����7�N�z�f�1�R1+xam���6��ˬJ�1������BIǅfZ�֣����3�����z�94�;��������v+�h̟"�VX!��B��W!���]3����_X�x>{�.��j�O=p���������ҋ~����U�7i��8�����3W���a1ud���4$����%��p�Z�͂�Rw]\#b!ѱ�\�)f��lٝ���_�k�}.C�4b���^���6f6z���zxzwF#���}ߏ����/���B,V&kd��ux?j�J��Ъ�nGm�{��<�zQ��Qe�L���L��\�+�(���f�tf��`�����d�5��&YEb��I��}��4��T�Wa����E-=��U~�y�:�/�r�	�uWa�|N��<����v�V�"��|�������ST:���А��e�S�Z��C�t����Р*eGS���, ��)Y�fA<�z2�ŝm�'�#��NI�H`1�aw�����#Akլ�	\�V�j��/�(�;}�) ���E��^�����Au���?�n�-L� ���>�NN�"�E��]ً)���4���zɩ\m#�o,�tD06�֪��9Ǫ��fJ*g�傥�	�V��ǫ�_+�j���Xl]L���<�|�l<��-�*�x�ٽ����E8�0oE"�e,GoZ�����f'�ZuD|b��̭5�[�h���fk9���-���"����￟f��
<��A�R�U1B�`ijd��jT��-K@N�K��ٶO�P����4^��5MK�I��k`�d��j��^i�;��ŒJ� �C��%9��G#A�\U��̞�آ�d��$m-b�̑D&Y�Z��՛ffk�\���4I��iF�4Q��4��l�}�~D1��� f3�My�x�>��(���ѹ�ʠ�)E�6��`�l;�i��DN1T�PPspS�y�ʻA<*4�,���P`�9e���H�a�KҴΌ��7��X�q��ح����,�@ѧ�{
Blʗ�[mc��}�m�л`�rq��Ĺo>=z�j8��=�՛44$�4u�����ƣ�_b{�"��g��)o��`��Z`���	�UWj\���<o=�i��:�zu_��=� �����u�Ȗ��{~�B�!�(�8W�ڃ�77����~�QhҶ@×�U��hԣ�a�_�s�h���M;uO�~���CI�Q�`'��#�U=34{W|k�x׶�̆ɉ�V=�'�Hj�5��(:�q��_��I1D7� �S\�:aڋ	���?���p��]��(_:8S�o�5�И�.�w!L�9*W�Q&@��-V��khTl_�1��id̔�9�B��(�������V��ϡ��KY�&� �B���fFz��{xt��M_X��s%�ލ��=�t
6b��VpT~ƟomAq�\���Ӱ
2r���^�<�n���Zd��v��-��� �ܼݵҠ�m�mRvc�6�e���0���]|��S`c<a7��L��������ɠ��Ȃ�Nn$���	�BO-8��˳Y��4y���Uͻ���C�4b�Ύ�������
��p*����R��m$Ck]����q;u�9{?��ߺ\�K=�h�QA$��,T?�1�we��MNC�&�]�??�_$�~#jw�?G�A1��W��DꔸֱN�Il���U�+�����}CI��&3i��|7L�8���[�	C�c�t=/�L�[���j����u+�P�.^bY�ڃR�ғ��!�:ᗉI�~����yӚ�WD�(��ߗ�Y����c�[�v³�z
8�0�_a���ʹ��_V���o9����Ov`��/ �����Cu����SriT���k����Pc����9�IK&4��s�Mf��z�HY�j���jrܮ���N�!a��iv\ J��V�B��w�����Ki����^�^���e�����़ː��椤�"u$�t@)��mw���J6P*�~��y�[�S����Ҥ44�d��ہ�`�`��: CP�]����Ӻj�*��;qFbؐ���$���1����($ƥ��Xl���-!�K�t��� ��z��+C--���'a?DPǢ�4]s{�\I��D�M<�n�.��H�s��@�~�' {�<���ϙ��}�E+� |�Z��� �Ky���z�Ģ���^�'�B<<�u�LHsf�.-ܑ�4Z4�I���o�ڕ�Z���Po�jj�Wv�b�i�(�d�J랎#2>�|��d$p_�7�5'O�+!�1^�� ]�!�U���Ŧr�t�J��
f':v��`8��`��p��8���!ڥXS>����\���@����?�x����oV���q�<ZR�\�P��2S��P������F3�h���׌��/I7���17�1;xy����yZ����o����Z޼���Y5����@i����Pg�b5�'~�Qp���9�^��ZIsQ���/S�4?�����q{����2��nx��#j��p@1�i�)��MEe:Q��hF��<�9*��O�P��
�.J�f5�q���0��	I+�)��*!��2ڂ��h9�Ė�K�7���/��:H5�|G�ow��14����|��=ؤ��s\��7	О�&ln�IQe�4c�'��\���.O:r��%吳tǾ�	'�'h���psE��;@�/Pk㓬�8��Rɒ����݈�O���Ϩ���)ЖX]�fдkK� �z��Gg�����د�H�Y���Y�=�a �Wm�GX��S���^��w�>��υ:<
�6��p�����)FP'��� �P��K���P>�0�1��V��m�7@�����!�Jw��6餪����L�\r��:�q�1v�`v�U�[�Ā��Z}>T`CL�5{Kq���u���3��
t�F�yo�bj�{cw����"Cۉ���c3���H{�����<���7�P�f*�$c8Y�{��xQ�;2���W�M��~�D�=���8�Wi�5�v���"�椯>���1��	8w��>#�YA �4f_釘�I����ES��J�b��|J<�[ ��^�
J{�g�{�%-�V	:�)+�3i���Z\�a}B���aED|h�]�w�~�P�l�:���n�>���Ī���u ��Ǜ�MNp�;d�z���N3�ި�oEE��:�������� k��)�Ay��z�y����l2.�s̝{.o$�Ɵ-t�Ӿ�m�6%�T,+ 5?E�����y	E��{��1>'���d�y�xڔ�~O�tIz�\��?��C�������Ҍ����҆��;���GJ�o��[�����1���<�<�H�Y��^t,cI4铀�4M��kG� �����n��N*Ӣ�3�o�B< �:11���v��ȩӧL�G��@e�d
'?�ps/�ه��m�{R�\9�ߔ���6��[��@����=�x����利��f7KĖk�K�$)�K���;&1X%β��q�����;�����v�S��Q�Ѷi��L%������) ��<��(����l���9A�a�U&��m6n��o'��+��B�x�d/�gU�#^��� g�;�"B�azo�wY��`.t�mJ��yw<����cn(�m�@�s����ߊ�g��:.�ٞ-���Z%[r�V�lx��٫�U���1�,���J�bӔ�l.kb��N��5ٜ�y\���[� ъ!d����d���t*�!�%{0�Py���/��5�6l�\~�$���0��a�\�NN�D�j���	E���s�<SdNn��闋�\}�'��W�n:���@S��ߙ۶�@�7�AT�{/�W���Ч@�SжDĐq���-��ȝgXג�2���~��;96�G�<�F�E�>�<�+q�}��@�.�"�9��|�Z4��@k������v
����;D��j�'>�g��B�h�'����d�2Y�4��i��V�y\��'/U����Z�g��e܆�Gn%]��%�߅��h%l����&�t@i�%dl;������z�.�K��{<۲�K5,�ʕ�ˡ����~�e�"�v󑔩�~�̾�$;����$�Y�}Y6 �Ivs!@Q�*BL����K� ?8�����"��(��dJ��q��1*B�}�vCiN���r�cN�RT1n�!���.�t��&��蹿z����4���=�p),,X��,�4,��m�p�:��I�z���DEK�q��Aq�n~_�0ٝ%�pv�^����PS�j.��z�
|?� ;+��c�!������<�^]�ĕ���-x֞Ѓ�����
M׫Ե��Es>�L}�]��zc �1a��d�󲯬&��E(���5���h΅Ct����}�6��TQ\�M����՜w�4��T�_��H���O�V	׶4�D�r�*�B�OW��6շ�+�,�:�WT�յ��/UP]�^��随s�+�'�+G�._���a�K���ݺ���"��;��#���Y� Wi!�HjP�i�rG�%��K�$��S��~9dѧ��]N��;`L�.���
d��� �@����� Bx��C�j��ã��B�jS��F��}��ʰ�"��9R��$Mo�@��$�8�� MIH�K7�<u�4�9��y������%�M@(T*��,��$���E��W�r󣺪CO����-4�OW��$���7靿���5�SU#���k�Z6���y�m�7�Dэ���{��7#nٌ��d��^\N�Z����z��r�Ck��
 ���v��#76 ��KG̪Ÿd",� 	R������h� ���)��:�q|^ٖ��gv�-��P�c��B�?�h�m�����z� ��i�h���+KSL��5���j?y�t�Rh#�w��TQ�� l����s-1�x^	�K�Y~���Q�ϯi\�F���v	���%�X���W^�����x��u4��z�yx���������) �����n�S^Q�ep G"%�B,�!��W�+������I�K��*���L ܽ��<�a�i�`�k�����q��=��w̓��S���'�%�߰�[�>���iѶs�,�M��- ot��?-	����T^s6?}Fjk��TSG�|T���FX��V�5�\$S�|	��I�{��[Ύ���-�߉�Z�8c����*����қ�d�W��O��^+�ba�ȑ�N��/��~�,.UL����QnQ�'����L��0<��V�������܏�ԑ���'Pg?*,dlh���$ �w���	"L��T����2���d�!o��� �J�=ָkpkgz��Zc�>FƔ��%D�;�^�st�Y$���T�Y��J �h����+��Z��B^W㌔��Ǒ
�|T!H|�y�J�e��,��/� ���X�B����ߤ9� �F|�k<4����%Z+��!޿_^2�����nk�]ӴX�����?kO�5����heZ!�XgJsX
��L�qo{%��+{��iC��[�\|�62���?j�:��o�7tԯjc�����d;Nc=��ÿDwF�g�z���9%��U����O��x$jo�ZSw��S�$R�ˮ�.�����!��u�b�x�;Z�{h:��E�^}MGv)��V�9qڏ��Z�[<�Җ��L��F&�n���Is9p�^X4�7?k!ӈ�ل�@ ]ٽ+���?K�>V���j{eLk �G��v4��&*T=��Z=;�@Z�޺p���������p��`H��vo����3�Q�ǡ&@%�p��!�vщ�g�x
K�
������7fG�L冧o������6�?8:d�E.�%G�~n���s�����e*̢b�̣DT�1!T����&^��T=�}<2���x�� 7Ԍ{�0�6�I#r��M}�!ܠy >�6�f>+7lZ�Ӆ3�I�bϐ�c5N9��KJ���dr��"i3�z>���p��<�2{#O��lr/�bv�>���*P*a����F����ea����ї�Jl�����bY�6�#u�@xR�.e�-���}Em�i�V�#�;�B���7u�lɶ�#C��%>����1�#�QY<%��q�K���W��‛�A�B�J���u��p��|IT�ŷ�_KN�B�Q�D��*i�ԝ�K�u�;�}.�V�X�yv����9����b\�A|u�i�j��"��z`�CR�ۈ��~`E���1
��?��B����ݕZ��R�)������q?ԗY��o�Qj����������QAL	�g����N�Us�䪷57Td�9id��1R�`�LT������(b	k�O���C�}R5Ҵ���Y�Xs?�e�^mS�T�Z5��0
�XW $no�����Z�P6�zmQv��Q����p�����{���C��GWR�K�j�A��ƛ"�M�FP�P��b�f ��ʉ�żh���j��n�FJ+Āb�N (�C�+�0q�R�o$��u@�#P�6d�)z~	�1��K�&M��=ݨ�]�.���:R�s���p��=��é;*�_���5P�;cZ��9^Lݏ��3.u�Ē���?�2�~��m@��7���$v�i�.�8��q`�o�?9J�� ?�����Y��[�Q=� ���Lw}��w�F�{�>ܣ�
[ ���|%H��}���5Z0���8�� >���<���ڡ0�6������{�L��o�r\�?�A�J�;����ծ�3�6/�c��+��]�4C��@i,�mϣ����#��2q�9����'�![�˳L��6�Qrs���J���=E6�1
�MjnQmZ?y|��x[��x�=��G��.v5j��[h�
t��q���&D\疰�@1zH�>��
"��n�I�3�k�����X�jPU�4���Fʾ]�ˍ��5�e0�cE*����U��r���|�7?��ϧ����x%R�1�|p��Bz>��e��v�� Xǈ�'՟q�,w�sǀ��Q�Mbҍ�\�\�j�F@˫����.$��l��Z��%��:i�Z�.$��p�ۅ����Q�(���B�Ӛ@���do*�����97�P�e\ʦU�\�j �6n��t>1�\��Ċ%:Tk�?��qr󓌖�ػJ��-I;S��Y���*O���m��f�p�ޗL\�f	wC�CkB'\����c#y�5����a���uN�2ʄn�.5�&fYV�@%�M4Y�C?�w�J`K �i��q��:�8����*Ի������~��@�z�#L������DOr�]VZ��m�rlW~L�kx��JH���T���m�љj	%����D�s��@{QQ�T�U:�{TW���j���d��D�yRQ�+�ف��X�C%�9E�2e[�����(���ھ�����c!��{]:��R�����)�����A
��V�P M��*�e�ؓ�-_뗓�W#)�=��T͑V�=CeW����0K���wE�/!��[���M���� �nUQ������f��81c�����+���>;_Y����G~C[����ӱ��x���!�ˣ���������a��_��Ҏ�#q��)��:ȵj{F���rL;��7.%`�Lr�	����aɐ��ʶ<@�!�����lzϿ߷U�CC�^`�i�Rr;)�><�R�tEƦ�J�IT�9^?y�ؚ��l`��"��/R�^A����L�������ɿxcV��#c�a�ͤ��l'1hd���;�B��]̵pA���8
r��w(�B{!�{uY��5�l)���d2\�>yغsK���� {$Q�v<:U�M�9бo�1#�R�r ?�Ə�A�~��^[þ��=�O/0�άX�~Ov.O�*�}�t�Ej���˧�kS�4K
|�%�)ܶ~�pv���\�B9}$ܯ�A�{G�%Y\
��:|��7/50?�=�M��u�ʰ�QI�����1���Y���P�g�(�ra�S~���"�~��O�w�_����:uA�.mΰH��$�~�o�:��#�+�*QZ�;��E���R�Dl��52�6���[=W.v��֣��rwR�;^���a�����R�.Q�Â�x8qɊ)��#�ɱ��v��O��5''�kΉ�O���Iw�I�|���I~h\�`1�����}l <��nW�B�f�(3O�)��k��E0?�a�xOG���]�;��C�����h�%�k�TK:R4����f�u�[�I���9ܥ��^�J�B�~-�m��|���9a\ �y�GJ�$�7�6g�R��DmԘ�W-����X�d��E�j�y_z���G2�]}����#5H�t��v��]۝C,A4F)���Q!f_A���{�}
����9�5�"���5H����m8*ޚE�w"����wy2)r*��S���WZ�/��(H�*7����r`��j{�ôk׌��Мv�گnQ'_~��;��=v��LD�����70 �0�X̪����e��A�k<�����asᦜ��:n�p	m׳����Q#s"�Ј�Rn�� �ӫ��0�'ۈJ<��`�¤�c�	������V;�j�M�������f�;��j�O����lfd�o�5��:�tIH��'��W��E�P�K�b�����Jp�GQ 1����m�uW�H�,�(~~E�l��t>0��#��ؓ�� Л��錁��	\K W\,p Pj��zoS
�a�����ѽ0hv���S���k&�,�+ژ~���͝���XTϟ�qR���n�P8�I
΀��pO���d4pt�̍$u�ό��֐@�����R���ߝi=��\�Bf�{K8U-A�g&���P)pe-�v��))�f��O�����+~�����b���_a�@B8R�!��fw4��O������[�I��BQ,�νIEsf�i*{2Uf�F!K�f���6S�n`·�p'e1�b��K�Z��K��`�ˣ���,��rF��2�H8G��dsaH=�Ki�>T��Er���t��̇UX�T�j����7��Pߦߞ:J�t�x�B�ʀ
��8P$��hn*�=�c��2�����s!P��N����w�!��bUw�s���O����O���m�Յ:�1�.Rb7�R�RWIK��n�~��Y#�kxdyO�xޚ�B��D�g2�NmܛM��	�Q�J�i���kɸ�����6���x፹�l8��D^�©��{��z�h�!����6�T�^,Y��X`�v��&�nkk��$"��L�?Qly`㐽^}U%���2�|3��R������r�w���Je�AWw�G�{�.����f�^�yʋ�>^O�fm<�ܨ"s/�k��Z�B�����
��rS"�P�*�?/y���R:0�R��3U�2 ��a�q��TK8�(����x+u��#h3xJq֓ Jƹ�uU��n{y�a����F��~���N֕�o!w&��@G=��p�E{��Xox[�85r�ڷ���@~Z=z,���&�,r;��t �"�Ȩ�W��n�j�{�|TY�������z�JC���,�Z.��р�>����n�랳L��%�z��#:���Y#(r@.��(<[��ƷCc"���q �9��o�`���e��?� w�YR��H�_Q��˜�Uۜ��v$.r�p%������>Y�^��Q)���b�?ƾ�ZW��'c���a�dH��n������dR�@=o�9�PB��ף���,�_�$�l�5� ���S��{>�l�t��f�-mX�i�.X���n%�.M��J�}Z�1��P��_�_\˹˳wD�O�34vo�:�L�l�&\�/o��P��8�^�݇r��޶$�%���9��f��Ħ�9D'�)�hA_<��p����cj$������&�.������o���F���քV-Y�U1��#��'MbP'T��=�F�=�B�|u�;�#���������1��ך=h��!a��7��.��Llc�!�w�&j�=�6�LgFǲt_h84�0�I`�эP�a������9�kN~�Ihߕ���0sb���&�Y�?B�C�)����F�-�z��3��c�x}���Y7V[��(w����>iy��,<�	��%���lC�H[�H\m�dO� �K�g�D��j��H��^E�㽦ѫGTJ̕�겔����Zk_ex�`ғC�9��~m�*T-��CfǑ��ת����3��{zId��w�n%�x�1���$�kH�������@n�/0����mb���N����M�� ��ۙ��c��9id��F�z ��BO��8���f���~3����%_6N`2c�3����|0AU��e Aћ�H�5�ȉ�>�u�eFƑ�w��T�z\1�d���8���85Tu�5Y ���<���eK�+���@��Lj�a�9�0a���<�1X�q��{����P��[A����6���^s��[�B�]z��fN!�ЪS�u?-r�������q�Kq|���z��nЈJ>�#��;��B�Cmop!qf��pو�����*�,�8N ,WU(�A��a[��hz�y�9J�Z
��]b�B�9Y�s�%�;��-�e[��m��*�(�"8L����i3E�<�wN]q��J�ܞ���� L�=q�a?������k�Jm1���ȼ�1�X�í�ü�{����[e+��kJ�MԼI���s��J��G�+�Y�N�&�WT��dS�lqA��k{-/@��e�_^rv7��xN���ԯUS��v��D��D�����u�K����K���K@#���t���J6)hՙD ����R�1<Z�f�@�j*�r�l:ؤ�������?�w`��3/p�D�����E�@�=N�8#@'_r%�!g���cu��y�b��ݛ�����u�sq�a���\e�f�[2���C�H�� �2h�f�J/C
<�sָ9xTf+H��"�'��*w���i�OG�ݒT,#���*�$�-R�T7)���D?�)����X���<ƌ�/�Q�~!q���όY��r�X[MIGEաV�,�u���6R����b_�`�Y97X�x�#ʒ�+Z��Y�d��*~O��s�J(��TN.� q��U���
f�v���>�]��H��|��[�|���b���E���D���?p@�b���i4�/�T=��-�V42۔x&�O���
"�f��#�&{��og���tn��z�Dw��ʫ�Q=��G�ģ_NM$dU�T���Y]��N��ͷ~wC)+fؿyX��?`Fк�.�y^��3�:5�&D�kX�R�ən�d��Ē���|:��~��愅K( t�JBq��{o,�P�m�A}ln���<��z
��>�Mm^_���E�l����ܥ�)�*���{�p��br�C�f3�O}5�xɔ���1�9��k }ae"m�l�6����%2���.�!,{�"؝�S��}�H��{�V�E��6��ݐ}���C�%�c6�f��������R���G� ��u�����i6.�X�d- 	I�������Y�I��?�K�5M�������
9�[z֧⼥��Y���]();}����!� Yr$7	i4�m�K���}�{��bU�®J��~�����~6e\b��%	�B��:�W���G�7���ͳ��YԺi	F���z>*�
z���B�' �lkKec�$C�(��[��`QP�S�DϜqֹC��g�:�	�mD�Th$�!�%Z�pz]fhӸP�f_<�AY����� �9k�$���΂� _�Rx��mZp�����:��N�+P(��ub^=A;=mM��C�s�{�������U�<����1�pǀU��<�n��H�;��j�pZ�o�ARM*�y&J؜1<�Ȧ�:�R�䲫hVѬ���V}%�%f�V6���5��{U7���W��=x�qIwm��A1�!w)�c��."F��X�-�`���K�78po�G;�ݝ��R&ޢ��;���q0�h�Q���M�����Jo�k�c��~��0A����7�曕����⯬��Qx�t>���-�˞7� "�(4�6,rv:�ݤl�Pot0�+�/f=]�^T9���nȅ�w�_���,��ݤm �{��u��ٮ����>��>}+k��f���½�5ynˆ�	T��%��]͜V�=��2�n"Å�l��j���AAH�o:1����-5�3$4�ظ=� �oZ����ʅ���LX�s��h��CTNI/��b8{�BuU0`x]�ɔ:�����h�pDAj�G�:�U�H�"k�N7jS�I�?|���U>�+
��/6��4̆�O-܀�:<P�z�&$q=ք�.�L�b?�v�,C�6@ֶ�ƛXou]��e�I������s��Ym�]'��:h�3�棘��+!	�ǁ<�����L���
�@:����O�Х��6�7����gc������J�l6pE�����2��$ ��P����Q����mڏ�hDm�]s|'����2�_�x� �Nrb����D�,"P��e=�ۄ���}#�'l$�o��X�<�n�#��Jp��,�N��IF��;�ϗ3�^�	����#�88�尦��,q� �Ѥ�Ǻo1�yZ
�����ED_
�>��!9L7��?��κ����=��nMXD�g�e� c����;6�^�-}X�-�t�4"��Q��h?%�<M�@� �-%�:�Q���M_�%����l��e��D+�c�#[��V~���t�{yJ�0��/*���<=�;:W� �,e@�������9KH&�HrH�:u����)�O:��ZR��<H'���rS�C�P�/Z�Z*�s�!�.o�p^r��U�&Ȟخ��&R�'���UbiƳ`J�U]]�@n��  `�E�fx��4��$"��U2��.'�+b!r�3U�� Cf���f�p ��{�p��U��њ=v®EJ�T?��v�-����t�A�o/�0�m��j��tڪ%�;I�,��(V�\�l4��Ϙ�Cҿ3��7B)�^�T��NG�_��y��ٺ�+;���z%;�Mu��b,�ˏ�"|�?[���%z�]\[͢�NU4��Yq��(���@�^�K��8f����_͸׳3K@����#���Jk���	�m�E�MQ�	��J8�z�����ܐbE�
2|�8�^ns�,�)�`��9��ޚs�u��W���{;�x����#<�,��iVAQ[��B��v�x6-]{%w�D|��i!�mm�x�-Q�c��D�}�"�^��*\x�AR��ȵf�����^1����&�6�v�6�0����+/��JU,LN����?X�Xc���g�S�
O��e�M�[t�%�T��B|�E.T����>��xL�9��P��I��9R�>ɾ�싞�g�4P��.F�2�%|Qo�%�Xt���ֽf�0������S�7�B]��מ����Z	|�Y���Q4�� F�v$xoVnP���P�,,��4/�9�5�]�Ȕ?t1��Xڨ�N �jjs�#������pU�$�ܩV�'�V#�<#fSpl2q����k�(#4��	,iQ�6wc�e�3b_��� ����@�p
	!k��U��������g�2�[��cq~�!���FzD���Π�}L�g�Ϥ�C���$Yp��:�HH���<���Ϗ�"���J�Ș/���F*�ݣ�0$?0�X�w(���1en�z0X�dػQ���|�7����=V,���i\��Qm�����T����������p�q�|��9d�G�[��8$�E���½�X�}Co��5hʫ4�ϲZ��~`�,����qO��=�- Z�xr��As����ؓ'�T�q�K<������Y�`a�s�,@�>�, �CL��:iLt7"���N�_�w�W1���4�Mk*W��)�C�+ߔ�e��0Vo_�@]�i"�o�Uƾ�py˫�'��sq#�K"�n*ܱa�pn��YR�Q�.��Ov��]�f%�UM�F Nq��z�i�}{l:���S��w	��2�+�7P;�]H����	y,���Q���;�����PYpqj���d�b�o<}�&����n�� 6ҵ�c���zm�I��	 U��J,+j#�!CR*��m��'7;�X���z����"�Xhc�&g�L� ��1�亮7�1�A�_�;)��r�qM���t[!�uE-��4��{�}�t��p�ًE��)[�o5V����T��&΢L��z%�\�lP?;���/v]�3�^D��!��������6IrV(_������@>�ͥ�7OW޲9����+F$����z@H�8*8s<�QL���&b ����u�O��B+�:JR�)Ô�<�{��^�1fH�W����h�L�L-����.HK��M��?<�L��cakw��8K]먳+�_��.��5l}[\�����zs��S����* ��k�.K���N5��k5�o	�dfz��Gd�0NKD��4x�Q�:���:�;�(�