��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aЫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��ע9�!�"��F�Wnb� �i��a��c��v�Ϗo@��Z2�[�Sh�+����,��ơ� ������:�������
^@.��/�+7�CdA��#+%Ī|�$3=;���[��%�H�����P̘��N�3���M�v8�;�=�YFz΅�ծ����-����]�Ц��J�����bgDI��j�6���Vż�A�&\����L�t�^�m�5~]�S/�����[�ɛ32ͧi�.�^�jWn�=�d�/vgRD�~��E=?Ȕ�M#
p��j㻵z�	ķ�X,�YzIM'7/Z��P:y\
���T6��,�T�x�9�O[���o�(J�k�j����9��}��c�=G�'�w� ��;NAT|׹W��9���ٞ�3R�n`e=����g���4aM���P��S�:g��d%I�,�M��e�����Sk+X~�~mg,#i�� ��LWt��mu�"�����]�cI�r�jZ�[��+��ز S����'�K)G�Kwom2Y���_����lk1B�ɾ��Diw'�8X�|˪��!u"vJ���|а	Gw .�"4*���,����L���;���rݼES�U�֞�����m#�f?��aCZr��pa�z�{��/%|��'m*S����@��v��@�w�V&�u^�'4sp�%����R)ݨ��\�|6e�d�����_~L�ո������jm�&`2ێ��ڼ&��᷄��N�����C�, D��(��<�w22��w��k3��4d�����zܬ�5�MyY���H�U|��7��l�i�F����"����:��=��*x<�T�̿�]�x��? _Gꑟ�w�X+����$�Ӣ������qʹ,��E���K�xR@���«j7� ݍ�-dQ�<�C��0B �q��X�i��=���!�`O����nP��/y�7�=�lA�Z�q0�3��#.'~���/�o�t�8�P�,�����M@ʴM������d�f\��D���0�#����$VZ�R5��)�DD@��4
w/>�����|3X0�j,M՟����'��
��9b����>q��1������ I@���8�0HH�rV�]�s�������<2Rڥ ���F8v�������֖/���K>~�֞p����r�������S�*ky�����P9+q�b>;O#�	DƠ0q2�p	�Ջ�0�HE��A7W�w/�/�6�\��;����f��h���a�;E;y԰���L����h��D����O*��-�R��OruKL+���9T�s��t���9�"X����Ck�� ���FƊ��/�c� �B��꿆q)�:p�7[o����䑜����J��H�����-��qE��^�ԅ�j�)t�,�c�W�gh��s�[c�[�\����KX����d�+BSlT�ʹ����u]�ۯ�8�<r��ҹ�&T�?ҏ��LՋb���
���䠖r���$%��?M�D�|�N��#cY�;�d@0+\]d��,��%��5N
�&�� !ߊ�_���R��Gx�@�,TY7�9U��Y\ޔ����� �6���V����Ӕ}���s�)�9���V�ϗ�;7��Zd��\^ܐ|���2,��y?�,aՔ����N�h�EE�Lf�8�f���&��u�;3�C�Syȓ_���x�j��KG!���g�_�Y�[���Hq��7��P6Z�*��6���ͥV��"�d��Q�ݧf�}��/V���5Fq<}����
�)�EFE@V���Ȋ�K�3I����"�ͭ�5#
B��' ��>�������'RȜ�<��5����+��z�{�^v6Eژ��tB�2Qǖ�=�:��#�C��{�E����'t���@L%��s��GC�o�2r~�	_-���4������f��j����v��5�ゴ�(�g.#ih�h����V�^s��ry&�M	]�E��p蟊�I8��Y�U���b�a�};��B\qg`;���q!�^��yF�H����c$K�J��s)�Rd�xt8d���:ՠ�N�&v}�d������Vj�SqT��4���-���é?��%��eL<���@O���S2��C�
娜,�����w)#�[��(� 1j�$pE�>�,���u�f�x.lP��`��:ޙ�lv�@��؃��ϿT9-�Ւ�k���.x{�ˌq~�G��GA`���Yv��w*S9b���z�s��������L�!��8�_ըIȩ�vk�f{f��ݩ�H�G�H�f�����5��tQu�D'��
&brc��i�q4�nVϤ�%I���t�5j��N��;�AX�7�p����+��J�V�t+��
0�JbQ�:�1=��|����ޗ$�_�M�+'�-��㦩���ߡ�H�;��K\�G��Dו1J�}NY�x���;�E��\�D�6ě���n����3bDoF7g*�F�����.�1c��9L=
.��������rlBtsx�Gb���̏��t5
tw��]��ԕvK?9t��f��
�H����5@����*�VT��)�P��K�r����1��D	V�����2�f�A�L�	�O�#��8/W�\s���1���2�O���4S�i�|�EZ\0�,4�;�I,pQ��ZJN�
AK$57���w�=����p�ͥ��6PR��7��Ok��{}�������L�d�?-����y�<�f1��A�����g���B|\T����[)/@�Y�(��1�V���s�	}WJ���W�2��mDآI�A���S��`�_άc��jB�o�ߢ���|�ȇ%��I�|��7n�-CR�(:���Y�� $aU����y�ٝ��~I�Ƽ,(~�	�`�}g�dx^֢�����U�}��ѥ����N��C�2.���X~��gk�9}��X���e��"gC����S���"���nS�Q4�:x@�83��&�on��ʼӋ��F�I-���-��}�iۻ����U��ڒ���.��멃+�ԏl�cc�����u�)�2r�"�Z:�����7+����z�S�I!޸����c/����ą�^��t�0j��!y��>]oޖ��q�=�T�cC��ouyB>��ޙa����ﴌM��S�_����XxL4���4��2��`읆�����+���1�pO3�_�E9�����pz^�	U4��2�� �����q��uZ.����/]
��k�� 1�iHK�ٮ��i �ξ�۰ע��ޱdc��?�P��TFR>���]��[���i��N�]tt76biL��<�>��Z�Z�"�X�E[��19��y�r��K���lՂ	 FA����ߥ����:�!�]�����I|�l�WW�E#���j\����ws���C=�G{��`�P��v�,�;��1eߋ�6w�{�K�Y ��VȂa��|vasv�	��+n��C"fH�>��)<��9J�$�ɟ�H�u6�I��=�z�۽���x�ǃI���'U�:�=#��r���VB��y�*l�SS[�5bv����1�y�Y;z��3z�X���ەDP� !
+��|j�|ZN��cQ�+Q������oW��ƱJs�CX�c�qS�j�2dUPCɮ����~�<���&�Ӯl�2��8"�o6� �V�ݧE�̲ry��;˞Y���Z6i�q~b�_k���Y�7{����)��
��!�Zd�	��1����1�F���鉶��Ŏa��k_�Hh���P�\�����#(�Q��9��R3�"�_�$*9�rMpU r6���$jq�N�\�۫��>�k#�04�:�Ke�0�Lp��-�8��ڴu��5�wI���?�?��(�����G�G<��N��r"�ml��F�����Ö���V��&c�_<���s�Dw�э�6D��}�X�S[f�8N����7ǹ���x5] ��gfp�z�FݗU��+$z*�ƣ̈́�[�"P��b}|��Xk��e7g���g�/'X@gՆ4��.�