��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~f�$L|�#_��.?L�|��Tz�:b�������U���l�u\yJ2�����t_ Ķ����/�µʐ��q��$�Lx�f�V��6�f�^.	��M^9�z^�C�	�m7�S0Y���WIc���&|�p�8�]�=IrL�ߢ��'k�g2��l��E��f_��R���GkR�� ���_{�����KYJ�~�]�P�2�"=�_���1�Y\ҫ�c�[���D���ºSt��s�t��\�j�硷F~�@PL��0Q�C](Һ����%�l�S��I@�l���� ���4��EUc�)�����*A���N�o��C��1�o��3��;y?��ꛩ��f���B�@����C7���2�`ɏ�]��m��o��4(�]�c���m�iHrdg5�g�B^���ĦCT�(@݂у�k%�Iy^ĸǂ٧h��gfi$���N�*�g$n6��m��G}��e��SWJWI��S��{k`�gqf�-��9�6�S���f#X�υ1�`|��z�T�e����GX���	l�5��\�3:0?��Q���i��N��K$��(zmCa���������r��؂��+��n1mw3�ݸ���E���������0~�o�_p�[m%��3�$3����J>2E���Dr,�:����(A;:�����p�<� U�I���E��uHTt|/����O��X�i�H�D�9���Tl[/���
В�v򶹡�VB�-?�3�!��B�=��7�����n}���>�����]��`\���'����=>�w#��Z�g�w�ܯ���itF�|]ƿ�C��O͹�~T�^e+�x�+᪌B��s~8���E�۠���v��_ֈQ�c�e≽���D�x��?��o�E��@�+o��7��VC��zGlm~O��]�2(�e��q�vm���yyZ�ڶ>����vb:�s��Ȝ�Hp��2�I����Ob��LK&:FL�&�.i�{i��F��g%�72�߻ԣV��*R%�=W*�d@����U���/#�z>���<���7)�ePϕf��Q��
I�عC��dXʯ�6Q�� ňQ�)��Z����.p�� \�4��K��~s,u2�t��G����"���8�������;H���)V�7�#y��'�/����)3��87'�'1�?/��RC!cv��J���U���hB�~f��F�w�}�G����8��aV4͆����w̧3���{�6��.�?k������b��o��1��愎RL�|��a���]�h�1��w@�0�%~k1Y��p�%���ش\cj��A���0gy >VR5כ8��;�XA&a���Ɂm��Oc���ʒy�Gz'�q����y��4��3�ߥ�%���WC��v����w�~���<�r�H�4M���󿪖-*m���'��)ʫ�b��7���Ti��<s�O�aJ��_�n-���3�Z���	" b��A�4�^Ԥ�EI3}�2��"iG�_R݂��=!�OW��M!\��>䩴[�8 ����HsJ��B�8���)�1�ا��ڣO�8���oP��<�=�F�:/t��Ä���؆w{����dw~y���K�`鵡�r�8�NOn�"M�J 3������R�d�JS�C��р�O��Gf����)�c�_p=g�i$�Baa`���/\ھ��Y�0�ԑh6Dw�+8��(�����6mz9�"�j�LUDCH�����SUһ����=��va�C�!164���%�[áX�K{G�*���%��U����ױ��X��	����\�U7/�=Pa�B*�SF52�V҂`�f��iw���ɺ�#�]5Nz~}J�J�h�P��=8�8D���a>0B�6y���|"���ǣ(�<����[2n��G(��a�Ry8�n��A^Ȕ�d�ʷ�����y�w-��������.T?������}k�:�.9�r�y�V +��Q��=�pű���KO�����bȏ�{�I�5c���;���1I�`VV��c����԰��j��Ç�J�$5��q�1�����σ_䣂Ӿ41����vr-&/mi��1l;���tr����>��ZnS����`��a�&�u����Z%�[�l�?��U3�!�t�SG(]p��R�H�N>4��J ��`��"�W�&�e[*! �.A�P(��������x;������$b0�D�m®ks[�mCdC�I�&h��N�^ِ�@t�c��l�����-�Մ�28��q)lU
m~n� j�j�TW ����.�"�b�l��\ҷ�vxĴ�5�.��T�wN<ѕo�r�H�T%�= ��Y{/����$���eõ3�j�N_��$tL[��<}��"*�Y4�բm�:��i�ǈf�#�k����ĉ{�|��=����!��ی�����,�� /a^�s��]E���Dbd�����B#�Y><jϣ[�#�ؤ��/�n[-�aθ�7�W���}���z�_苯m��ZFt���ͻ�d��Fg�66��_�$�BDcu)�_q�+:�)kUv�]a8�8���L �	�a(u�.��Lƽ]}Z���R����e��슝!�Pd_X���s(�����fH�����q�3��˴�nP̈́�(���zS���+R*��p;� ��r�w��y��
�N���MV��}�8
��K��
�[��-d_�h�1����0`G����:�_��|̰��x	��o�J�3�2 *)R����mH~ǰ�]'+'��,��>�@�?�Sl4Mڢ4�J�����e�6`̛
_d-7#SEB\/����9�QΕ�N6=%d����1�Fz%���[s�.��^��0������Y�sb~v����;��T�s+�z磅=�R��r��o�[{�(Ѽ����y�>Fa�7�f���j� �u�:�N�9��brH�7�̙$�6ϥfzK�\K\7e�}��6�8*#H��V���|����