��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������f(�7�u3����a8r�˳n�rd���7�i���@L��&׳=��7En�����������M����e��Y���GO�ʎU�n��a�MT �H2��]��D��w�3&z�PY*}ޡ`q��~�����\>�'�(����0O�]Ŋ���_�H�G�88݊k
�V,$5ۍ��,���`����9��:dl%������Pq��M�zÖQjƱ�:��e��r��g@��䓏})ha謺���~c��-i��@=��G2f�hT5�=P�!�i,��J�s*.�7~E]�|�������0�e��O^�;T�ߘs�`�+ �(���pX���"��pR"�I��?t��2�?�P�� u��4��#A*��'섓��xl�sɁ�<�q�82�;�&F(�`��E�!:Q�*a=�9��Ve,#��}%�Mk�,N�z���b��\�g^L5��T�#�Fi�h�
��t�Z4��.�
�'@�ƽ���sN��EX����}tSt7�SX���D?��hП�9�\n>1�S�kQ��Ν?�ಎZ�Ip3�8\��
ouf%��
���HN���K�.��w	�~�OON�2�$����Pm�`�b����j��/��RvF��ݡ�y�-��ۏ���=f�ܙ�|�@x�w|(��P+�����c4�~�NȍPt9Puk7���ߊ�b�+7��v�qG�B��E_�m1�2K���0cP���'د. O���y6P4���[H�9�i�6Ps|F�um���t��3�.�o�wUux�=���=��b�E���O���G!��꺟��W?XA�CҼ��ޏ4w;ӫ����T�FV��V�~�ę���B&+��QZys��s�u��	O���q�"O�w��tR#\�β���d�'���`����E՗��X��u��ߺ���@X-1���
�f=0n��ޟJ9W��^�nf�l��v�C������24-C������Wo�h�i�Q
�����`�j���w0e�x��sv����_<�OwJR%�w�ݑ`^��RK$�89Ճb�% d�\X@�f��j�9��s�ǿB��X��T��F?C���#�[1�C��%^���-(�S�j�F$o�<KK�{��w��-�L�Z�E�IH�I"T�f����X��5^{*Lp�a���q?���@ZD����7׋$%ϻ@��[_��ˀ9�����Z���c�̢��R�e4Y�ț�N*�5[�8^��7��y���Խ<�0����F@حo�&!P���㩦H�ǃ���"R�{]5��E��8��̿�9o�h	�?�_�����	�r�Ԗt��Onѷ��V���1�o�j�yi�壘�������T�[P;FE]Tv����R�rX7�55�y�����GYUG�&e�\�%H+�]J٫����ZC�#a(��y���v3�m�Hb��g3�I3�"HǜOۢ<���7}�qW|�+}/�����Z3.r�����̽Q�����lN������N�Cޯ�S* �v�c�(ȣ�Ud��P��K ���ķ�b�l�>f��N�\������g�OT��,0�~����-�N�PC{��*:�: ��i����ց�<\�5�oW��ɏBvl}'ө���D�f�y�^�0_���X��j�[b���Y8������AM�;�ZY�a��
A���?��ns2dSx��c%�ڼj;�*>�/��Z$����]Q�gh�_�K�} �0;�0�QvZ+ݑT������7h��j~��ԅ.���"��ulr˼���߬��gE��#�6�<<i`�Q���TJO���Uܦ����S�\nJ��ן	��ֱ�|��+Im����Rcr�1L"�(j��6����=�-C����:����Vۺ��9���k�opj1{�'O��i�Wq�U���!4��[�#>�1��K1qb�C��92�kk�0wJ��UYC����S���:��8	o?L.�s)ϱ�
BdEk���"�n�)�)��u�y�o��M��}!L@e�D)H��������l�-�Ðvu<!p��Us%iRj��M�J��*t���v�)�Wף�i�5}����O�/*[�����S�+���/�G�ϯ�w�DA�,{�P���W���Ѫ�����<������cP�'!�I�����΍�	NA�a�� �5Vv��H����烌�!�Wp�J	��{/�,���"U"��8��F,��Q�'�ɯ�fв���������r�g��.5�:c}k�ikz�*�ג<�����7���C9�|RdgH:`u�E�w�sfnQ&�V�u�*\���� (���8�)�Ӡ�Et���5=��}3�MX��=ߋ�5�0��1��)g�D�����{�B��)�{�F��!�L�},t*+F�b�C��t�"�2�7ٽU��Db�����U<�q���3�1Ar[@ *���ᾙj$��8�����Ot&���8b���
;���#]'cg��YD6mَ�������5۸/3/��ϴWE�~���}��p6���Y��p;%$h�2S�g��V]z����bh�X������r��t(n��ԉޓP�����#��E��t�K��8V���e��xlV$���@�$��11�����9�`u�y�z!�-���qZ�����.�c�(�������Vhe��YT)]���3���n�^���crA�u� �7�)̻a�j�$��y�CA��0�=��;�N���V�tU=.�0���R�?a��}�"c�bo<,Hez�OG����OVܡB:�'��жל��ֻʥ�p��)�;�����V�^��8d�wN����=٫z��ޭW�_7�2��°�����Q���j���0"Z�ŕ��������ZΈ��%� %�"�̽*��r%��&,��!M���[��jp��غ�{��g�{�[��^1_�9d̪v&;'d�<��_�G`��^srG߷����b�F�����Q4��͔�r����,�>(K(?���a��a!$oܹo9�l��,�=�p�k"Q���z߆��c�]O�xf�=����B�RU*'oi��{�Hz��o�ޣ���4��r�y��#D�;�i�pnE�gWF
�Ώ�2|K�T���M���#Ax��#�o����ig� z��X� ���8݂�Bi�=� �C�6�휛��JQ��%�k���܌�q)��r���N�fޘ�`1�Q?3*�F�Q�a3���ǹ�)̑e�c��Qn�I��"dg�Fݟ��ߖ�Xׄ.��vj��*N2�WǶ..a�f��;Sdh�����TC��+��#áJ�8��ʞzFV�p�����r5Ac��a|Mtl9@}������pa�"ֱ���#�I;�ق$SfpW�'`�Ec�K&0f�k��h�7��$<�i7ыnbq��)Й�?P�(1-pJq�12���P�b4���J�CX�� �u��(O�n�M�<ND�Aɍ�%Dz'�%�Q>�)[8>� %Ek���C���}F	�k�e�e�e�Z(�7۩�G�E4Ք@���;�0R)�`[�(��\7x��,�aּ�=��J��T���!I5��:���E� ��Y}/��TV�/�-n�fM�+ ���rVt&a���1���nS{n���Y��s�x`�ۿ�+�np��J�a���;�A���>�!�v��O��A�|T,xd�gP�	��4õ��ㄹF^ ���O��������_�1YO�W�R��?��nvձ�qPQ��q:w.]�kE���ˆ3�?�7iJQK���`<$�+d *�4,��V(˭QW�� Ⲁy1�.Z[�7�����/UP �����XfK�~>{��Q����~H��K�XMFɹ�=��u4\�7M	�C�Oe<�	s�5��1�n� �~{�>�i$��(��ip���� �4����q<w�`�Bp]�W>�)�Fy�x�ݓ�}>c=�Ah�2�L���c�<�Xy�>O��P;ԧ}�vҧ>��ȃ>h���?MV�0m��nǵ�_79sFM�4Y�"b���Kz����xk1���6�ֹ`�0����!��h�7��T�D:(7"@���Ao)|)�r�3����c�P�~�d�mrA���:����CMe��9�}ԷF��b֯�TJ��?;w�l�o£y��'��(7���4j��z�ǖ�ҟ�D\ívm5���9��++os�+�ӈ���w�8��F=�����ݧ00^ �
�^�$5"p�m5��giC9�Ҡ4jbX����U�V��.�8�W����"Aω���������v�)|�[�Rpd����Ic�S=�.���׉���S��Y���"_q>�-��j���9����ȹ:zc,�����#�P�������.����4��"�q�K%c���]���C�),=�Db!1���\ٻ ��@kA�����p&d��
4[
��출P�n�l<B�,9�˿�C���4G����|(��������;Hl�n/vJ,9[�j�\�C/K�c4[O����ԴV539q�&1�Q0��}(��ǟY[W�u�h�
��5C �3�8�(�:��e"��:�3��d���B�c&�U�� �ߥU���Z[W��M)���]#���A.�/�u��$�/2`�Ò���m�\�=g�Py�E�T�s�2���ǊD�Rq�D�
��w�6�_8�~�AL}��b�8$���q䰻��Fy�*z�H��Әy��:�I��4���YBc�[��c�s�CU�H�_ug*�L���H��fg�V���7�5��m^t���O'/����a(�xugG�c7L����T��f���OǇ�%�1/f7�P��l�'�k۬��x�ù��q�5 3��1(K��Ł?Ĭ1�+ �S��ƇF5�1UΗ{����.ҭt�ݞy���Aɸ�0,��S������;����JS���h�kl�	ab��7(lJS���t
Y|�j������Bc;jA>~�j���U���LD�P���9�%��/��q����D�������f�S���˝L'�rn�~Ru~���ߖ^�� zm���Ƨ�l'��U]g���<����Z��\ �fe3�F�vw�k�	�Ǜ�kd�W��Z[7���P����C/�B�}�O�L�݊��9�"4�m�Ę޵r'��p]$��[X��@}F"�e��d���%f��m��$�pc��w�tP9%DruJ�+��D�L&�zoLV��)���Ї���ɐ��\�B��@ۘ��ݏ#䎬��m� �e�M��iK���P�>����KG����+U�nH�VY�Ċ6�w�~��'ӽY����������?w�]Ԡ��`\"-�P��ݷػG�z���˵RW�k{�@�橏�RT)ߪ+!XR�I݇��#�d��p[G��}�q[Z�D��d�f�4�k�R�&W��K��ɿư,8��znӮ�	��:W0g%/U��\DC�ǱO��iE��x�l�)� рܙ'%�u�Eo�y�.r�8�OR� B;w����̉� D�"<A�7�\�B	8��R,�&/�Ͳ�c ��pd������e�C�������o�+ �\#\Y�h+�<��U��͞����hs���/݄�B����D��b����6��>]�J�>�^xȔ���i,��v(e�^����8 ���$ӺKu d��ڴm����JS�Y�W̘P���|�]PU	�s�{�N_����Y�V�t�����`^�#�(�q�K���/"��)&�e+��O�b�����g����ͬ �'?5=m�vQ���ͅ=�����SY����ߴ������l%��ٵX?��5lUF�����m����ӑ礎���	���fSmL��s�����?�O:8������?�g[��ۋ��(׼��FR��I��1$�ӧRTݐ�Ü_�C��v(�<'R㚘]�!�vB�N�hEp����g!���;&t��P��t�mf�>
^���C�Pt�9 �:��;�����8���k����S	�mU�6@��t� 
�L��s���:h톛��둏juB�$��WA-[�"K�||D���A�Õ��:�l������w�V�Ybu��	�c��fv�v�G�u���l�E��J� �c�6� -Œ�hu������b�꿢��=)$;���o��h�q ����h����yU���}bkJ������i�}�h��DA���������Ґ�7s�E���P�\ <�{���8�N���#�_�>�WO-O �|MC���n(�%`B����G���m$�3���.�8CR������̸@CV権�7���3�Ӻ�Y�9K>�F8��\I�r��I�Q�$25XmG���n���s��^��Jx��v/�ِ�VqP7*O��g�uy�,q �1���imE��8�y�S�8��iI�خ�#~b�_��>�����D����$�R�K��z�3~;� g�;LvS+�1��e��K��tKĪ�RV���[��#+��� {IT�D���om��@�ksMJ�x�C�g�Uf�a�֦~��I�zP��D���a ����U�:���]Z<�#�q*�+���;n�X�I�`vvl�2O���l-�ԟLK���?���S,�ʢ�����>O"؋+��tt1�8wJ��.[XX�ᎅ@Tt�g�oR�1�ʇ�����h��K���H��i{��̕mq�/ǩ��>��	�"+9��J�.ā	o2�8L�@��:K +�9�$m�ο�W3"��*Jn#md�[��=5l	$�Q�Fn&y�IKCJ��*ڨ4�uo�
JBX�Q^R��7����'.�r5�Ek��|8-a���m��ՆrӭdΈx��b�8:\O�o<c��$�}c�U�k�I֘���|^("3��U��S��ړ�n�@�VT門kA��{��UaNS�3v��#ɼ�[i�h_F�ur������O��{�X\�l���V�[���VW�]�ߦm]��?�BhC�6�4�o�m�5��38�W��n�\�  �g��D�IH����x�9qx���D ��Fif����P����.
�g����:hW?[s`I��M�ןK�;D��ը�"t�V���{:���R�x�ߓ�ɿ<@�A�C��8�>�]J���r��?>�'�l|Qi�K����!�P�v*7�;��ΐrB�;�432�5�69�>]��͊�D�f��L� >�I��nx(�KGJ���v�,k��y]��w��0��˗�J�
��qa6;����ѹ$^�i�+$�i�گ��N(=�-9PX���d��\��)�D���nܿ�<@��Cb5��5Vv�C��8[0EA«bυ)�<���+��s�b
�K�VU.�[�3� ^I�w��y��1��o�h@{�,�@�hD��U���	$��dU�kTl�������G����cKo	�C˹�dϑ��>f�[���w��M�-�%��7TrVb:��7',���a��G�1f���HB����L���oM��B�f\cd�0��fL�5(���Yƕ�Gے��8�B�fH�chb��z,N�ob�����)��X/�Y��"A	�3��d�  Kp�{���t>Z��;a������o�b���4�5eG0�d`g��-�"e�ɟ��-��e�/䝖��Z'�x�k4��P�q�G�������|A�����IOP&_Y��3A�ˑeUiZ4��K�G*���Z�e��/o���ArI���Շ�o�:�_g�G�|u湉��H����1���sk��\N��˔�]<\t���M�9O3�����������k�)���1����O�F����������I��q��Σ'���Q���|ų+x�p��{��'�{������[��P-.���Կ֤����B�6�.��r_��۷�P�t�:^��v-��������
����:����t.n���H��S�e��ls�jl��#�/A��^G���WM���t��|g���Z�5���V4�U���7Z�||sZn��>�ex�ى��:��X4*a/S~�� ���7Mnɶˌ:V��٘��(�����"|Wz�<��ѡ�c���r�����rH6�������-}5dv�>U`��#������j-+`��tl�!2M��4vsO�����k�NY� �WqI��*+l�qМJUՆ��y