��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e�ҍ��
�$O#��E�Z`���P5L6��P~%���4����x\ަ���Ij�õ7�co�V����mJ?��!������А�ӛfD�| V0 z�W�z�}o�C$�^S�VK#���/���-c+��Ȯ6�V�7w�H�b���	��������)ɽ"�G�衎-*�T�fQ#h�+���ҴV0��]M�W!xO��B=HQ���>�〙9t*�Bi�� �Z��	L��=�Yf)�y�i�j!LX�o�~z��;h���A�z'S�	P ���`�[P
I��:P��`Ouη��W�x��b�ɢ]���_�7��(�u���B�y��Р���'��**����\�"���p|ۯk���dZ��*:�?�7��.�(���+����Z�!�Df�++�[�SV(�u�*
��]�t��ڔ�!�h�\\�K��u�_�$���i�����8����6W�(�A�����ß�����gM�m�lo�0�pR�ac51�਎�����(qPh���k����vj~���NF͂��%Id�y�Jrv��C��F�ᴯ��CE��5�H��8/2�T2���c���.���/��a�#�c����Ƨ�#[���Ҿn�-L��(
C����-@}̔�(J�2�䯱8���Ш�)�u"��U���p�qD��<��[�X���M�v6���&�Yd`y�����d~�m��ݺH��7�V
t��f���B�N��ʈ��laQ��q�����[�e ���ߩ:��.���U>������|�>�^5ه�=���W�댾7�t��A��[wR4�w�Q�ݮ�,r�<K�5f�e�9�u��{��:��X�=W?�;�Ò}�O�f}J��Ӯ!%RRw,;�ۻo�a�[�ڑɡ-{��؟2ν;�3ty[�氋MDs��ǧ�#<?N�UᰊDU��o����)ϡ����S�֎����UV=,�j�x�˖�O��-�0Z8;�`�"�2Q�x8�k7�z�Ӌ(��U�lT�_���x�)�gh3)3�,<�8\n�WE����4��a�o�����+Х����(�<x&��x��*n�&������|Z��D+k���E�#q=0��CW�^?+�{��{lİ���ѵo��:��(>ن����Ӎ\Aĩ�b]�[�D��G&3dQ��ݎ@��u�C�\nCf������B������Z�M���{��.M˜M>�&k,���q�s�=q#F�u�kN���N0�A	��#���Е]�cX���>hO�Q*=��{㭃G.+��!<����Q�&�v��Σ�����z�Y1YŇ;�o"�W��	άH�v���^�)Qd@&�!Wo�{g��M��\Z�������8_(�]��ԋ�e>���@	}�0�ؐ7C=c[]�`��*����)�s�,��q�;󬅒�=��w��?Y��F�!�r�\��;��^Mcy����@�	0�!{m�#պ�����&��iMŕ
k�C�Z�p�d�Åq;�R1.�F�s�ϛR����+��M�L"���Ti�}���� zuip8AVD�N|���vzK�^���}������0�f��W3Tл�&��y����G�둺�%IZ}v���|#���(K���m|�͗։/�fZ*����ݲG�AYh��-��U���L�jf�z�®���Z@�;�������jYB�I�c=��g�UI���}�XB#��s]@;8q10Q��*.���Gr�lF��Ⱥ8��Z|�h!ļk����Ƹ��K�s2�&yu&��.����a���܋Q	7��!��	�,���h��>n���|+*�Nt7Ygz�B��DW��J���T&�ʪ$z����ŏ��Q��m�x ���r�n$���I���7-`��Q�����Ckx�bX|��3%ޚo����(-��,��:�]ھ`.�/ȅejީ0Q]{�k;�K^I@���y;�@��_>�a!r�s6�v3$ɦJ�13R}1P��/I��dՓ�:`�z����m&���%:�C�cg���]1{�ʔ�ӽ������d�)-�e�;� � ����puz������5!fh��ӱZ:��Țo�Cͫ;�.�S4&��$X�ٕF���C��)2'�頙��M�h��MD�~;r:f�B4I�T1�RBEW��`}��s������'���3�%�S�"x{?zC��9���P����Ӷ����WIK���;�g��c��A�A4�z��褆G�j���f�� ���0�k�d��je�
�^cw�Gk����y��My�j��u^���A���í�²�q���� ��N����Xᷕ*���Qp���H�/��JBL	q�r���9��({��g�tXM�*�Jwi�JNow[�dmv�*9���F����wb�)�W�2L��iz>�_�(�)׺,-D����/���'`�:a���1�Lu�Q�#���M��ێ���4	C�(rE��*����\�[C��c�q�����iS��S��	[M�PG>����n^���8�r��+���s��6!c�P���k��5�� g/s��Đ��Xaq�����C��'.�fm�i����/����l�/����l�'���={����h�����i�U�ĀY��5����] �,�L�mc1t^�KطC���/ǝ�Qh��(��U���J=+ �\LE���cO���-�%�^)��{�JMt�J�~���1h�$0He�K�T������3�\�:<@��5 ��K�;J�����Q�=e���co�G���򆼜�jۻ�e@�z�����o��N4����V��yJ����yD*͹hF�oi�.�:���y
IǖQ�XzPm4XlQ�dhteiG���JH@߉��^���hm|bw=�v�|�8_���QHh�NS@�.��a���S �\&Ϯ��7Q	ηCI�����]��jP����+�����8�����a5A:ـ���ʷ��3��P�ln���W�Y�6A#l����^�w}K�z�^ŬgvO���Cs��G˪�w}���Ӛ�ƈ[���;|'�X˘?@����MG�z���GR@�Հ�Hx��Og���m>`�
P�����3�ꖔ�U� ���&d���υI��J�MsT�*A��������_v�TiJ����q�N��Z�U�@��@6>ӝ�_	�&9�e�c;fdj�hKT���Jx嘤t8{������x8:`�ٙ�dN0Wk|�`��}J�L��5���kS
,�7�ؽJ�N�Rڻt�Rț%�.�w�s�X�������×�6؅�I,�J����2J���1�muQ���2�鮶�n�Z���>������{ĸ*Cë`[p�p�$AN*���/O[{Rd�� 21������ �׉)jS��x�i�R��m� ��Q��$��!���|�M4O?=p?�C�8�����=&x����� �&�&X�Tz}0d$E�"��,F�Fjפ�����颞��-��2|ϩ!��kW��}T
��cj�P%B�4�"�`=p� �����E| �=|y��j8M[�Yӏ5�J?'���O�'��+j�וL*�(�ӷ!�z|FTq{0��U�94{�-���u�a�4�a�����IQ��+Y!�^��Z�p�m���On��r��Y�j<"Q���u��u9n���mk!-	�H�,}1��F7ZBoU��<�3��v��{���l��Y�d���$J��k�H�9�--��[�hv����8UP��'��x]ԥ#AӼ*�C�?�}��p㯦ϲ3'�[$A$Xum����޵�
$+�>wfW����Lp�N>Kv.��w�0 ���y�V��?����_"����t�y?w�s���j���O_|�`�����N(�ͮ���s��� 쇗�jH�@
bEj�.I�����4P����U�� O=�H�m���ϔ#������.����K5��wF�E �WHl�<;��|��y>��>D�����pE}M���v��F�f�JR�$�
ma;��}�)� ��տ��ZJ%T=;���*`�]�:��P��Nʇ����Ed#�����L�ϊO�0����^K�9��~(7G|_��sɡY�F�����\�-�Oq�D����c0nl8d��:[O�?D�v���d�ƶ��G�p�Ne�h��Z
k���:�����5$�5b����O�ْ�})�>+1n�|�L6��E�ߕ��ԅ�FP�;�B�ۚ~���5�������H��`4ս2��q��M�����djlF�G�Z3���ns�S[���+�*0]��dT��IՇ��9%F�����gu�e��y��lD��c�]��7�#�(��^@p���{��+lq�K�Ԝ�<㝠���g�bH?AX���e
4͞�X���7!�x�B���Q�B�K��1:	�B?f�rj�q5�d*"��Lҧ��h��+>��b����H�ʬ85b���8�N�|�D>29�mn����� �bp�e��;�!�����&W�?ȉ�~����Y)��]Ђ�޶������z��*�*�<xd����k���z�+0n�;�u�Ey;^O��|	�;����.x������Q��j���~3n�t�do\��#&4�D���)`�ae�]���v�ƫr��F�����(g�G�G����щp~)���\|#JX��a���P4�/w����V�-X�0TE,�܉����"9�(�ew�Z%Ƨm����C3�V�w��jGt׬8�g��u�35�?2�@-���Ǩ�5	�	$:e��H���>^�6����&�!2\���軌F3�R�����Qk��<��R�)���\+0���s�!W��a_[� ���p�����Ta��a���ͷ�CH*�+D�i!�+��O�ݎ۹j�����b=�/7� �2��t���0��%n��3v;�W`*g�ɒ��&me�T �I_9���F[U�yL�\4�yfvG�����<�w KA��"�����V6A�����]^��<^�Lgc3w?U5�b-$��u|<��~Rf�7�Q
vr��P�O(��%-��N�jt�{�5���UGG�P���6g.���J�8�Q���P�9����3�xY��^b�mpƾ�;���f��!"�;�a9�^�������pH�d��oƚ7V�m��� �?���E2x��=Ḑ�螭R/l��+,e&�o�hlUʠ��I~��ZR`>��ZF������1ZƳ/��8�zR�V���S���]�I,Τ/@xnxe9pUi����LWV"��;b,<�̹鬪L[�����y_ Q�09E��VY��86�r'�-H�q�/�_���Ԑ��y��#%�_kA������*��.S9���w[��T1�F��pAѫ�`���o���~���f�������S?�y����&�e��*�mv)\���Pқ�J��Z������0��M��pa�(\�֞�,
}�qd���E�m��q���C�5y�p��b2}��˻_��`���'�*+��u��4�۟��]||�#X�գѫe 9��[��z:5�����9�|s-�����!b/:i�_�s�m��^,��N%�Ώ	e�˧.6�⮞f/��GV�B������	��`w��D>8!��C���Ȣ:3߲Xde�����,�0}N5�"��}�R1�7i���f̺�9�x�yW ����g|=��a�-ۄ>uu�t����Q��q2	%�n{���}��/��g��c��1��UI����3O���Ʌ���8��"�19,�r��VH�:�C=l �܃2�:d/�[=���[���(�Z)ȬR�zGy䍛���s9l�H4
�	y�F��p�4T�p�/1����9UD�q�3�kl^����|�� �~F ����p�O�xs�.��͝T�-�S��Z�I��y���~�?�����������:���/�`c��T(5�y�z�AȈ�5��N�BY�&���/H8���i���̒s���İ�ݯ�H��'X&~���o��E�����9�B����Kǜ2Ѻ�~����i� O���E���r۔��Q���#|�3��^T�;�\�+'���v���L�ʯ�9�C:j���6�bF��خ�n��ȯ���lLs\�)��`��<"��H&�\۰꒚���3V����Þ��;��He���6|H @ߍ�|��E�5!O���(�ew��An_ܽÉ����h��ss���PU��:+�H㚀`r_�-\��Mvw�_�t�I�tzC�%�x�l8/�󖬎�W�y���̈́ߤFσV��(-Ôg�^�[�v�=3)��g�����l� �% a�9���E�#v�Ig}���XLv���ѵ�`���·>�;�6����D�F�M�b�GϞ�Q&�>qg�T���}��={�$��&B���-M�=΀�������ޢ��������@;XM�X�@�JS��\��d'MQ�*͹�p��_4�k6csƿW9��ު�~L5�uP��bG�B�x�ǳ�/㢯@��`E|�]0z֌���m���	��P�❇Z�9�#�IKݸ@}K'����qM��@=xY,4�	�R2`�Wc��u^v���'�kWp�Ή��5>)>j� �����ԋ�<I�Rم%p`�J��G���4F�kwB����T	P�;{�䁯V���r-�"U���f���l���{X�B~���PJC~'�5ߐ`�0�� ?9	y2��	-�k���~N�w���2���+�h	2A�� �mɷ���;3I#;�T�{+t]�_2����f�̄U�6��*���:�Zt�;�^��8�E�r�����0úX�8"|p�y��yY,WH�B(�����e等�c^U`�<�G��6���S�+�� �=8'6�9��N�׾�_��l��'��X���ˠy�%r��zL]O��m�N�J���/va��T
��	����-e�=c��+���%��W)Ԉ'��A՛��n�	���8d�6�Eq_���"���������S��I�e�1��#��9<���q �׼�rh���\�&�ИԳ߼�0dԃ6�J�P�{y���hJ~5���x�=��u��g�[��v.u�V���=K���û
�5�"'<4j��"�}�PF-XՈ��N�*u���J�T�N��?���|ڡS۳��g��	d��o,���~w�y��+�[sٻ���V��G��7&Ԓ%Z�Ҏ�,:���J$s��ŕ���jg�_�<����_� 2�^`2k��2?�vIE{'���ҥ��m.W^�: $-6c�x���k���&��.h&_�GR3��2�/	���Wc�j(��e(<�z����!@�*,�:훗A���N�Մ���3ev�R-��U��N�p'E3�*�a���d}ƥ�\®�xizzډ�I��Q�cTE�q��~d�Bu\��]����c
�v�v� �r�zy�t����Hŭ��?�Y/���e]wy!���F�N9�Vp[!Mڋ/m�D�Pu����23��c�O��bhJu��r���\/)�vC�'��nq<�=		d��E2������}o}�i�X	���T뙞j�"`	�j���20��v������RI�6�Yv<���3���H	G7]��/�R� ��JԴ�QB��������,�2�-O۔W�K��x�����KP�����������$�<��'���6��� �MςmO��F����w�_�gm)|��֒}&,z�a��:N�%�q'�ܬ�	���H^��)��l�V+�4_��s�D���/]D�H�g�O8%?��:C�Յ�`�}��ǚ~�&��'(�eW�9	<��\�L�;�	4&���6�=F��iG��@p��ɓQ����H�9���ͽC��R���M��u����p�&n"�m�)x�v���}<�[�pcH6צj�kB�!:\.,]z��MM�|�m�0:�F㛇�E.D���껫v��?�O���k�H�I�2�����T��SOV	���9&6=��R���6���FFm��ï�����<ʒDX��* ���([�5i}�0��̙t�~}>g�n$َ�1DM=3�W����,g�Sⓝf�����G!���c��,j'S�w��B�_�A��%Nk6t�3��Ħ೙&25�c���#p7�Y���;���)�{5��)���J�u^y8�f0�E{F�L�b��8�Op"�G򿿟v�~}'��ղ!�z%ᵀq�����55����`1W���� �`�_v_�W��p��Kj�T�^bk��Zk��L���z����� m���l�Lb�d|ϫ�n�0��b��D�)U�2*tKO��9��0M�H��F��6 %�Ă9�S'�ޘG"��q!������O@��Y��.�*$��'�2vj�N$�J�̦C2h��b�%p�
e��/pr0ҳ��O�T�J���o��eyQ�v«<�PNc`Pfȕ��j1��1��[�9@�`������nP[�Þ�T���!��t�M�h����YOw��؁�� Mg-��e�S߰ 5��MiĚ����/�����-�F���m]�u2aT�h��z3���N�%V!���\�6[�)�<7<u����qk>R{ �@p8J?����.v��`P��n���R�8���L���O���natXi�Y�&��dW=�a�rc�	�B���@j?y�o���v�Y��]��~�
��g�2�	���Tf�vl:H�G������|�ZS��[���	|s�@e����y�v�+p'�J�6�Z�w�=�5�]N#�N�ޗ�qi���ਡ)���xq�� ntFT�f3e� 3'&S��7���1�a����Q���{�x�G0��覛]\����{^;>|e��1��%����D	����K�>��`�}�2c��d���g�qt��z*Tf�<`<Qq�Ej,A���\p��\��t�w��GJ���"���8� �����&�"=%��R�jIΠH�ۿTB��K",Oc���T�{��U�l_8\���,T���������5��1M-�+[��k�F|Δ!)�Kk����0��(E@ lq�ޅx����m<ʇ�᪣Z�/�/mj���W���%o��L�P ��H	U�\�)EY�y�]W�R,��t	�@iF�5�F��4�)6�G�����Y��g��+bO���R��}R�m:�(	�{]J��W�ʯ��o�M(4�G�z�}�f�ԥ�D  ��-���.�'���¤��=�
"C��`>%x�t6����4��������mJ/�9(�^臰<�w���s��'g�e� �>��Ue��$�p�N�&�w-}��~�0��o���+>��J�/+�e0�E��<>&��;��L�LV�o���l�����>�k�vo�|�s��{1r_6����ee���9�֦4L�9d&��%�O*Ȃ#at�T����8�[;�*Ҏ4L��?\FA/�gD�.���?�X�ܑ�<I*�s���U9����J�y�l�/�[�	U�wXOR�H-q�`,t�w�z|�s:��@�X8���;$�~��!�4Y櫽�zǙX%�h�.D��Ppy��)�V��S��F�s �����a�m�����w�Q{x�$�G��#r�t���#���}R�"ڕ���)�$P�čO?��2�&Z��pmʴd2%n�V��Q%���� ��t?r����R�A}�AW�wF�Ա5�9/�<�Vޝ�yI����p#��"�2S"C'����=�,���5�	�(J�)p3��9f�ty3:|��O��W��"L;�9�J1��`8��:�3U{��":[��U:�t� B���v�Y�|��u�L)R�(��"�1�w\D��*��@v������z_SE���.����2~O���T1���~�'���K��NDv��@�%+>=�Le�j����d������巁C�+m����%մ9�b�~bۜ���J�>4V�پ΂1�/|���p�z�MɁ�hz"����fcD�z�2�͠��i���
��i{�W��F���ǒ�Z�Dt\��Pϯ�f1ϡ�+���c��z��KE<'��}X]�(�b����>A	=k����Dto���}�!s:.�N�����B�U���4��i��45��!� ��5H���^pi��90�ef"yR��xZ������������P%"�j�6��(3u����/�
��	�>;��-�����t��em�>ߘ�M���~�{ݜ�d�O5���ʻ2BK�2yn��հ��d#�P��B~3����m�C?��On�AYc���r��}�ǚ��M�qp��Cv�/���7��o�����'Ц��b(w���N"wX�p?T4�M�����EoZ�I�S}���ٖ6|8SJ�!j�a]Wn�Y��9G{r���/�_@���W�]�2#:�A;c���;u����(��y�� ���3���G�Qpա�����*p�jX�9^M�L�683[�|����~��u��_ϡe���!����	����o���I�T�̯�}?&�ƛ���o�y�C��Y3D�'&�y<s������-��C�(��F��}�*�9�+c"-[ϊ��҉�\[�Gb�_ʊ#�}{U�F�ϛ3�~J[m)d���g�4�\Y;��:_m���p�fU����\�Ur���6�e����B=Gg�f���x޵0��铕��&m�~Ĭ��>�&�Mc�C�<N�y���Y�7���N�{ d��-�/����ԗ�4[���w�K0;\-�����,����������S����J�`�VwU6��t9Kk��I$d�n~J���'��g:g�0���a[J`�m���J@m�pp�C\����*��TxP1q�%���AkŞ!�m�-����"�"j��YWz}W����~�tʨ���ͪ��:F�XZl|X���HU��(�3��u7�K�C�qO�~ �G(���. �7/Ѝ����톙��F!⿥�3�Uw,�?�8#x[p:�9��j*����^�K�Yv|#Ӵ�W_yO-_j)�7�O�9����;�"o��_�?�p�0V��*ه��dd��%���VRmP�֡%��}��p�ጹ���$�ը
�eJ������]jޛ�pU�*#aZ���/w�?�ք\%^��L��2G����e�q��5�IC��&.��o��E#�C��MކS1V4�)�����SC�fL�J����C@�u���'D�j�R6X�h��,������%�l�G,����?��9x�@�g����%�QCH������Mg�z�W�����%���W�AR�B��4��� �c�g���#,�h42��hx�Ɔu���i�y@erlk��zk�q�v�wsR�	x�{��}P�-�29w�	u�Ĕ��A)�7�@��+D�I<�p�?��x_\����6ߌ�Oa�		}�����!�򉦤l��1���!��2%��V����:�~����G�n�r^rbT*�e����fяm���rړL�������6}g�u4�dH��yj�е�2�r;�c��6��FS��#i�V�g��lm�wO ;�XC[���`�^�Ӷ{t�L�́�a�1��r�Cu�:_kr�8�������'����1T���dK�60B�5� �5v��Ы?����A��G�I("#.����D�ƺ�NNl�1�i�Y��?]�/zp�;���i��B��+=� �Ṛ����KC��Z�r�a�M��	Wj;{�a)�o�#�4
V+�)7������pY<T�=�M#���ǰV�\��L�B�_<�nH����c;Id�1�6��=�Ɖ�JX��ۆ�!Ʃ�~�}���P.���*��Ny,G�1��=�~%��"����޼R3<�H���kt.�1���t1���ǡ��_��}�m���Y�D֠J��m�����㯋�Ҡ$�9�#��,iQ�P~�Vʊ[����=o"����u�2��t��kW�+cTH��
� ���B|Y<RB14u�!���i��������G���.X��%&�ͯ9��Tj��������X�m�����7�J��p�ܸi�6F����֣�Y��C I!�i�E�ݖ�b���0���B�h�v�V\pS	Xf��/1+$RZUq�3	��Ɵ�ڔZ��=`;[\�;=��~�����E'���]����0�{�͎��@V^��X�Q.6����=�FI�S?!0ނ��ꮂT�m�nv��b���!�9t�&�36���d�7\���Z&N9�+�#Xf��p��K�ĥ�v�����<7k���P=��~a�����_߳M�p(����%���"�m��N^�o��_���/�lb7�%���5Q�#����O�S(׍_�r���V�1���l�*��-��wȳX�<a�B���z��e�79�$�Z��(IpTymZ�cX�-fp�@l:� >K����1�@���
��oթ)������[��V7b�Ɗ�J~��Ϳ��/��"�?��P�n)n��T�qb�?wn�\��]>^^Q��?<���$�B�3�S���;d�W��Zd�F{�{+�e�^^�8���o�\�@\�v��7)��jC�ߕ��@��|K�F;'�\��i%\�d.���g��������I>(�3.�F������n���lEWn��3v��$���������!���t�1!�[{M�-[lIe8#DK=a��'~46b{ɾq(�͠��IUл�7[�ҽ*3�R����(��*E�o�$�d�x��'��j"�'�7��`M�U%�j�����ϛ?��Σ`7�_B,kz�4]�X��@7��Ex �SҒ���5��l�w���o1$)��p�@Rĸ+���ļE|���N��q0���R��C�&X�Oe���X����0b��Fɩ���L�%O����0Ǻ<,?��
 a׭��~�96Qf�'�h��%��R����%Km���N�%q8+	��AU���31g�n|	�mf�//��S�h�����z�ͨ�+������'����,����|mv�X����@@� ̈́����"_܍�aa�!�#�Р4Pp�����V�m��O�5C��!����g/׈\4'������S,��q3_��L�WI�R�&��tӍ9T!�G|8#�aŔ2E>�Z�F��Uc�{��^A�SB�ݍ3�9���tpkF�ь��*0�[�\�䖹1^�՜_���q�D�]�Y��&�j�[G�N�����[]�0�ɫn�~:p���F�1j��~	�L_v�և��O5����65�Й'�0e�@$��:xB&��B���Moeuh�[�r2}T=J�*~�V~��l�B�ǹ|�7��
�� A�������,ڿ{��1S/J�謊g:dج����S��e�p���Б$�<��w%}=0]Eѹ�23�y�x	��� L��rY�[���yB;*��l�x���C��	�7C�:��,5�7�D��qw y����ŰK�"�-��wßC��#7���?(t�7:��C������C6'�G~w$���ա�g�{�����:����NȢѹ����X�n�X���Y��i�5�pQ�-؍Ã�K�j+K��'�4dg?U�3.���@~�"��؅@g&��_� "*8^��び�;�S=�ޥj`A�gbt�KP@�DL̷�gEr�:Dz��Gų�ӲcEe��}C�!���m��� \�6l�^����	�l�CDa��}�H���;�X�� Í����#��:f9�/�#���5��rD��������a���3���FP���u�Z%9�q�Ũ�'��	,Iqa�֙H��;����qL�ycn��w5#����Y�����Bz�S<m��w�CmF��Rp���dRM�.���"���p&��rm�5����s��j�g��/,�!���m�g$�y�.-��,��?
�I�D��>hL���z+�ՓD{&�ٯ���S�P0XA���V�������o?��&'��J	ҫ�K��Z��<n˜�?*���C5�t�k��[t��o��%�]�3�7�a�ž���g^��L`'�m0���<W��Kw-Hji�%��o$p�T� !\��An��UQDu܈���������:Qƚ{���ؓ��e/�O��gz�J�Mm��(?�##���5��ޏ2�W�W�X��������2K @�{����>Oe�$c���3r�����1���ҧj�G>�����f��(�	#=�FdD؎��-0�X0��6Í��v���h���! �S�4�v���	��|M/�A@��I1	�]��|��!�CdcsM^�s2�&�����ZL�(�4X����bZ0xO�B��U��*�3���S�4˦�GIa�_� Բqa�ц�=�R'	H������β���q�$�L��HH��s�v�1Ӧ�ߪ�3>6��Uf�"��X�E�u��'��N�{��p��l!с?�PV)-
"|˹��)q�T/Ë͠EOaLLY�;EeI�XV��L8�er���$�Ҵ��b��O��
cʻ<D>�5��r��_�޾'�/:F �U��J큺' �y�_�|#q�a��]�zp+c���0�D�8	��,��Z���? H������ ǈ��ٚ���9N~!�|d[H���4��uQ�:r��+���.�>6e��ƥz���ձܩ�6��-�9�?3"��
��[�YI-=5�P:�r��Y�j2�.�'D��]#k�ZH�b�I� >/%�'`��ĐʯL�ش���q9J#�I�.QX ֞�Fm�dy�8M��C��� �!��x,"jG�L��C�f��4��ഈ��5��6�%���R�p���x�����E�|�J�*���;��d�9 |!�f���_=�T�4ĈblƓ΁fP�]	�˿:�d���
��nS��ٌ�71}�d=f;F'/E����j]�~�.{�G�>�I?_hF�R�R:���\Χx �vi��LR�UaJ֤у�#hO�2~��)�/�T�Ԛ�Wm����U�-�B% ��^�I�r�]F����Hv����I�!{ykw*����m��1�������	�)gA�2-���=g'��KPv�xep�A��xӉ�k�~&
4n���d�*���M�J�O�������);vL�/����DV|�}/�	z�n60� K�m�$���{������g����U��_��d��@쀒j!���U� ^`�*�������q����Qz<��5�S����?i84S5��=�p0[k�(���Ua�d=s�C������Ê�>���l�X��82��=�9r�~l?��v�W˛?���/D���qҡj�� r���@w�v����;~+'\g�8�}N��A+<	�k�Tr%]���~6�ߖ�4XI�^>l�p��ڃ���B�[M��I��x��*<5�*�j���71�7���4EBe�q]E�e�Dֶ,��(7B�}���|������?�5"��Cf�IZ�ئN�STD�Nf�J\�����ӛ{�B"�� ]묐Ե�4X�$%	)��������)��M`x�f'P��Uo5�0�6��&�u��9bȹE��T�|��9zz5+=�<��:��KQ��}MPC�G)�_��ɂ_�s�}�L�q��H��6Ƀ�j�j���<�&)_��Y�a�0�qd`�2��C�ݱ�l8.���]�,P�UT�l;(�
��ղK�����V&=̛@2��_�i�4��lA��ÈY+�?a�v����kϭC[���sQyȳ!5��iL�e
�܃?rxO�P��_=��P��Ɠ��0�1�vH+ƿ�3Ѥ�X|m��{1��j��J�%*�Z�(r�Q��'l.�U���p��`���v��z� �dT�c�ǽ~9�|�\7���Y������8]FB��h��tf�� 9���P��}c����4���mĖ蛼������{��9s��P�Q����\��)`6Ӑ�{8f�6��`�=C�KB�&�Ì�M|�m�'T��mx�Ӯ8M�.�ͫ�����D����'���bM�!�-�3�CTL������WF����?5~��S��kjۂ�6�!���d���B�&�gត7�5��^����-��.���T�V��@2Z�}�x!��5���k˲����S>U�;��˨�o�_��ࣝ|��n�K��$v  ��I�k�cmS5E!<�Җ���Cugz='��?����~�����o�W���xς���G^�H�j溸)ppS|�BMDBh���">T ��O�X]�����s��<؃�L$���p�x����p��~�L;i�&�z�6�`�&�4`¶͙/,T'/e��y��@U���Y��i���ǣ^� N4���"w`�	��t�R�/�������_9zK0Q ؾs]�}�CD��B�c��V�v�~ 21�e��IPB����
��������ZHҾ�.*r�\H`����|T�og��=U�m�W2�� M��I�;�>H�)4D�߸�˭܇Vj�1@7WT����C�\x����A �?:irz1��o}	���;O_(�+�2�٥D�Ȇ�̾�8�~�7R�S�:8c�I)�"+�e��QE�If�ī����<f �r�s��f�_pN�I{4 �CJIi����i.��c���to��i�)���=h8��4ZJ6�Z�S"p�NX+b��v�;����k�����r����*��f��ab�Q[-��aw�:��R�0F���e�����Y���_�,םVܽ߀���e�K�O���3�wˏ{�-,n��B��Kr�,;Vb
[?'=��LeP��a5�q6�]�6��ٽY���f�H�q�K��u�^s(GѼ;}Ȍ��$��Tb�/��?h< ��]������t�\��i��sd�gM�/9����AxĘ�]�^��`@�sX��K��hX=w<l��/8o���/�b ��b��
�D����)աӚ~Qd��!w�����/^w̻۳��>�CX�p�=�XN����s���	#�{3�U�E��b�l|�"�圣 �lHK�����X��%��.I��.��iU�M��`�w�C3��8g��y���[���R��A���5b�ыi�`$}�u��L��2��y /*�0N�RMy.?7)=�����h�L��j�~�u�8�Gz��Oek���I�p�[��ԍ�/�&�K/�Y@�~��D
2�a*�����c�~wĈ�#���q����l^���(u�9��H /�6��Z��󿰾\��Y��<��;�����#]TM�UҞ2+b�;$���ƙ�����."��K���./X��TAs���3�j^�s���ՃZ�B�n��kR�\�(��f��.2n�����jb�b1D��_�0�A�ܓ��
L��#r%xR �d��K<ڎ��υ1r�%Q˯k#��0`T���,��L�����F8�Uh�DMD!*�O�oj����E�Oy�� �4
��[���'�qe�cDc��OHՂ�b�j ��~aD�Wzm�h;��Ǣ�
Ƥ����ԞH�: ��y��yqs�g\(�� տ7�޽�c�~�ӆ��4sd���k_��p� gP3�	D�a���q�W���=1��ԼTx����׌�X>���P�I��ȏo���|!˒��bp�wb����.�n�D��?����,�4���<�0�.t�:5P~׸&�#Y�ds<���R�d�^0U܃Půc�/	'���s���ї��� i:��xW�R邼^��4�t� 6��i-<q!��Y��+C�!��H��l���q#4�ިٞǂ9n���nT�w��	*�B�uBepy���I�m�h��0���ȝ��z���׀/fڛ�kA��{��BUI3eԝqO8��r�\_���}��D��'�&�b��HJˈ(����r���Mq��qe�T�H>H�$���8&��֢�+����6�[��(5����/�Sp��*�Qx�'+�|I��%��@l6�Pڰ�,�z�U��t�b��X��ŧ��A7�ʚ~���6*uh�.�7&��
ZK�wp{!%Bv�8���P@}�����k�� y'VY�r_�`��E�i[�zQ	h~u�BM�7���c�6��q����?bG�"FVpu�o�fܪ�Fg"���XO4?\ц�p�R|J�������D�ϴ,�Bk�.X�t��?�cY�Rm����L��P�0]G$�@3��q4�D~'�3(���v:��i�_ɤ���\�+��T�ư��hO���PV������L+(��9>��ǜ-B�{�M�F�E���+,c�>��eBd����Y�[����>����D��x��;��0����p�9obK���i6p�ʟ��5Aї(x#I~������'�;�  �*��cNGr*���K��}f��VV�MV�����B��)�K����7,��ʫ�>��˯M�,I��F%B�����f4�f퉥���:>7�T�@��ok*�V� �F���H�c�oLn�#N�5�0/��>���_v����/�nmoI��)
_<�/��7TN�&fjj��Y�T��}9RZ������#�*>d�i
�^�Ό�t�æ�$kK����>,�o�\�Y�M[��C+�[����c�y����r��8�Jv"���+����-6�$�u��W���,:7`�]�	�H�;Ȑ����qk�| �0��a������.��4M�V��i�����%�vvl9]�mB}��o�Ϩ��w}�-��b�\a�<$'�>H���s(��N�S��.@~�1��>�q����A�^m��HB�/�
��[�jG[Ek��~V�{L_��[��+�F�0ˑL�8C�n�U*��w��nsq�|W/  a!ԩ�Y�x��k�nſ!Z���U��ߥ��+�l�)��~<ɷ�vJ��qI��u��
�>*D��	)����p����F�A	��$�9�$̼�m���˖5��m�c[����p};3�W������
R�M��'=0��܀��ɔ��i�_�Ba^yz�y�3�O4_t[X"�G��͒)O�����( 8x��_� Ch|Y*�G���ܽ��L��p�gr�Z?@GQ� `'�j(��ylK�:hO��_��B-���h���C���{�M��2��f� �	 +M��T�	x�[�u�BjCԐ�k聊�;������j'�}� �t���
�b;m��R�ꗼ`H�)��,,�����Z_]!Z��.���E�ƚ�p%���(:�6�1<m��آ��|��MM�����>���7i��l�7�v��u�ϛ]�I�"�cr4�"v%ˋ�<<I��4�^���_Bz�q��{�AN5VMúA��uW�`�/E߅ø����I'Xngdش�sc̚�/@��׶�
��)r������-���}�BK���}��&g`��	��%2{T=Q\�KnQ����St�/'�gx����nv���Ra{�zw+�1�{��H�����|L@
J�#�ё-����e9�z0�!�x�f�.[!8�'��%��+x�1qx�҇��7f
D�y _�*}p�6���3ͧH����-�m���DQxP�o�kNoh���>I{�U����1�F��72�y��!�6���v�ܲ��i�(Ssg�T"�~�3Sn�%t���\��|��9�;`��^�GI��I ٲ�ߕ��y�1s$ҹ[�9�ˁmm
���2\C�~r�6����K���W�k{�(S���Z���PԳFP�^@�E~�i�@�|;g�>.8��U�x,���Fm�.�7����&Ueln�p�;.���T!�?� !g�~��d�#KS]���ln�ENd���j�V�5�f�s:<��d�*���gWN'0����˯�����ԭ��4k~�ׄ-�Bz&
�V�ϲ���[g�^+O:� B�������@����T���x���_? #� ���n�DuJ��35���[8�Ha#&����d��6V�n���k�wp����o�x��1r�_F�v��pwE�����Vxx,T�J���-�}����c�x-{��+(W{z\��y��(˛
�%I-�3*��J��-$x�9dE�GM�Y��e�g"�BϺU��4r�I�!�r6�Ȥ�� ��)���*�(N�%Y.9��J6��y�}�Sݿ#{�r�X�ڊw�!�x��-�\'�yϣh5��c��2�mYe
��ym, �JA�A�4h �ƕ��B��=��:��u��2��x�:��~!G�ǆo�9�N����r�6\Z �,�Z|}Tt�� h�hQ��Z�A�V;�ٺ	���誦2U �t"�Ќ'���^!�d���O��j1���C3���<VS$a���~�]�@��D*���'  ��eF�6m���V���9���nj���p�L�QAP��{?�1{�%����ڶm�C����]]��_t��d^U�AS;2T84m�:M�=�_�M�D=uNcP�Ʒ:<��o�����&N�A1{���G�DQ������%2v�����?%��;SDSdMJ%���A�^��c#[/My���y�/f+��^���ҏ���l�Tj���4�C�F/L5��!�WƆ&�{�h_�;���:r�v���o�a�Yc��ùW��_�,�������F�ZT��QC�`+���"�&Wsrq�z�jI��%�9GD��	|N ճ1j�&Aˏ �~ur�L�k.�W���Cn^�5F����_û�4���2�Ы��Zߓ`z���
\N��r��m��� v۰�{>V�-��9L��v'Cq�夗�+h/�^j;r7��x
�&�_s�VM��+�F����8�E�l��h��&pǺ���.��f��v����^Â�Y.�%�]x�C'|�Zg�O�Zȩ�K�lܳ���کE�ͥ����&��,*B�D���%L�5���7�YV	��~��?7����t�?7V�.!���ސ��\C%�9�N��dV����\tDG�{y(ɣ���C�[Z�����3�,3���ӻ܀�Oi$5���;��d�W%��D��=�U���js���*T_,%_�0��Y���(Ā9���R���}�}
�t3��\J��Q�4۬)�z`��Z��������҇����3�'��ж�ǡ5ԅ�9p�:�D�tN
L��Kt?��5�+<�>��5�w���n�QT�x���(�%㾝s�ҡ�m���ur;��C�V�{e����%b|m�Uf&����'��CbNKԧ�iw�<�3�k������?Q<�s�{1�=�#M�.h�a!�)_N��F��4���,�3����A�,v^��#G�C~�E�S�'���bMl����5T�ܺ?D�2`�adT��)V�	^��(�ѳq�ߨ�]$���N� |�I��&� ���^�w����([K�5�MU�g��h�`/[�/yK��V�`H�����)�/1B�t�,��s�Yfz�����j�Lиš�٩-���h0�s��@dS�}���mU6W�zT,���b�kϪ�t� Kҿ$yc����j�p弍;Wr�JH.Esb��6�
-���v罠[�u�*�E������a�3�n�.
~�6-���������e:���ɁϞ��+�v�-�So�J���8c�V�4�Hf���o�<����{��#VF,�c�n�f�J�?j&~��a��N+��t]����>���A����}�)%�VJ&�ci��U��h����t*�w]��T�2^��3��?�Q��^u7��fTZ[gy�%a� >����]�$E=9Gwq����mbҡ{��Ys��`h�a�zWԽ��/g*���Sϳ��nS�;u���5�Ӄ�\�{��8ii`� KްB��Wj�0�g������z����l������=�����}�K���`���2I�߸�ӱNAm$z}�X����R�cc���׻�a�{6����5T��n����ĵ
dέ�����+l�������4�=K�,�~??t6���h�^�}������� �XB���7p}�5n�+S�ABǞt�����_+�k!k���>�/ %I�j������ ��@���A�Z9������my8��kې����)��ƴ}��A�}cG{���n���'��Y��rU�	�ev��ﺐso[np�B{�~�к��'�V�	1`
����x��h�.=�K�iR�����:2@���a�$���@��)��r��k\
	(>� �?ԇ69�OA*6�O��W���t.`���ư\\��W4���U}�Zf6d���epЄ��m���$#е+|�Z<�:^ý�I�xr2�k��ִ� e�`��`4T#b`؆��f�#������|���^��7�pl�VFn
"�¸L���A�IG��I�cW�B��\tTym�	���8�4e=����0�a�
���du�)W��x����~� r�_��;�Ō�)��#Y-f"=C�y��T�'0(O����ۚͽ�K^�B��F���{h7��Y
CxH��q�`��V�㍸�nM��0Gm<��@kX��\�h�G�{Qx��B�ԯ��L������6�@��I�)�a�=�o��4��"�g3��L�M�pb:.O��?�����,rb�[p �{����ei��}�}k���E#�Zz����*|�� K&C��W������1�rb=�=�&r�T�[ާ����ȳ������M�B�NR ��`�m��J�;�y[W�"Yby�s�@�XZ:��yɅ��c�5/�~��:�b�-��EI�M����M��<�6V;�B�
s��]�,�x��t�
U�Xx��݄��O:�ZMN¤sp��	M���_U�
��p��8~u��?|($��c��kP�w�E��n/��?�1cK�U�Q�P\`�	oB��ufe�̤���렏|�� ��,���i;����a(�)$��7�fV�L�G�L�~� 5A^�}
�M�	+������B��gT��N��;����WA`n�� �r01���f<ӈ����Qvp�B��ۤ�i-�6�j��0���{�ۯ����1�?���ig�O� �ሽ�J�6����X���#��
z��u���j(���g���]kV|�G1޳����eQo� ��DԱk,�dD�ca�:B�0�t����ʴ���h��$RD5o��]�5U����
��"�/ř���)} �����28G{��P�6�oF���K{�Nɵ�B؅������0W{!	j�;xPׁuZ Zw���	�k����;sZ0b�3J\�Cb�E��?'<$��t��)�(9�U�"�D�\�s-�M�a�Ө�h�B���S����Մ�}˗�࠘�p9_kmb�0�N�`Ŷ�����36O�rsqr��K��И�NF��|�SN��IKe��%ɏJ������o�`+��!�(����E�D�U~n6]y�pm`;I�jv���o��*<S�����[��@��s���`�dї�m�8�����$N�����=�;J�ˬM^t|L"ۊх��3jP��ݝ��G�'�Yly[��rc��#�Η��c�X��#-�ͫ��#_��!,�]�=��v9a�(`����Z6�i��j]t(#�k��3��0U;揲�&�#�'io!��h���J�2w�!������Y���~�cCJL ��gV�0@�G����xBB��P�?Q�~�����bBpd���tVؖ����Y�\ϋ��W�;"���UeS���P���N~�[ �eb�@�Φ��E�-Sh0���J@�rA�3�W g��$zϔ��!���9���i�Ğ����WO%���3%�Q��P*s]���ђ���X@.���إ���>N! �y`�B�!��=�7'W����"����K7iQ�hJz:�������й�?��ndz@�N?MJ*��_0ei���*�����W:���щdPm?���S����$FL�
fs=�q��X���u�s'�iL���G�(�*[#{� P���T!Ω�v�U�Iz
�+�գ�F�&�9�'��1�Cǋ��{�T��H��e�Cf�0����_�?����Q�އ���9E��ޫ��<Oi�!�6�ڪ�\?݋�Oh�Dd?^.{�Uoe�6o9lm�GvE� ��$���C������bQ���ݷyK�H3,[ک���J���o��XY����C���p2Gd��gj#G���~�� O���	2�V�ט����&�����>��d��J��Q6P�´��H��X�",�>ۆ�}u��+�����_�n��뻎
�τܸ�(�6Fa�|�t�sRG(9~돖�7����H\�n��+��%-���But@��*N�����!AVڏ& j;/�nx��� S�ɱ/�����x{h	������s��7��b�J�d謅�a��^LeO}���+�~n�{q>�Dp��	%T|}e!��2"�pY���A�q�'E���:����Qn�>���xd6�0���*�n�t�@6���0+��H~o�-S���%�X6��^��K���i����>�MU���j�J�h�:k�׾���JIE��K�<}��� �N���|tX`���D�R
aT�W-y.7p�u�,""(�%4�iض}��5���p�[�"����h@hZ*!���|
v.��@zvz�p1��9+$W�Z��y�_n5�P쬰���Z0�VB�Jv��ؤ��C0�9��VF��F�V��zIL֚Z��nO����{��NGi��[S������6���d"d�=;���X�%7���D&���9��3�5���=~����8:S?���-]��=�0��c"�t�@H����H�]�1�o� �,�����$�.> < K�n�/�p/X�Nx���C����a���������f�i���A��-�-���ӛY�9+-'>�̈Z-�TvY���2���A��8���f�1j�S�CS)�\#���.>"O�@�U���:�I,�ӝZH�4/�PW`��-��,�E�u��^5�"���X��Qp�*��u>W�F�e�c4sѵ��1yu��{GO��8Ne���~���[�Y���I �O?���D�G�ޓM�-MĎN0:�t��=��&�2|���������f+�Q�"�=u���<�����h��_���,��O.��0�up>�8ہ�_r�[��T�u��S��?#��V27O[���@i����2>~��ί�C2@;n�<i��^ve#��އ�ѱ���C�C��u���߯w�E<%��ti�
t��b~^0Z�q�"���L�J��lπt�d��-��j�E�E/TfU.�_�zx<��f���];�5Ǐ{�U4~(3��yQ��W8�(5E. O� �n���4,�l0ȥ.X%�$5�c��Y{n,���/�f��-����6;�^pS��'@����� X]�-E~��AT����������%Q����,�I���C��
��ݒ���k�c5#V>>�ّ�`$���%��^\z���C���Ť����i�>6���L:6W2Zs��n{bw?6�Ad8�⍆�Wi��^�����T;����x���n�e%;�nO*���5�i�����nS&H���?L��Y��?	�ڧEu�GJ��R��W��t�Ξ�~�#��z�ڐ��Yy%d�y����C����8�ό�Y�t��՘֑�eD.8~��n�;���h�CQ��.돔L�=w��?��cì�	6�@V��
#�h+%����n�@M�R�[�t�]������%�Xa-�Q=cꃠ��a��h�O}�pr��� |�Q#wIz�~VP����PM��I���پ�1�}��hVO����*��
;"(BZ�x%N�5��KR�
��#w��/�W�r�v)�����+���@]�����x� ?A�2-��^LR�p�#}̯q�_�`�'��E��$L��ͽ�#V��=E*��8M�@�;h�%:N��lx{Fz8)4j?�>��	��pIx���O�-��V�.�A]S>Å�i��{z�.8�9k5JU� rX�ӏ��f�����} ��""[_꟦�8I�*N��&�6;�'H�������x�&<Z��Z�Y�^�;%��Ӟ��s�@Hs�I�����$�����m�rO��ɀy�(D��_m�7�U��Ns��M+/�i�C��G#�uaí'��>t6�U(�OhT�ufC�3����Jy2ݢQq����$%��́��H��6s�(��<Qz�� F�>	��f_H�8vf�ҩ� �()&���;Z�nc�f�/kI�&��G���2|uR���Y݃��],ٮ��a�,rz�g:������kg�a�����!&�����d�:�R��v���0�G|�ȕ�T�5F�����	�c�)$W�^��v.��^ی�X�TbaT���{f�%�A�Iw��ƕ�d���Ev�6�{g�	�����Ж@.������:��6 7,�H�.;����#¦ʡӹڈ( W"�T��D^����K~|z߰���W�(���Zg`(�B�H�y���t#ƢL>��i��C�U����DK�f��	 ��˨סSF���~�6�b3&�W�q<�A�s�;��NW�IB������o�/쀏�Z���|īʘ.��j9v�9�x�n'n=�J�ZW��'�Sx�@��
����	��B)� _q����~��J��{b�ũ:�].Le������>�w��K}�����O(]�{���Z=��Д�,8�ު�:h� �r���,����S��[Ш��@-�^�9�4a� �oz�l���z����)�ӣ�#W��ܬ"J
YQ��d��Q� 	�(�J�J��[��>z3X�dUW��ol�#�������|�	�$�����s',Ra���N���9=N���&�o��3��G�+$�Ѽ���L.��)�#��d���{��!|8�k�jzGk�n�Nq��z�-Q_֣H?;d�@�i��h��}ļƨ�NL��VjA#W��N�hlWX�^��{6�%�m�م��T	�%bC���=5F���D������`��p}�Ӻ�Q�m�8bN
�ŕrl�<��F�4(fO���/���ۈ8x�ԇ6����nւ%�j���Ȓ�^6	F�H�O�VO)�1�klP �e���dfE���v���m�"�����}<�ɋ-���2��.��������k�;�~<�����%d��t�]6�7x�����<���D���xr�5��9$߀�	=�v)�-R��ߘ&u�,˄���<(fbS�j���u��x�3���n`9�-n���$��b��	"����K��[ݖ/��8^��E$�@ךV���|��א�BA����t2͡*ɶ��<�YP�V���N����\�T+��n6����">�.!!��G��O�΅�)C���
)��qC���_Wc��u��c_ɤ��n��z��c�Tvg�2jeW��+-����TTF�'f�X�#�-���橥�zzZZ(�߂��ǝd����CzA.2�(���tf�#[�Wu�8����rv�k'!�-d�;�L��Pk_8J'��������y>�bh��*j�� -��d<��&ˀ���u�tj�p�u��=Y@�BӸ�TK��e�$�RbL������$�V$E�fh��@Gʔ�7���D�v���\Fu@�R_��2�h'���1=��f6�8ߵd��k�r��X�Tc*LB�b}tD��"�Y���|��q{�U���l�I�=7�U=�����u7J:1��VX�©A�(�l�x�_fe]�Hh��=it�����#��݌ܔ���Yq�+�m{���O�*�/����+����fZ��0����ߞ�?�T�|���d�7 �w������
��pDf�Q�=�������<BC��{��w����Z�&�P�y����J>�3��\�4�<n�u�D���x�x|�2`��y�������;�ZU�l��A�Y���B��q3%Fр�o]qGN����q9˳�`{	"J�i�K�D�Z�َ�l;n��K=��{&*�(B2�W����R'b���8�ſT�ξߗ�rиL�i�N\�����խ��Q���Q�#�Z�V�qZG����c<�nw�wK.���v��7 ui� ��P��̱}�4��[��o��ĸ~�T�_�hJC;%�Ns��j��R�"�E��$Q���KA��0�ş:����+��$p.]�	���+�+@��аy���߬}%��;��v�1=����W]���N[��Gu�8�Pn�Y�'�+G�p5�*��
����,�o���:��?^g\!E__R)�t��+ڌv�y�b�F�6��Y΁Q�ғ�/���ߨt Z.�B7IaYd� ��2���f#�6敀]���'7����7�T��m5+���&���))0��W Ϯ{s�J�,:r�rãy^;�
@t"
F��$���'%�� 6G�+�(}5&���M��@a�(V]e&��>q�Dӧ�𓈻H�wU��v9����1bk,׶U1�o�"��vs�X̟_$7+�=��p*�ƈ��=p�	��[F��|�ph�GZ�LX��c^�a#�����\+u�Ლ��2�,o˵_U퉊�4��*셔��]r�����i��8#y�����m,b�ut��$�;�di��.����ް}AKb��-�/�Hs/mN���Ӓ<F����	`.n)�����܍���Ar��h�k$�ƔyGy��Ŕ���A��ܱ���HfFB8{)���7�o Cc6����шG阀v���p��G���w<�zJ�bol��Z����U ؝C�o*##��2->>���ؕ�e܌�o\��gld�a^��+Kn��۝�m��o�%#�-I�A�,�Q: :q@g �¯�K��UivSjq�N����KG�g	*�$n#ihf�8�w�Z[���E�a�����c&��������*[)jI��*#�쮕�[�'�\�8>Wxm�'�8aρ�3���3J�2<+v��VЈ���U�[��P9V�e��|�N�|�d.\n��mYf����$��[��+>v��'���B�܀��C��V����� ^�CE������EE�Z���]0�s[;&Z��ϣ0<�_�
U����0�]=�ע���π`�[ �]7lr�*�)<�j� �И�+Kv_j���e�/�se~��'�^�`k��e6�e���oy�JK�+|WAH_�8���}��d;[~�1r"of>A�۟B���ؼ3��bԌg�У��Wۛ+�O]B2P�Us��h�w�y�.��v�X�w��S��%��-M�d�u�P~�������.Z������$HZ�amL��9yveX���>�İHY��6���s���n(F��$��<|����oZ�Y}�~��ǚt�vz�°B�9.O�}�I�������^�W2 �5���1����L`�,;g��Ϝ���s �����b�i�����=�(��Au��@�����aO���j�`�\�r�f{�hQ���PJ\�l0P���P�<G����4��z��4���y�Wӕ�u3v��2��	<*�˓17*���u�
��o�����6���Q&ݔ�FWߕ�U��Z�����౼�O�'qU��8��m�>�٘���0"���6�0󡟷���o-�Hc&\��䂟�M����U�:+tTax^%���Zt��'�}�跣�}�-&�P�2Xpi���j0�렝�2m�R�[�����@A�q7&O)�3}�}��Sq���8Y-��b�;��D����}��Ib��x"H׮9�������~��{g�@�9���p���l���C�RP��0����|�Y��fC�Þ�-��m.d��⊐�q��������81p*]�����l�������挡��.���עnQe�O�f�ڲܐ�B@	n�'44˙�4,���7]])�wU�\�"A=��t�,V�����{w@���	�f͕-��	���.���4��GX
��+��D���Vy*x�i��1�7C7��q�kS%u"�BH[�:�ǿ5�|(:GPk��ik����AZṠ�I�]���F3$G��̈�Z����0sAw�a�ɬ�gI"�*Fr��
�K�=��p)���6Ef���q�* �~Ѡ/�3i0�d#ǂ7�`�w�7�]^_*��/Z����:������-n�h�����2\�-��\�!��s9��}�-l�?�X��8/�Q�F��_Ax.fq�� �Z�,�$H�t28 ��O�yzvfb��N�n\��	e��)P�$��8e�:K��N��X���[�3��7�"���y��'Q頻n���;��(��ӥ.�4��B=t?�z�ϒ�0��Q�0�*^eB:�0v�D�w"�US�r���@��5�ڎb���Z�l�����0���z� C����ծKe�S+�+�����-v�η�D����Yx��%�oЌ��� ��d�F@M��C4�ԇ�hg(�Gw{��U�.��-l̺�;Kj�VʹXͣS4^��%��h������j��H��7�\�LNM,��0e�\��D(@ ˈ:;ek�r��wI��)XmMys,�;VPqC�b�ɂOv��0�C+��m�ڽj ��"9Ȇ^�6�ajS30�Iϻ}�$��J��T�L3J��H[=�j���%xNG���b	��~�T�73F��.E�炽���]�/YE~�=T��X7 �E+ �I��h;�^u~���N�Y���& �uD��4���ܬE�r�b���F�d������I���b��`�ӆ����$u��ֺC��UT������	�>uBumr9Ӛx����Q��S�#�O��V��v�Uq��9hH�lT�5�O���ġ�j}�2K�b�5�rf:��@6mq5J4��` -$��xm)�(��ř��{�|�(�%ﻬįd���������f= /�\f�_?F�������Z�����1�󶍤\���q>�����U�e��
%*��S'\��xa���~=ّ��1�P�w9�
<%"���"�?�9�;K3g��%=�='Q�y��
S��
�]�o��fWY�*���K�Ly�[4�ϸ���?֋,,J�\��(E#0�2��Al��$+k*�%[�G�Y��agqI��2EA?���,<��i����U��a|��f�oۧ�Q6,lA=)��P��zC�䚵�1��u�ɖ8�>锵���9����9w]���55yÓ;�+t����%8hoXb�B�2χ�"t��]�;�����G|K~s"o���Kv8N��1U��X�u.#gg0�� ���k# 7���n��I.��U��& ;t'�����������'Cb�� J�� 8~�p��۔��Hp��d���a�Hg����vq�$n�t�O?eW��B������]��zF�+J�`��՜k	���`̸�Ĺ��K4(�y��WΔ{��3\���%��W��;���5�C�IZ�՗(>�������gϷsڃ�F��_��VL>2��\�<"�l'G8�$�J��g�Nݙ�����-��2Ƞ7&��$��t�����8y�2)�?	g�b�w�Іd��#���pr��>Y}�8�QDw~w�O�s��]�*�uO��e��3��6"�����D�8� �w~j��6�k� ��
�N@TE]��}u/3WMs�i�ۤ���T�/9�ԉ�������rޑd(L��¢���k�7�k�dtMh�h��AԹ�JJ��3#
�m�r����H>1cV�R�܌�Mj�1�^؂f��ށ[$����@{��k����$c ���� ��|�<�狿��C8�D��L���񍽥�)��,�D�:��dn�K��,p��Mş|��]��yp�p��9�J԰�h�M)�N)�H������"��b�!
Tމ�9m��F�z���N��q��Sl�a _F̸]c�s6�Mac�%FZ2|��3��}k!�ڶ��ֵ���h��j/`c��\��U�(d��O�BԙZ�:P���i�<�9K��H�7��<���尫@�=�Vv[h#�oA:�g�^����u���Kj�?�1'wf���r�yb��`��IE�U�)3,䂵�����6�
��/H%�G�����\�A;�|N�| ��� �yO��'}���6�yYl�?��ti����ڳ��z!��k�`�)o/p?��탛�ǳ�T�x��:����nA�F��:*w��+����h*�	���3Ln�u9�����Q�	��f�]��s�]� q����ڬ�@��gohE���־Z��RF���9~Ĥ썟{�t����g��ss������!��-�I�R�F�wA�X0}���\����&�0�����<�! �0�߭��h�ƙ�|6�%�u>^9ۄ���ڹ��`�svE�Γ-Eq��<H�����3�Nz�%C4���|��!�4�D���%t�f*@�W�,����C�NE tIn�.M�i���G�M��	��;
mORv�:G��շ�&�)^��cV�$����� �� ���e{Tr�24��QgBcyQiz���^ߥ�e��Z�x@f�<�F���1@�>.������G����w1��l5�1�Wd��@u�+��_
�4a|�����W��c�0�h}J�O�	ê _h���/���U�;��_9��p� �*���Lk��z-V��q6�������w�Z���a�h�QGW� bB@�y���7��(q�8:+"`�c� 63��,�&�d�.���ȕ����0%���Y�mWD����[��H���Y.�4w�蜛���5���j��ʊ�-��>:�m������} �b�Ϻ��6�H��*�`�$5���e���� 4݊B�!���\��H.hrɲ��Uh�Q�Z
u ��í�- W�t��;�򙦩�6�z7�����7�Þ/� ��{���Z�Q�T]W��6�P����%͉�[�$D�m�RZ2���0-�
Mc�>��^$T�V<�1�dj���5H��E0	���.8>�ڭ8_0|�����d9�����ֆ����^�ؖkd���7�c���"ބg�<.�3��T*�q�E�n��Xˣ?��0�f���Y�!-|Y	��*�6�&Q@�,k���ꧨ�w��jL�CVw�i\�.&�۟N	��d�s	�|��	lr���ʹ�׼`Zρ�G��@����nم�i�Q�4i�F<�6�G�-u����1.R�J��BtF�6�S\;}|���4E�c2[��~E��=�YL/)ǽ[i�g�1�Nox�(��u�:H�Z�ZQ������TI~�7�$�;��I��m�X��2~��il�y܇���Lq����/f;��U�M��-����1kȸnD%e|C΁nn�ov�ޜ���W��_BСJr"��lᚲ[_���#��Ǽ�dU�h,�n��b�/�r/?ɉZN����h�r���,uj��	��v��K$^:Jٟh��5z�7���y��Lu>� ��b��ZuY�H@��L�;>���i���DS[/Cg�g�c#u��[�o{�j��4W.��o%�-���̆�Mw�we���D���~>^
E6\ Q~��`���n�K�P��=�\L24�[&�������u�|ϻ��i�K�O����^�1L�-R�WY�_6�����i3Y��y�
1[�w�3����v�h��_aZB�~�|�J��15��I��F�*�V��>���C��2/ڏE�[g#.���ыb�t��)��
��Zu�5����;=���m�����T�; R|At�0�=������K][ A���p���hK(�S�Tx��A$hϫݝ�Z�V����?�L��S�d���5���T���9�	J�s�����0�@�p2���&P#6�V�А�����7򊹮q�& �����1�7!��|y�)�_��%�t
7_NH=A�r{xo�>��`p�%�N��KYW���	й��������Tuc�̐�41� ��)s������$s��P]�@h�kGw-���Rt�⛦�p���3�%l���,W��qݲ2C����̬�55�� B&'@�|е@@��OS��Uu	�H��ĜЏAf�oQ�`��P��#^ ]��	~2ל@1;�0R���%����f�ohq4gT�7���}r�������b�8��M ��:^/�Y꿼s�F��S���t�:� �6����W�*�6V��%�^a�T+j[�R*��T�?]�3�����9T��G^C�������������/kqx�8!�a&�)��j��-�-ۓ>�F̅�Ad�4xmR@�Ĥ xҨ�qj3]��a�1�(�R��=�1�~6�FZ��� ��a�TE�@�weU�U^�f{��8J�8�V��S�P�ji󥿊����$����W����0��|�Jע4;���m3# ����P8"�IDRwM.S*�Θ+��B���!MM�%߃%xK ���3�k^g*���W�l�q0j�i��WD��s��8'@u����9*7�=�3��-����a��2�'�%���V�M�΍��5��|��i�J�z-1�w����:y�.�mX��ޏ�P|a�12�U����L�n���+�S�T���e8�;K|s��{����Є/��d��JT�,.�m���Щ��3�Jg�\��4Õ�A��83#<�v��ؾ�M4�������t��y��3H.��t,h?X�0y� �ꁹѿ-�+�>��_�w���x�-4�!���hi8a�sR�'����C�	Y �}���B�c	C`7L͕�wku�LjS��F�=��7���i�� �7�zFu^�- {�YI��j�77Ab!��vx�3ur�Io|v�2b��l!��	$��SN�̨L��oQ�4����=/"���G�9��%�~�U�=��&�i��bնxy�vyV
�e����=͕�����-�۪��@霶��8,vZ����`��ǝXۮ��3�s^���t�*1j��(R�`q �B�l�ڹ�A��U+J1�.E?*�O\�P�`�C�]qb!�&�!Ĵ:r�b�Ǆ�:�&�~5��e'8%v��{�z��L�p8W\Q�G��P�y�)%b�.x!c_�)�2,�B��E���y�6 5��<�IT��`'*4[!dڧ�U�u@6vjk~ <ڗ��?e$p�^�W"1�%��0��#2�  �h�S��Q�b-�J�$�Ъ����Ӆ�;������s��4�Gq�1m/2�Z!����!;���~���+�HC���1�[-fv;��I=ߔi}�I�8�.j:~G�����B��0�: bHĖ�\�������uK�8��g�ϑH`�\��=�gf�lh`�?XX��lW�8��SDS�@�6ە�"a
�Q�8�!E6��5�¥�WN���)��ȫH�K�#�N�:ȇ�3�5h9�{������P��`��7�κ}��w���N:��)Y�h�R�����;�����M�I�M��P:�ѭ�R�&˶>T��g�����ck�=���n�Wa�gD1��<����,�9������}�
�R�7��]<�yVJ���2���Y���
���T��+�T�yY��h���̊�4_��G�n�p�@2�q�/��<�N5	n��y���[�70�U3���«��m�n�N �o�!"oR����~:�7�_�����T�&}����g���2�}�o���&}�QIx2֣H��	��6��I.6���u����~�	�1up%lGϵ�Z;m��/��L]�c��~7iU�j(DX�����q��}>�{s4����ʁ���ӧ�i!���t��<Y�c�C�KJM�8�ONU��op�3����ڃ�ǅ¡/�Vu;��}�w�Xl	\LF�XA��6�3b���x�m}�Zx�@TL��������(s�)�?x1-��J����q���	���(u"^(5����L��̤	�kc�;q/L�6NK6�T�|X�e�K��N����#�K4ãTi�Zp�T�֙�!n�
��)3��ۮ�#�-���;=שM�x2����OÄ́�J���hA��u�#K����7!�I^�l����P�%S�u�gA��Ny�G�&�Z��+O�o.'�.�C���*1`�6�@4*��&�D�,�>1�TH	����9�8 J�+i2�lu54���7�V�@�AG�#�/��Oڇ��)0�ӊ��>u�&$�1�l&����`��ys� �f���vxY�v
~�^XԽ{Lhz��G�G���*��#�ޘ�Ϡ�X��k\	��t��	�S�RP��y���!1�
߭����r�'.ݳ��s�Ix�ժno���S_���>k��v�6T��1�-��h���Y���W�&dȅ351�G��u���"���B~�3�]#Z�f��A;���Ӄ���э��[�+������@m�Y �������{F^�����P��$�Z�V�����g$����i��w?+GuҦ��l ���6���+li���I�/�1GH�q�@dr��,��k-s�5��OO��>:�0j�_�6�p�ǲ�H'=5}p��duW���u�㛁�<�.��E���0���3k3�ႆB���UI���o�z�.���P�A���H����sm�҂�y�\{k��^����1����7,��%d2�¢�&�S��D�=��>���;�C�8pͻ	N��v�Q�A6J���<�R��:����KUA�x�{Nߏfi��� 
\��% �>�覜��qgv�o�%W�j�2>��<�k���5��s�U���f1B��i�r�/��~$�fwzP�퐌�w�c�PM�	��.|�*S�ȴ����\f֑t�o���q�r�x�����>*�@Ha�ؒy�5�Z���(kW��CK�v�j���>�4@6�P�T�|�υ�S�G��'�s��f�A��>����1r��'���^i�
��w�U$����J���2���@�>� �&^��s�`�����5/��6�QsՒ7�eR�~{���%3�ʓ�D��3��Y��S����D;5a�k� ō���_[(��Axb�D�ox��m�m�T���t��݄,����N=P ���ZRt���(<�gPόW��0��`���nN�	���@�F@L��	�[r�`q�	��AŐ[�*7���g��M���p��\��v5�YZ����5��ୈ�3E��I���˴����q��!��m1_�"N���o�]�Sn�����	���b6���A�������ж�r3H�4������"â�+:5��f[��|�m����?t�{ �8��#�X�eF�΍G	�Ͻ8�S1�i֥�'jy�	Ě��������6>Ѓ�������H���0ߛ�����b�9��<����͆�f$��ec�*꫇Q�̫/?F�:�V,%z�qxJ�**Á}�7)��P�~���hs��12]��K��y\-�C��}-4��u�:��T����Hx�)�;�]�ۈ]�esF�v�7pt��b�@�GX@%�7sa�%x�9\�X���.[=g�Ia�3��i�bk�>�RV������(�����0x
�΃Ⴗ�툗D(��~����s���'Q�!��>XB8r�f�\���<�����){�� "	_�,��������/t���w�����wDt	���h�: 똒����]�
B��Nv��9�$�/�Y�0t=f��dBI�(��r\lm)�����Ԝ�ەp(
(�N� N��(!�u�g�M�[M�[�t`�T+3�z�ø�T�@�Ѹ����o��.�itB�)k�E{�vɍ4G ���n�4�)��ؖ���޴m��EU� �c�:S�T7�R�\_�Q���2��s���ZR��j6w5q��K�{�S1�x�����}D6���zM����Ɵ�	�}A\���.ϼ��`��i_��� �*�KQ���|�&C6�J>�@�}��9�c�+��^s���p��T|�ϪӃ���ޡ�sj��w}{��;##���� L�.����Z���U��v$Y��.5�LVx�!t���t�9o���S��vb�@�����f�H۽dr+d(��o"ٽ�$N����j���7�q�W��"{uH[�-Ǎ;���g�ft`��)�q�%����XH�q��R�� Z��B.�_�%��Tr�9s-3o¬�����}�fe�To�IM���u����Rw� �G��b�RR�n.\�RW�s���]�9a� �btS_�q@D�y�%|�"Bɉ�����!L�l
�@V����S��7(t?tjz��sڶ��Ѯ%�}q���K�|�@�\bl�~�KJغ�;��x�UD�G��?�YQa�/wSx�5�r^QD��U2�����1
���S(>M(mR6UQSm<�$|M��Lyc_�{�ypivv�x�:�6R�t�oxU]�Έ�l�V� ^k<*X���N)��@i�2l:F�&n5u���\΄-ڲ���7YK��@��9]�i�cX�j#�,���H��|�?�`F/٬T��x{��-��Hz�:��z��W�AX�8r��z��J۝��N��l_3k!���Eh��6�?Fv�]���s��K��36�#�7�����4c%@o����WԩȢ��
�BBKU**2^|pS�9����R@�/ �o��?\�'��UH!V�'`�iӥ֤HDk��v3/��B_(���"�v�Yߘ�Jq��_��Qi>�,�)�� Q����p�h�_#N 7&_4EOg*�|�_V��.>]6���n���ǖϱ�e640zJ�j{�Ec�1���o1*._��V�l���K��]M�;���g���KVʇjb�|����,��d����U���PϽ�2���J!��F����H���S�7Y3���ᵔ�gZ
$��?6Pj��QuWh�ct��ΙYt8�  _N��7X,�u-Li�c� ��I����/0�[���JW@ʊ��K�!kV��E6�7>c_�]�4i�|S2]�\d��'���pR�W�iBq5�j��PYZ��W7o���?�����I�TKt�	A���u)��x��ؖ�+��$�7!��������T��8c��+ⴆ�&"q���mXD�_w�Ȳᘬ7[-K������u�A�Phs��ڸH�Q_��ĳ����}���Z&ꀾZ���bƕ�<4d�cHE���3��\O�J�!�,B��p}�k��G���6���m!5�������b�1�b��wm�>�c���3��H� �ųc�,�b��s�M0��?�����U����L��D��R��rB�H�e��ᳫq���!4J�?�@"9z�\��-�����ĸ��A�T�r�|�vr2d'��Gb	��d]��}�#9J�5�M2I0�\��\���xE�xC�������7�f��;W�)�$�N��\/8�k�*�X�J��ր�Ք��y_�=�6*R{d�����Xq�o��,\I"u�eTO���D�g b�o����H���X�g��5�'?ʽ!O����(�"���\��Q�dy�;wV������F���#�)�F�hf�J�0 ��mw^��G��3�=
�̺&��	��v;���$X�,��[9���1�6ۈ�8d�~���x���� bF��e�&ȯ�Z�)�[p���_��|��A�������UB~{R�~!�Ռ!�o��Y��?*�#�Q	%���9_Yp7x���/mc���­��<;/��Rr�=��H�
(�DB�v�fL�P�/E(�ு؆�/���-)�8�7��y�OX���Q"�9�L@�(���	]������&�-G���2+e\Q�Iz�а��K�>���:7@ �5>�6��H�Q���>\V+�[�g8R÷@�o�ɂE���Äh@����|��7�lssO,Z�R�	��t�lV��t�:���] �鴓��gH�,�j�ϭ�	�,r@Sxg�Y ��U �f��q�PW�)�᫗0�4�y%�HtCLR~�2z&���o� H<�)/�ᜀ� /����Ȟ�@��=e�t`�z-��E�oD��'C"$�F��]�m��5oM�Wgt���}�L�������NuN:�v�S���f>T���3��������J���c�Ef�N�*FB��d��,J��3�������Ud������I�(�7�u%�O��RLZ�6��yz�M^h�P�F��J/	Pm����y��8�z0��J+0_"������!��y
�w�P�L�~��J�Ƃ��z�ͦ,���mN����ʊ�T�\�h���ׇ!mHc�l��9�I������GP��6u�+ƶW݀����'��U|$�l|�}�D�e���o��O�B�{�Ztj�c��`%����TH��-�2��5�k�9�@��@��!N\��y���cc7���W��A�c䄃���V��s��;ٜ�%;�|��o�5��J��ڞ��&kR��ʚ��yw�hx��(�3k竛�����sbN���s01�<ʟG��I"/jM�,E�㲢��H�� � f����k$Mr'��A�u�4ؗ��z��*���zM�nn����b�����z5B�w��m�F�Puc4��f���l�3���i��	��0�1��Xj��$n�l%��W�X��3{]v?a�nV~i]��|\���y���Su]�Nk#�Vc��* ���8�Cw�؆!/i�߳8e��@�����^zY�u�6�׺>�9��  ��M{QQÀ�Z%7h��kK)��Bzh�́���&��N%Ul(�V���U p�1/��L�P����Cu,���Պ�f�K�1��`��[�0<;;����rT�T"d�uB#�� l#�7n���?�;���[����Y�H-��D�%���@�9c [���������r4�x]}�P�� :�k�t���\�E�aF4���,�UB+aG8��ҍ.��'�J6��1��*������
�Cd��� �A�)Ã_��l.���ׁ"l�sIȉ�&wÛ̦��4]�n��;�t�y�>%Bm�^%�e����$��}��^���lj�.�����H�Ncl�9ѽI�℟H��m�IЯ��_/N�=����9�G�*%��#�E���9QH�^kS�ǃ��H�n��fO�}�����E?�j��s�nR��u�.\�*�,N��JP?�9 Fi]�~H�e[���X
�݂��D+�K${}����&YH$Ә~6Ϟ��^����s�q!�`�&+�v��5�G�p*�%*d��ómm��+�W�M�ҕ��9��6d+'�TK�zW���G�=@��,�Z��ﶾ���<�1��O4a/'4 hs:�VgA�F��@�ث��)m�����ٻ'Ő���J�hs"Ȋ�SZHG��5� ן(<�G25,�Ò��$���ІI?���}8,�Q�*�BcȞ�m���\�<{5<��ʡ�ꉶ�[��!X4
�y������O�%0���)錏A�#���"���A��H�lH��;a230�K^�3��y}�ԇ�)���ʇ�ze�� (2�hAo��L0�̓[8�˚���kgh� �~�G�!jڦ�� ��=i?�����"$������C�d?�Ap�¸R��M�.٥'G�k��M���9Ee�l�w���	��k%/u������@:� ��E]��|�j�5��d	����Ƀ#�S\�ɭX�,eǮ�N��m��w|M����W����um��:
fI���s���oP7���VV��ߞ��Y[�nlq˓�x�N����8G����]��r���0-I����<�n�Z�OTf���H�mnxm̏2����d����x��,��1�����	�9�r*Z�K�D�7`��֍&�JY��f�j2R4Qs�E���a���/�qe�н�M�����ٓ��bϣ��ޥ�\��]��1N����6͙�yƊ��ZĬ���Ԙ�L�R�G����}�B����6�1E���ĀDj���8��yrjmǎo4����j^�,��1t/���/��� �&��-r����Q����`3K�p�#�[�l!�Hh�1�&��i_v����[W*���z,�ߴw�3cM�;f6�uj�t@�4�5ۙ ~[��Z�2	�}����_G>�DZ���/���ղ�Ը���c�|Gb��Z��&��)Pc�XO+8ge�Vk.D0y���_��)�C�N�^����B涯l�
" �b�t��2�f1��=�=�#i�i{�:4X(�=����A�@���0���ͽ�����P��j��-�O�m�L&5�m%8ee>gqk��tp�^�V�(�� ��1�K��Z�5; �]����ze �[��3y����B�<����Ĥ�"�E�e�k�= �}�@����V]\��o�Ԅ�9�l0j��	LZV
�Z�2&|�)H>Q�\�hK�GfH��=��3�CR�����a�g^����@����^q�$W��#�񨭟X4���]"�kSb�.��ngG�#���rB����\C�=�}�(^�%(	ۭzh�1)IН+	��`y�,?|��~���8a�v��a9�+Z�:���P��9�Rr�6���U��N].�&�Að[������i�d�OOs���X�U��:/i���o�X��H�[bF@�x����B��BD���D�4~:R�s�ʩ��	���L<�ۍ�[��^����oҟ*N��f���'��7�B<��ˊ_|w�M͵}&^�r�|��Vqvc~�����m9�5蝁G����Bx��ט�]�Oe�%��	ѫ��D6�}Ŋ(��z&��4���[���V���q%���u�Lx�<���΄oFj0=AZ��m��#y�y ����	C��/���Pm��ii�\#Z?�����0aoH�e�ˑ��ܦ�����!#yz����Q"����H��<`��T�b�o_�q���q?$��cݓ��齁�<�}���Ǚb�i�N��U	s�D��t��`�;+� N�{o��<0�pթ����}�̴��YJ����h����N��-�Y��Y2,t���'?t��KH�ϲ7�w��K4r�·��=�ZwO�6�^r��3�������/2&�n���d���$l����'S���g1j�5���d:j�e��]�3�y���gc0�$��'A?��	��P�a�fy�q��'V�e�,ir
�\Z�-�53�s�V͊�>��������hў���^"�+�T&m��`qK:m^��҃�`����1��W�X���%�B�sC�I�A�9���b���\p�l�|�p��#��,L%CH��a~���
�����#�u�(��aS\��y��{ R��сX�ukQ}�h
��G(R�y͆}ho���ɻ���Qg�(p_��K�_���=h��r����H&j�YCq� �M�h�ӣ�N��Ǹ�6���B+R����/��A��� ݏ�k���Mp,V�-$=�(��D�_,k��H��� A�S�s�8����~귢��u��e�R�l_�8���Nк� ~E�_��ݠ�P\g��S�p���:Y\vxF0�L�[j��?ȅ�k��Ps���6��;��
ۯ��'7�M�g�l�������1�BI�V0���W.��%y�wt9�x�{����@��N�e*}�������
���F�R?zy�`�A�w����l�xm�^&��E<��&�h�y,����8��u����35ⰿ՘/�����ZhA����ʧ���(+�%��QȲ��Rhq��jI�d�a�F�c\�I�i�T/�c��ѝ�sޯ���ܽ��Gω)�Y�P�)��56m�/��2N9<V�[�}h`)!��� mv����z
�cݛ*�%V?/d��/_(�ى�g7gJ�|�2�d$��m�v:�3<���1�&��W0���DlU�wki*I�;��~��Utu-��rd��a\g�V��M���ܛ�,�U�����]�#i�2��3f�A�kK
�K\����<��*_ +�؎�3����c��5i�<9���;X"�x���f���<s6mR�wKZ#Ԫ�<����2�����}�U������h�\6!�A[f��ܒ3�V�^uQ��2�{}�C#�����(��vt����|E,� L�V֘b5U,1]�i�c�ǜ{kW#4a(�����7�A
���m�3��e�(<�<|�O����s���-�N*la��I�|��>��Z� -vJ����,��I#ΰGu-5���ߴׁսg��4V���λE<UG;���[8�\C�A�\�Z�^��+6���B�@��I�{%� ���ު*�1�
F���l�ҥ��@����z�����~��*&�oG�F��n/U e(�	t��8f�T�����:��t����.���v�;JI�e�]�����;D8��FB���K;T\�k�/x�"l�9Vn�[T���p�) .��T���[������2�3z��x����Hî?h���l�ދ���|�[����y�ϕ�$)�����;����А�*��$�[�{]^����
�<p�� ��\��� �)�sUK&g���x��%��C۔�:�I:� �eFcw:�^�>����kO�/��z40P��$�E�J�z��4*�o8����5k�N��*��"�'N/\�/����e}�� ��m���\���r̦�6S�fX�h��,�[߃TW	H)l�EW���V�qp.DI 2�i�s���m�{j��p�hL�8�cj���*Ƹ���W��7l�0�.#O_�ś���t�D���2�H>�ZHY�~�q����h�% ��&��.`��˪r�y��1�1�o�Շ����k��hH�@��S���֋�O�N�ۂ����9�Bzu{�]+?5u�{3��Zb]S�o�[�S$��Y�ҒX����W(jA����MH,w��Tl��H�оI�<�_b�V��\�W��,�⻊��6�
葧�o��hΒ�}R� 	d���nh�UU��>���k�� gWiq0����e��
�����Oӳ�"�a6��coF]#`�ظ�ɧ��4�P!,V>��;o,՟D�~�g��1jc�~�Ici[)0��ݯ٣d]�@�����Iqq ����{[�C��z�.�W��d��X��mD���1$r��	g���oG07��0d:�N:T�L`[m���[�	٤�FA����u����Ś����omf5���
Hp*�����!Hk�����h�W�2��ޘ��3�����cV{z���:ݑ+m%�r�y��]�Hw�I�wX�C���3¾��K՞��{hi�/Br%��ӊZ�M j� � N�Av�h�P�����N�f���ef�9����w�-��Q��͛��@���
�m]ѶA�q��f۱�_����������X׷�@�S��N/�L�yV�'�yj����0�4?w�gř������O����[+������9o�e�E-������
C8��V�,��@u&�Nɯf�����q��@P"޼T����k��lmfՅ�딱�!�i#��Ź�G���H�NAno���+�C�
Iӛ2��(X��b�C��͆�v�����M�^Ƨ)وV��Dy��6ׇ�Nz~L�)	#;}SE�mE�w$�׳�r�6��
�B�O��`����hni+o��s�v2w�Ԥ�\���&R��A��S=OO��u��zE�*R��b��V�e Ι/Й�gc�0���U	V#�8�;�]B���#�@�9[R�$�V��P�_~��k���;�=?�͚%�}Ik} ������C�9�(��$��PD $��O��JDZȧ�\�J�e���1��D��A�o󅋈�5ă�3�6�J@[qt��/�p�s ,�ή���zn��U�f���S�
�PZ}��O]N離�������<Q��k�q>m��Ju������v��a�.w��a�ϟ�<H����)#�i�fr�h\��4��?�q�j��cz�:���vɈ���(����C�i��%��{N���h��$̒�*R5�T(@�߹��/I��z���L���˵v�s�n�k��Z�#.��)�9�0Y�f��Z��e ��bC�V��ƥ�0r��	�#�8�G�;z���L�ְ@R�XZ�����>ƶ��^��"�������s0"��#���5���;D=]��@��3Mc�}�'�� &U�}˅�h��lM��d��b���5b�*!��.њ�T�X+�r���v)B��6�Y�6�!׋��I>@6�%�����<�$��f]�"2��4Eo�T���8��l�ID�pnS���M���8p.��I�k5����9�V��v���Ex���ˡ[�Z<���W��g'��-Q��9������2�xaۭ�粖�)ސ*Ȕ���x� �� &!������*x`�˚0T㠛$҈�A�~��c��L;l0���z�o]����"eQ���F���MBZL��i-����aꯕ]A3�S�8�{�m��Ѐ�D�$r[�5�f�^�	��U�
��^b���
��F����Pc���<��-n43e����?�a�򼉺[��Ek���2|�ѯV������Ħ%��̙3��%�+�R��`����7й�=�'_��=]�������;��v��h�H�Z+cȅW��bL��5]}�'$��RXx�ܩ{e����eWڟ!DjW�~)B�R�ӆr��]�9'@������:5"��g�V�|���c70$�s�fq�p�'��rz�E~���������[+W�
l���W)�[�I5.Ah�6���`��`�n=<�A���r�M�Ƒ���f:Z�����L�K.��	��̱Ghp���U.Z��N�_{�Jg�{-�O������V�Ps��m� B�4���i'����LMa���,G��d8"�`�OX�7��c5㾀"s��]Pi�an*�,�v}W�P����(;
�����7^�x�+�z� �{>��"3D�H��z!�������׃�l��q�T�����-�q=_�J�j��+ￆ��J^�^��i �9�@�ш�نd�u�#@�|!1w�>�w4� �̑F��� ꇍ��*�����g�w;�+2*���aP[�2v�1�	��zɛ�wz��?�\õ�}"��4�5R�
�E9$FMl�-����g��Dܿ�3�Bv���;�x�z;r��0B�1�z��Sv�U�y:u�Jr��gu��CsԽ]%�e�BϽ�(�U�&�)��'�ьُ��8 �b�q��OiZJ�ǁ]~�cظ�w- Kq��a#:���J��q;�u �H����x�@��)lŒHvtM ��x���]&Ȕ��h ��^P�����?{�̋��*�]�$݂\(�y�!�.~r��ߊ�AE=O��G��<l���ۧ�ו(՟��~��������ޘ�YP�� ���#�(��N*ҕ�l��[?�����;Bi��$�ף�q�32�\��&T���%����:�>.��LO6/�H�ݍ���S�l�d �2�̀��6|�G,��A�$ˆ7�X��ɒҽ�x�o�e�[t( �)u]��B��vM�'f[T4Y�&�^�Y�$�o��S(Ҥ$���~&�nvj7�d�\ܲ�轒f���P�;邕%V�[�!k�;���_�@�[�%Њ�z/̂A��������v~#��$W38��c62��f�S�|��畡y�)5ݽ�������*&}(9�M\�=~r_E�.���ɘ���r�It ���8�R���4�Tl��J�	~b�+�-�H�m���5�g0���0 vCRW����p��i��ƾ��B�����]�s��R�*��8��Z� ��ikD���+�:�E�.�}l�x���<��,@��� ���' �o,�+�w�Lw��0[�<���|%ϭ4�������t#wqf�]l�\���r%w���g\�ӈI��	���/�4��o�[|�|� �}��C����+TI�	��֦�ݴNcʡ�#[��q�NA�B�BO��J,��2�&��X@��I��� 	��B����ֱ���[R����]_K�#``ۂ�K1�7��x*����s=l�3l9`��2� �p�@��2���/W���F(~FjU�l�e�eO��5#�>W��k(�0Ի��#d��W2���Z{[����$�����^�*��b�S��Bwe�J�����֕�F,2�@Ha��Xbj�cA��"�"�r$.��-�Ss���S�M�T��ߖn�e�l���_Xu�YF�uU��z�ACWC �O�@�s���v����K�b�=
H��� l'�I�%{2]�����/�7��+���܍i�1p�bVI��ӌ��W9��7[�:z�93u!̀�}�'#@U�g��t �����[sJ�Yx�V���� ����|�D��)(E�3S.IT���Kzc(�,PZ����Q-���Ez��w�R_�W�`Ţ�{��8CCq��U��+*���EQ4/2������3I7V��=Q�)!���3?�d��*��rE�VvD�z������Gkح"22"C�3!Үǫ�K�cgם{�����֧Ͳ@ƀ|�~���<� ��՚m��[��o?Je]fQ���Æ����!	n 3�iKv�o ]z�"D@�/<`�4t"�񝥲	�Z0��pq��ʹ�����X$� �<Қ�3���e�1�T.R�50y�V���C�SD��1�f+j��b�.�e|���c��x��X�v��1^`�m�S�����/��~�9b�p�OU"3�Om��N#�(T&�`&];��K#���%\���6)��+?�ѻ1P?,q�w^���fl�������@�v��z�X�:(��$��d����;X�� ����/���� �k�yݞ�2ϐ���WB��s�o�N�;��������}����r�rQ��_��-���De��k��l_�(%�a�]k] �7����{4�����Ĵ�a�Q����4�<GJ�\}'Y4��'���I��2� ����3N�Ϝ�:h[����G/p��������6�>���i:��܁�������p��_D
��-\۝m^$!�:C�^�3�T^¯���PnAC$�7LO)��O�L��2��"�h��,�Q�9<�1�~� �^W{��L!E^~�Y�TIV[	0}w�-j��΄0l?�e�g�]�u��;��IA;q
���=�������h�@��u�7����.j^+�nlϯ���Q��!�o�.�-��I.��Jr�ET��E�d�A���ݖ�T��ˑ�����r�0��N�f�"�M:S'�e<�Il�dB��(�r���o�Zv"w|R�|��E�uf��?-�i������!Q��;Z�/��ޔ��U��✔|>ɝA�d�R( 9v�;Ú��.���k�qb.w�N�VN���aa��k��CW���e�?���1��hM]ߕ@��.p�V��/Ak�.��z֭�S�lP�1����vp5y="�3R�U�m��}PVԖ�\(3���W�T�W�����ຳAy��+�����う�{fO�T#okcj�;D��7w�iǎѭ�u*�X�4:�z�V���+{-_�^���kM�C^DPw����GZ�t�h�,�}� �u�Ct�-/!�~�"�Y*�J.�؛L��S��9�����"}��gx�_����x�q@�H�D�NH�b�H+�	!���7��p=t��B3֭�����Ӳb�d�'����3��u3��U$La��*U@��P����#����Q��
�g���ٲ�Pt��7"�����z���:	�cL��[��@�_TS�[�`u����m�29۬OI��A@�bB�^v�HPy�;��Χ��Wz�rNm~O����w��WmøFm�\l�W�4�6b�d��Jll���:rۂ�*�']��}g��Ly�V�B;�I��R_�<B���އ{{��"�֊��Q�S��p�f�h��tІ�l����	5@)��Ry��ds��j�g}�� �[�W<pߤ����`�Ef�e�l��T�x&�B��9�=�������Ӭj��!��Rl\ʶ����
��v�O�-6랉gc�'y���g
EPW������c]DT��b��Tn��;��>u�)z�X|�@�=�6��i=�d�U���w�^J{������Ө#QϷ����s�9՘ፅS �ӳv-�N�teP�&7�������y�S��Zq�Dwa�������|Y<�����j��Ԭ>��kg����'�*��V#LH�f��ztn�A揌�������u����~��}�^/o�GFz���t:���b��2C�$a�Z��3�~�'��L\�,��_ V=�[�6�F6g��ۊ�>��M���
8�&ԅ�v�P�>��{J�MS�i
�z?e�>n�$҂�x�Ж�&�
w� �$��ߐ���Y�1a$Sg��+�� �M�o5Sf���~��üD�2�5�P�ϑP���-�Vr@Q���V�w���\��<����̪�h7�%)�[�D9�X�jŽK`�A@,��gd<`��!+�}��)!��P�/��`>�hww�1	�o8N��~c.I�����իA�I̍����jE��G`��&���+�<�sW�F�\Ľ�5`�� ��?i�kҏ�$6�*oI�%�)���l�NC���}n�<k~#�{����˪%�S��:��ǵ$HnC��c:<T#�t�X ��,%-�s�����bo�Jo�XM\JW���AIJ��H��2���z��}͸I�����������\Pp-�d�7�:�9�9�ʠDN�=��������P@�4z h��c՝P���.i�R��1���,�`�5Et��a����U�&�mm�tL��{X�0�zq�NO��w���u���z�hL�r1����u=�R|���[�u�mY3�a�JSF9�D�	���C@��45�'�MT����\�	��N���Fp�}����C^�~��VȖ�l�򠄷t��Q;����x�E�����D���_�xI�]��Oei/��׆�F4����7 +R��X�4������9(g�R���n7�M��u���� ��;�Ղ����.��}�)<�!c73c� �w:|�7���|���H�?������x!S:�a���F�֪�| ��p�h�[��7v�,�j �m�eP=��]�l{h�+�=��9�!�d��BçJ"�k^|u��?o��{�=o:�P��9�Kh1m��i�!���%9$�5�iU�ev��P/9��� 7�le��W���q���X����VIdt&QJj3�t�X� �>��P1�9�?�3��ٗm��#�N(�������z��	�F�U5:YJL���@4�����27N���B/��X�Zu����,3�?������2���%��.���	��d%�_V!�:v	
�k�#�&�I�RԷgj�G���N��j�?�w-!�����{C _���@�`��[�S&[%1UVYԢb��сE@AH��#,L#?��}<�Z�Q�m��ϸ��;����8����V�0�J��} ��Z��|-qPW�R�a�L�ێ�G�	����K�ٻ��ك.A�-�N��i^c�� KX �,��A.��T����px�ʵ@A�W�yw��7_>���sCÏ����&#�s�F0�Mݔx>:�#��(F�si�(�* �gw�)ǀ�츍)r3_����J¬��d��@<[~�j�i"�w�;R��n=��-;��2P����.Xťv��"�N�d깂A�F[I�7�C@I���;�����t��y������UO��oR�������|��V���^�%e��~S����`��Xl��>����pLO�4�m(d��>X}\`p=�g�;����j:b:��4�ʪݝ^g�xe�H�c7�B]���E�Ϯ\�Ty��=EQ��'�~��r�Z��*'"R�jj�[���Oׂ���3�Ξ���hX�xu���>d9�g[�d����>e��}�,��\�:Z ;�Hց�å�m�=�!�*���Xp����7^u�1���ᵰA+|�y-��F�m�������⳴�P�A��u��@�_�9�P�̷���A���f�E[��n	b��Ēd7J�a����Ǖ:_v�a��5\�gac�E&�4�Y
�4Ӊ��;�,���;k����j=#��G� [�uGj��(#���]�*�U"��啧�OE�f�Ơ�)Q��A�V�=� �I��]A�O���y���IO�ښ�:RYP�s̫���	��f���ٹ�?`B��?�׸�G�FL�r�W��<Fpإ���`�ѓ�֣�	���Af�*'�����YaL��������T�z�hoC���8A���;)��H�<�.6]�t���*��ɛ��}SrEa�~7{"��1�.cL���tw���@u	���P�w��F���z�!B��y]��T!�� ���8�bv3~~��Z�����У�&h�{=�=�H� "ޞw6��dj���$%�۴��qH��w���%ι���Đ����	�{�ʀo�#�����#%Ǫ��槬��!hg�;��C-݇e�N�������p����Ew�M�"��$}uj��ԁ��?k�>l"�@R�j.t#A�@�fS\��c%�h�o# ab���/�H��>T]�w	�d/M�S�a�	'��bS`���h�F� ��v0IX�#JG�������B@)�3�@BQ��B�,
���<��ɣ�� 2|T�T�v�,��"�7ND��-�p�'s��26���D�.OʖJ>�b��D^�um��h��m>{I1$r���8{��<��#'*�[��.�K��]��&��MO�g�mb>߻^Ɍ���g���1简_Ǌ��i�b�<	t���j���~p�L���UdG^I��D��p��m�Ts�W��[p�پ��ą�@�v o�6w�����8�S�e㸌j(A�T��b��n���,Cd^���UJ  U����bP�bڳ�O�f �t�'x��fn�K�"�G��;�R�D� �.���-��I�s�5�W�������Y�0���&���3�֘��� ��~;,�=BG�\���. �^/~�j̜hצ�)��:��-p%�Yx��>&<E��k	�r��1��f����8�QѰXl�fp�2�S��d�p�d�<���4���ѳO<�ׂ(�Z>�U�|�#�]���WH�!]i��� ��7�t��Lb���ճ:�Ҹ�s]��	�J@� �,%>���7��9H�k|�*L���&t$Yqڥ4Ë��t�ꩼ	���Y���q��o�5Pϓ��'�|E�8| ��8/���R�]�X���� b�{6�7s�|+��J���VoO�s�بm4G�7&�������#5��6�y!d�ϭ$hZ�(^���G�ș>�:W��yQ�����\[��$
�S~~���'b1��%wK��;�����(��I�*̔P�����b9t��bk����J��_�h�{�eO��[�@$ƿ:�L�yDn�f��0�XF��"��x����(���2:I�8��g�����^RAG�Ӹx� �ߒ>�-\�M�rr;�{�i���\���`���`r��V-�ˋ.1#x�筺�5��@���ڄ��Qc�8�&��v�8��SӶ�Xe>sa���ªp�����3b���1�et�B��0�ϱdi.�έt�
��S�F[��b������N��A(��ʹ��)ƠiWTp8��ȭ����%��i7N{��%c���_��,�|ԣ-��x�6/��F��م�00�1BgiΠ�d%Z�_��u|"#�A���i��"QÂ,t7�����ao2��ʞBWc���RJ�~e���B�Za�&�]�o߂���w�|	ޏY����};+�5 >�R��d����`��Y\Hi? 2=Ym��)���B������)��⧄��c�g�T�D�4�����j�L!q��?�?�2����UGv�]��X(�I�oU��U��h(Z�J�o0�P&�2*��3�f̯$��xk#<�ݯ�ӆ=$X-�`�|3�m���w}�|��]r�%�����!8Ԓ�HU��@">OClҝ��F�ۯ�NcQnR2B�s��&f+�[�BX�+�"���c�(�,Q�B��\�{�(�H>qewuN�/v"s��[4C�MD�@��-^������|��ˬ�7L+Y�A~εu�aZ�<ٍ,��q�{QU���������R�����2TwC��cbD�.`�&�p��،XM���}@U�v�6<���2ˍ�6ѷG��>��`[��y�<@�H�������9^�d8�m����lu�>�.�N��$Ҁ���֥ �Mh��6w���u���^�����?�{��@��N��� �T8S���RY�'��o�L';�\�'&��zR(���y?��kh
�M���j+]��<�<��{.�@���1���iy�m7L踏��?k�߭E8��,�U��1z�7zܜ�occ��y�`��K�i��0��]R���S2���~�^;p���?=9`\j��ҍ�%a&'rō5�/E�^9��@���+����i0>+A;��2�ۆ/՝�ғ �}��W4�L��4CbF�1o����$Q���٪Qy3�Ԅ�&�OW���j��������I3�VQO��<E��J2��������cRRX�B]1�/͖q���b��FYA�T?B�������E��=Ke�$��>	+#}�:�[3J�B��z�⟉�-���D�P�ӟ3�Cu��x�VL��|�F>���4���ʏ��Z��7����#��m���9��gDX��{'�}\+�ƌr������^r��\�Un��.�R��)��xI$��+�,"�:v\��mŌ���1��P��_Î�y�/�N���T��n��B%>�\~$���B_!� U��6���K�����7���Լ�X�|&,�]�,��\
����X�(%��*���G�pB����"��R�{e�ه�-����`�h���͙�p��T��v!��9�
&� ���7��soDF0����<A��٤�Gf|O|��O�yH3R��_�e�I�`�?��๸��`��O��L�B]�X��Jr!^�� (��n�Gӫ����4��5-��+v�G�t��mk@i{�L����b#M�[�m&H9�r� ��yۯ�v���1f��h�I��O�p3FK�˟%�C�z.Y�]4��K(dA��y���9��V��2��v|��9�_�\��^�җ�bi1^�<f�/� %Z�s�f9�!�ļ�;�G{8��w�����T�J�^��u�U�N�m��@�K�kIL���8�G̫�s�i�����f�O�@���%�a��/A���_��W'Dj5+B�(��3�KZ�'�!.?�dRH]���*�c�Q�����s�о(g5q���9.�j��)��kS����֞��M�o��"P�U��r�/�oN�v�{��s���X;S�ҢT�E|��<��@� �a8��_��s�K�6�}:a$,����F�9�M�x������������UP�{K��L�C��R#|d������ԤQ	:WE{I�m{5�4�������)�[eM�
�.!�&\Y,�%��;�e�\��p9�$�#��FKD5����nh\�|*X�pX��P<��O248dc����iZ��jo�w��;���)*��ӟL�I8j|cx�")����VTЫI3a��jB���t���l��罬�vl���6�4Z�k9y=/t�#�DG�E��b+u��}���}*p������~R�8y� �K��8=�;$Nx��K(�������S�<w��?�}����P)��
��( ���`�([��I�A��������?��l?zA2s3Ls���t�y�['g�T�82���䔢^�.��D��`�SڊSs�����L,40NǯP��M�l�%B42�^b�O ��A3�䥵�r�s�e,��L�R:4.�w���sx�$9-���\G�`,�i���ّ�����K�f�����̄
MT<п����(:�O)_�~��ֈ�8z�%�a�U��Ԍ�>z����|j�]�6����j��\�!d%	a������y:>����nʤ�~;ܱc]��[���ٰ�����o��tb¿�P����w���Y)r��k���q��p-Hy�����E��^��x���R,&����$����2U7|5~��~,E�	A��)_f��UZ�����FE�������Lr6(����X����B&~�`�]i�G:-�l��2��7�}���zWy���Ŭ�c��F��Q�|���Upo��5�	���JA� ������k���2�����w�l���c���L]6���"��a@k̷Z�~��=d[W�ɳZj>Abˢo'��@�(������� ��Ƽ�I���vά���ഏoc�|��NM���C�����#/��Y��o�f��O7�#-9�Ѩ5�A��V�Z�ڪe�#+X�R�^"�\����U�}�6�Q��/6͍/3)e��#n���;u��I�iv�F��;��*}�}�}�>ʟ���e:oxw�>c�e��?]PA�PA���y��(��N�^�v�Yɰƴ/���Ό��Z���~�Эu,�%�S��ؼ��� ��y����$��&ZQd��w����ޖ���/��G��9��]"a�yw0�Q¬�˘���f���Wx�QC���t�Y�U�g@n�v�+l���l�0@P��ny"D7���+��D�<-�U�R�C���D��r�S�:;�)�%�t`
����"�^�[ʸ����ܜ�^=z�q\y(k�0�a����4���f�$��)��r�b�"c�e.՝vcB]]�������� *DU#��ӢM���x�w��Х��m|k>1�a��v $!�z�3fDM�A<�K�Kke���������)~�o��]����[�z�*Z`�v�V>���8����;#�"��nX�S�ٖ�H�=O�C�ϼ���#�{`/�_�9Q>��\���NW�R�"� ���������s��v�Y�DP8�t PF�_�8�+�eiuU����=[������^�� ��o�������4�`���j���Hݥ�������-tF��^���Eg8nf�WR��=�+�C"�[̞ҿ��%8g:�:eZ�"f` �x7q������E�����,��Qf�c�7�q�)�~L9	_a���vG�߄�"����,�O>X��6��fQ��b�8+��&�y��T��fRy'x�xZ�h��So�>��]EУ�!��	]�����Է������;D�Xz^��L�۵�����r-�P���n'}Q��dB���Y8',��ZN� ^�(}�-_���/����*&�z25-����c� rӗ2��T�<����@g���ԃ�F�$@2%��.�oꧫ>�W�#�`O�ިA8R{�K�NJو�HF�{��y?���Z?�q������c�>��缪�6���Nn�H��b�������!�����m���N�����Zm�uN�� ����k�:<_�0�M��^��� �s.i��\���z=�~��x���[�����(%�SPŤ!�yL�"�Lѡ8$����r��"�4P��*�|��ث���V�,��0B�'���s���>'����o�;O�`V�s�)��B��N�H�5z���
��2F\�ߥ�c�,���T�)\^C��CB�e���ω_
8ح+�-oY���
#��Z�&���o%^ܚݗ���>2%��&�U�7|@�����h]��JF��p��6�D���O���ې9��?0j[Ep L.�~��WЩIv�<-*��T>�	}�.?iV�]DJ�����iVӅ^�[�P]^��4X�qF��\ޕ�t[�:�����Λ`}�Pn���i6G���ǧ;���8�p`���b�,"4�F ˲����].(���K��2UG�����m�D/�|���b���E��&���=Ѧ��όx 0*m�[4X�c��ο�֋c
ج#D��i�	���;:˵&&E�������5�1�4��$>)W�[��0%�%k|��'_�4���j�#
eno�;3�]R�~���!5���Ƥ0���)�Q�v���v�^	���~�stm�������e*�jl�|y�^�>����8O߆�4����l�`?]��D;���5"L_	��#3S���|����/a3�2񍈞#�{,a�0���ɭ�E��N�6�4�	��T�*��$`1&�C�M�8��T�,�Z�i�q�)l�KT���_.Y��Rl���ai�=�ø�M�#E�[�si�lK��q�׶�c�c�K�1�/n�����g�	�ca�2�\�2tR�[���冢�=j�]Z�׍f�E>�e�b�slh_i���� �ƏO
�i�����>��2��x�<���w�O�n��K������m�G�e{o�:Ktԯ1�4ܱ�ަO���J�<�MU��[K`���.`IF?�.�1ta�G.Q��&4��T�C�]��������F���K��Z$�	-�?yWڳ���JN�n�
����/�I��kUݨ���c���1
���Y�p�ھ8e8mF6�]h`Ѿ�c=�����Jnr/��(�Gw��7�J�`�O[���Z��b!kza�ي㻞���?u�n�'��o���7B�)��>a�|,��(��+�r�ⰿ��Y�y*�>��L����u$2�N�a_�L�-�9 �^��ȯt�E;i9|5�њ�#p�1̮<���4.�t���E��	:��]_CY����0��Xn2ji��	����5srή�ӓ�(��\=8 �)�v�& ���PK)5��f�+{�f 59PM���3�M�u���(I�HG/֝���s��%w�G�+�X��n�2�g���fMV���)eZ4� ����R4��u�G��#��x��X�ݑz�8Nǒ��.;����%ڱ���1�	bJ���?�?��H'W�yXݪ'�(��O������$:2Ľ���/J�;ݞ����La��i�!����ֹ!��'�ͷ�M<TەE���q���F^�|�G�� M�)l��U�h��#�,�_�4c����p4��l�A�E�8[nťց.ٯ\RU�nY�Ǐ-\�Tٳ"�8_����dw��<G��Ӳ%G6�΄s�3��n3!�y������2 �4�+'����TYu�>?_�(����b�HY��<䧥��j����MJI��N_���?���:��<��.T 4�0@��ܭ�ÚBT��Ja[ͪ���5{o(!{�ݜ2�g �z�����#8^�o�!=@�S�-���+{fdV~Z�P��O��P��P�U �ڍ�vV���
2a؄�7���.6n���uƻO&���)^�)�o����o�n	��X�}w��{�2�7���q����2ʠN]�6С�c��������{L��"��Ȫ�T�5b��B���`T����:M}u$f����1O�J�?mU�ҵk�N�TCGp��jQ��@J,����/�C�]�NC��)����� U���3$�QW��ꮉ.���Ɉ�:�"� ��g�vG����O܍Dӽ �Dkj�K�P�	k̵~, �8!���}�knX�X��`R�F������9֪�X<,Gͦ���\��%�F�c��G*t�@m!�I{�((��	vr����8��܆�[p��<�9��{�C�b��x2K� ߭~���h����_�6Ol��(g)��M�*�����>����e�8����7>�5���n����}L��j,����_h1Zl~C[��W�s���+����اWvd���]��F�/x��k^�q~�����7�yX�QD�ϓ�vM�DY�_�c6�1���M�u��T�Y�W�}��P��D�>ΰ�ꔼw[�09��o�9��+"͇��M'����V��T%��@�-^��&'\�3�,��s J�2���h��gT�C	-�d�Z~W�.)i�7~Q�잨��\����߇�E���ld{J[�����ַj��)���c�Eˍ�.dP(I�"��(�W�a; v���&��4ҷ���3(��Au�RL�@��N����vJ��!�V캇9�/�㍰/ܞ��6�zRj{BE����l�@����$�S��|�6�%U�h�hTuF�d��AD%.���",u��le�v�G ���N1Z9���ɕ�C\�Ѫ�ql�mi��m�qn�~W�#V7u u&�/M� n����!����|�q��S�)�+�쿥`]X��A�K.À���/�OP;Y�SYb�u�\�SCu�th���7�nϡ�HA�|$��Ƞq�*�;'ιi'S��<��a��E��[F�#��i�$Xx^4���U��(��ه\+����o�1v'd�δ@ЭJJ����δ�.\���]+���n%�P5��*�C�1q$�n���ev!N�'����T1�g�8�%;��y3��<��F�;���4��7{�6?�_5�\���ǆ�}�P*C��Ifx8�<{kvՋ'=�z_�'�.�SQ/��|:���Q �Z��L�X��E�V� � 3��.͸�u5E�Kΰ�D�vF������lع�d�Fq#Ue�w���ӥ����3�x�X�4qF��h<��B��NF�{��E �r�S�C�Wj�{�5c�h��ҿ<3-��Z��)N���%<,pt�+W�[���:�l�)�����Ő�K���v	P�[�q��g7���#�K[���O0]Y+��``����o���4��kr��_�΄����:�b�D�X���E���!����ɚHf?���Nj	�!���Hg\
vN����W��O���G2<��$�����*韫�Xꑑ���:gg�n+n��}Q��9�`�eQ��W!{�+�n��-I��̐ɔF��c�5y2{�����d!���3F���@���)�*��G{ߤK�����q5q�l��>��b4�9�+#�BO�����ݲ$�u�w	����l��aM�X2zC�I��G��bĉOOq�K���u��]���7���ǟ��z�@b�2SW�Up@�j5���wt���d�t��G��ҕ��x�߆����*�~��m�~a2ù�����'ZHX�����q@(Pޏ�`<m��$�m��jI�zMurT������9��TU�R�K��^�+���#���R�k�t
�^C\OI�����_ӆڰC�L3��&d�ˏ���5��)��f�F��_*�YV;T 03�Ō[,�:��۫/ֲ�#�/�_�Ԛ�#��dw������D�o]�WC�� Ҿ���U�@�&(P�H�@����X퍱~�቗���d^.��QG�2��
cj�N`˪��SXA*{L*����<�7�����s���r�q��Q�����\H�#e�9�[g�9���E���	2��4ڮ�y��.f�m�~��>%�62�G���ָ>+ur��J?�8�����O�Q��o��T���F[�RG$m҃���/Z�>2q9��q�r �Ė�\��)��F�>T۵#����S@џ:E.�O�h�����'�c�a���M�d04���Ǵ����;1�M*���t�w�zyȒ�=txZc�'0 fhmlߚ֓�K������R͏��i�h�fF?����ֵw����v��'�v��ev��3�a)����*P�g=�~�T��p��_H�4[��?���0��$h���ҿ�����e���U_���wsT�L;M�)��b�,f�q�ŔF�t���fU1��� ����7����M�*w}�%���a�9nE�惐����\v�`Î��B儲-/�guyLͲ���(���q��������|�4�[��d$o��԰猃���g��x��7@!�|�D�;IE�$H|caD������] ����14�x#��>����^���I�0]G�j�E������nk� �fq���/��o�Ć�x2=A� ��.[��/9�0�B�m��K���@�J��&M!�ΊM�V=VҸ
ؼ.�TN�!lP��m���
G�J>!]����Ut4�E�K�#�dc�����>�Nժ?�N*�1鈛�?����B�.O'9�E!4�a�).��<��i��Ɛ'Z/ԭ̡��A�#A,�4��J��]:�Tx\����~���g;���
Y?�:��s�?ChG����Ѣ�铲HP-(�mA��b��=)�D���h�_$�B��7�x���
<Jp���p�+*���f��I�%椠J?���(+��S1QY�ƹ?�r����_�?Cǥ�e��8����}&p�z�).|̆a�0��0�� �\��_��t���1|c�4�C����ԉ�>���j����r����4�4��k]?!֬�3WX���Y�3<f��GlL�f���e�����z���nR:���]�i���0��{�=�\d��G��m�������9��[�~�-Z��b�p`�.- �ZP"b�nZ�|
:hjlO4�$ b X~��n"�ݱL菼zsl��[�����g�8�:}�7�Xh�TVP������Ȼt���-�q�RZ+6�k:Rkz��@�k2b�#���<3mT�EP�Se�
����3]�6�S|@��:�1��G\ׄ����J���56+�l�oT�}�	n�{4<B\&Z�SL4���û=Cv��7�9F}���K��~q�ի�a�4�ӃFsu�n��Ph{-$$�26�c����M�H�p@p`�_:�7�u��b�p��ɟ+- ����a�0%^7)�g��Y%	ɨq���h��i%KCcF"C_F��$��f��&��xD�6O	سh8]�Z��X��N�g�4'6�1�1����Y�iv�OBI��h|Z���Vf�l��S�rX��/�\/U����^m2�h�����-�<Ms�a���Ï��D�yB��� ��  I��H�2���ښ��0�A�LR~r"���X�����zet~�f[�j���h�&����Wa�_�V�a�"�T�n]o]Xr���-5�Z]^B�� �RYT��M��m�ϖ���
u��hc~�(�{���ۣ��<�<PɣP�$ ozM�<����㸊1��V@���9���)�Ϳ�H���>��>�`�#`kF�u!�&v�M!��K�RђW�z1�Ј�h�`�m���U�-)$�J�ɥ0Gb�闹A������뾀�j� &����
�q�ب?�F8.�}���>%���7ֹ��Ao]�$'6p/�u��mc����?�����r�]�JY@�TWō���'6f/��gcI3�^1�ԵX���f�8Q��wg��.�K�V�;�\�W_�[z�ʈ˧Gn;j���Y�i au��}?�3�q���"ksi�<�W�����,S����#�j[w�"UHѰ�ILAD.��E�����?~L���F�E��
Q�
�~.��k��X�*��\)��(�b��9��b�-?��w�=����e<����z�}6�C�(���A�w��*�����T"Kt�0��7d��N3�dhF�_����"+k�
������yjr��4���A�j��t˛\j3����pb�o߻�cx�����y�L�ש�p��	
0��I���H)�T��g�(	O}��ZE##p�[��_̜Z6.V�����5��$�띀�����ӵ1�H�nلٱ��
��I;�nߖ4����6w��)8�O1��9� ��μ3�y�0��N�c۲'
�#� ����*�E�P��E��=��}�A
�nw��,<@~>���#!��Q �|�Ӌ�hv5M������1��y�-Db��롽)�P��m�_�A�h_6��j��p!��p7!�$G\)]HG/{	h�.8*��	���0���k�)e��V��OC?� �� u�H�6k(h��X9��O���	H՝�|~j����	�8S^҆�1���X�:�5��G���Qz�΁3]�W+rǨ����aC�n@��r�o����/8��߻Y�:�&�-HI�VX�P�8��ā�z�݊S��4o����Hi��!��.,*�4̒�ч��/���AÇp��>?�Aţf:��%�B]*���Ӯ�Opr�|��f^�b-P������:G�l{���q�ࢣ<g.Ճ#�j%��)��̶b#lV����4Kzk�=?B�$ƯQ	Z�����Oh"�U��^�z�勞��Q5e5b�eĳ��-�E5�����:�PwV�7��>��)*�� 4�-ƨDJ�d�� ʙI4����R0�h�g;43�0"T�|C��$юc��M���G`�4��>q^���������Z�{WB�|�ȴP��6�
@iP)L���
�ʰw����i�uq5���soe���Z1�oYD���J�{�|���<2�[��Y�Q3��F�4�/k�`}����}�� 2�J��Rue��$�.!�#?'6�D�d�EL�")��(<J���G�ƷbA��B=�Q Xά���А������[j_�ѩ,	�}%v}�����;1k0�|A%���(�%kj{�7�m
��5L���@G��9(����r�ͣi��qߴHT��.(�h�F��E�
p�{�ξ�%��лP�{�N�`�ˈ�-���K.�N�V2��6���dV�h��'�?E�L�ޥ������2���c�m��QQ<^�;��b)�Q�Lwzj%bi�Q�Hx�S5�nI��W�'O�nH�p�bz
adO���|���*�Zk1� #n"K{����NG.?e:l�u��dϥc�&���\P�?��وvx��N^Kt� l,�����Sf�n�c��X�n��F�YL�+�6/�2�4nV�m�(3�$bwG� �sݨ��E�����Ɯ��-#ϱ���Mo@-?sAu� �0l1}ȵ�7����}'��ܓ<������j� ~=ݕ���Hf�oheN�)W��9|S�9�k��n.����S��������I7Y&�M�r�ț����Ӱ��Ӊ0e���tCY����f��T��$I����{|�"�K_����N[�_}��f4���V���ʘ^�����U��RƉ��q�d��\k{�#r.l��u�s`9�A7�n6v����P����r�.<|�qz!V�D�V��� �PU�on6��S���q�n��3�G�n?�7�jk��]^ B
%�䙇��ȿ0��ŉy�4#�pN$��1�0�aM7��3��CxB��SWh�w��[�@D�K����4 �R�g���n=�흩\M�����T�,E��Z��m��)��Ơq�gZR?|֒[�C�wV�^dn*@#���V�0�������4�S5nHBEhݾ�o�Dǎ��_YAI��GDF��i:� ��Y�b:���c5�2¶�Wu�_���<��`�J�*c%iРw-�$ ��pf�0x��rmI��=!{���o��r(C+�XO��]|RZ��S��[�<�ݘ����?&�p|�O�	�tyΗ�N��b��Ѓ#���7d���%�E뮤̵�X" q����KK���e�&s=�4P�J3�:	υr����h�~�R\���#	��25p Bc��gna��M7F:��^�+��J�wρ��۳�A�Zi���.�hw[߇��m��2	w{s��;�t�l����3f������KP�VپMJ�O-l��ࡅ�WξiU��8l��&˩xr�>����H)���Z#��7��U��c>a�g%�*V�G���#�i�daYF
��z;�o�$���Oi���sA����k�V����dj�܈�\t���E��m��3�d�;�6$x�VLU�I-�^��T�Ak�~����
ze2���_�a4 ��Gu��Hѻܕ#���\s��\�I�C�y[<[>�\����?G>D�r��+��@B̩����Zó&P�N��.%2�������X�3�^�'f�����(�*��Y�E�B1�T��Ǟ����@�Y�A�r�ީ	M��}�f�F�v=�����]
$Lwf�>�[�ڙ�ç���g�:"�,�����.뼈�X�1���T&��j� \� s[�L�9�'�>0�f1�_�p��-t�ٹ�l8��ؒZ(�of� ��D\P��b����]T��F��ܒrv��,ox��@%�e�A�uɅ�Ee�L�/�A��?ȩ����d�'�&Z�|����R*'YF#DT�lD������T�(Oz��}��Ō���*e��8w6fZ���(P��S*
j�v�R_ȝ����֏�㗑LK�p��h� =��\�����N~0P`��R$�Ţ{�.���N+�-	I�J@Rl�'c+������-[TN��٢�y�1�Wv���;Ļ����ϰsl��\��U2�\�:ಶ�9�dIz����+�{�@�\᲎ ����ˇ,�Y�ٺp����qJ��5�^{�}��[��-"r+!�
y��7�-�I�_H��ճ,n��m�	`�Y�]Xz����>~9͎UF�~�=I[?$c�5��É����N�;�ߪY/NzT^r���g�פ ���t�{����⹒�'a��Lp�6)$��4������I)A�sW��&��5\�-$&ҡQ;���Ռ1�ҭ��L�n
:�C�U�c[�8ɽ��&rI�a�*K-S!Zn�ٷ�����!��S����<'�R�?������U>�
�Cz��h�3]��PYu�f�h�<��3*|�Er 9��p�U-q�.�?�������%����|�,��N� IU-v��D3A�8?��z.��۸��g0ܺ�Y��)�P�;����G��I�j*�x���ծޱ���ܯN�Q��0�\=��_��{jO]VD����4�8]�z�v1V%z��9	�dȼ��l��n������Aʿ0�˳����m5�͂Y��d_�|)��aeE�q�.����A�}%�b�ܼ,7u3�1�p��6���W�ϸ����3Dx�����Ɋ2�m��w���� ��οr,�ޅ��Z7O&;���ۘ"���KR�d]$��z
�Jl������M�/���D�U0%��&��[X-bh��tO�����zΞ>RZ�1B	�c)"Mg�K( ����V�}n��2,��G./�xV*$������4M~P�ƪL�t;r����ʿ������5��O%�:��9eVE!ܑw�d�/��]��.
d#&����!BX��y�g>k�j�8��W�+������K����e�x�7�ܣT�����VID��Dw2�R�C���83�-5�VJ�È���SU4J����Bt�54��i�IHD=�:��lx�£�!��\H�E�#&</�-�-����T�*�{@x�"dF}"��%�*&�EP�V�R�!�`9����z�-E�#?�M�W.а��z�-�Y�;ej�za#/��޼XÞ�2*��@����o�]6iEB��v���2�1�@
���c��Cg_�U[�2��dD��S����
Լl����<��s�9���CNz�&��
���'��>
���"��Qզ��`��($��웎�.Iͯ��_ }���l{~(R��^�ʫ�RiN�{�ԋz�f&��]�(�0�Tغ���Ń��G�~�)��X���qo�i'٣1��m(�V�k��{b��#�=�=�d��^DV�+*"|�*�FS��J�z(����8-@���R�� �U�cAa�?Z�H������_Bײ�H9�6������d妑R$8��#Ѥ;|2�|x�x�X�)���ӮyI3Fl+-?�kΏ@����B�W+>��4ͧKK��L�0J~ c�??��u��F��/=��*���6�n	G�G�Dռ=���`vӘ�RU�2�<�M}�B���_�R��b�����x���_]�n��|�y[Ѩ����T7�U��/�͖Jy�A���Y���#DH���ޓ��ɤhEd��]3�R��|�闪�%��%)(�%�a
k���h�����=��A2i]�l�߅a�@����������zi������$0�8m���4�E����������zQS�7��QSl��T�F�ϛ�~(�Uu3+�'lU�_�#p��2i�E��ޥN�Z�oqa�\W�e�TA�;��J S��TA��Ƌ���f�A{���D��ul8l�8`~���X��s*No�AKIF��]
�p2��<9��I���x��Z�hx���%�:��%���5�VK^^l.1^��>��<(�t�)��$�`ե�Ƴ�^�5݂�	��KJk�t/ޟ8I�ị�����.a��X`�	@�5����!��Ua�s>q!>����� Y+a	��\�e�1�����O+��"�Z4�D%��!8J��z��d-��o2Rڣ����O�����Զ6e ��ן�}��7������⇜�*~��I�j�K���PPv2jL¯T���� ���4,Xv�w�
fw�m�S��o>�5?���[�(ӂ�#��26rs9y-�����0��|�~��!Lq��\�h�4��*���Q��I��h@B(T3��m4���� ���#&lR�v��9��l���{��1��jMy��2�S�������n�ae��Ƞr��&%���e���=#�>���tQ����mz ���O(`����f2��w/���:��:���+����֔�+]���'P�x���8������g�/�}�Fv3P�m=a��V�FX�%�*.�=���bO$�E���Q2Ƙ��g��Cy�d{`�%��˼(����<2!l#,��T� k�9�D�~��\���O��$���G{1�k�T�9��zE� :�Y�@SU�܁둆ӯ�B�hf���Ĝ����TCd�.�o��#��P}F[�l}Y�/��0��j���8�C֏"|4rE�`��f�Y"�F�G�Y�mV4���F��Q6o��#˦Al�䵯�e�Fv��D���+�+�]�`�^+�|R|g�9q���-� ٺc���n�4},5��
Rڞ���f&��[�Gԣ��hj�ł�/&���7��[�v�ѽ��8t$$v�ҝW]j"��4�5sB����bNX ?�.��<�J����!�3�=0�4Oҍ��[�`�p	��7� e�qBz�o¦���n	����GA)��K�-�9��,Z��(R��Ƨ�؁H�MPJ,�9+aLG��!���
俢D>yy�T�i�S���H�2�A"m����EQD�������ÂYoy��D[j?��mXun�u-�����\Ss4Ԍ�N퉼ƥT���p�x��m���1��.��pԔ���kH|[i+��sJ68-�\��,9��X�Z$0�&�JH��/=��9VhT���Q���J�"@?.UJ��g�W����,mog �W��.g#S�h�����C 6L�S�L�����M�{��o�\�z>���d�&�;E��	`�nN8M��U��jx @�g(��:n���h���@����z�[ p��̾Tr*�%?t�j����1.��#�_T��7+�P�+c0�BƗ�n&
���?��2ݸZ �Vgf���w�p2~�d�3jh�%��;+���)����!s���a*ZEh`�1����/N�#%���޻���I��(�18���w�	�ع���'�3L�Ѧ�P�m|.]ų�(�_��=�ܷ�ŋx��
%���Ջ@����%TAd�0ʻο.��^�� �ʡ���0D96�KdF���-a ����e�p���7H�3.� M��`U�W���'�5)��'1��b�L�ZN����@��H�f�=��Ak�&�ez�4�~A]ѹ_��q�oY�e#)�WE�o��W>��<s������(jn���6���S�t�,xܼ��)�%l�oߖ (/w���6k�s����`�/jz����	��H�iB4�i��iN���Z�� :Sh�Gx�Z����j��j��{��H��vM�>���F4�`@����2��2��F>)k�Y�(������$��d$$�g�T�B��)��A�+~���V�}J�M�����,��㝀��ܥ��u��j,[Ld
(oF3���,g��<2WQ*��y�X)A�l�a/Tkˢ�R.(bR0&B��`J8���|t!����m֚�Wt0o��>��QB�XX��J�ވ��d�tQ��X(`��S5�؂�I�^�{c귨��H;��?�	}䶜MX��8& uMhB�d�� X��v��B��L���&hl�0�ʷ@�H޵��g%y&mUy1(�����ۯ��bSXw���a���ͅ)� ���ب!nW�([0���4lSj��.1���v��l+,}x��Q;�L0�.���'}���V@��
@sn8��"J�y푶��T@K`�&�[�G���[VC-�O0�Nq�+Wdۘ��Y�H2�q Z+#������2D�f{S���#q fAHʵ6��d�����k=k8��#^�%O�g��cf�|�Ç�_۔�T� I���D�M�k���H�Zjy�ʈFA���w�����U��@���Fi*�n����H�-sGwy
���f��!��p`�(7^��D��m�F�T�򤶴~���mv�\ڙJ��¢�ru5�)�@�5���G�5��"ٶT��`c���n�"�B�.LN��xy#��c�ܤm���ؚ��3�0�u)O��`�v�� K�c��-��+�i	��ʖy�I��KC���Ha�+�R�Án��ʸ�Sd�/]�04lj��.'�|ߜ!Fj�Ex���H�ߜ�	�BiI��{en��}�k�W���h����UQ��%���?�����I��¾;>C�r���y����KZ�'A�3�x�l�~��9���А��Tb}g�|D�M�O���H��O�X��nx�'\o |\�IW5���z����T���{�p���;j;!�+�:f���Am2|D9v ��bM
���޿���x~��U$��]��X�ʭ�i�"L�8�)(��SRӈÇ�焣�a��t���A�����2�z�X�G�������[������R�N�����e$5u2]�U9�x���2](S�[G���:��B���H&�:n'3�T���#l<c����ܳ�n�iQ86U`�1ql #6Dffk4�s��w��K�<�E�&��L-��R�8�Z��X���X�_������I���v�d�mo��f���N9ܧ��˅���TBM���J:�Pf�n������H)qAv��#7��^U*�F6�RW�@L�(�^�ж��M@�=]�^��|U3*;��l��р���x�>{�����Y,�4���&�~[�B�g��\�&#�c<!o�Ħ��-��p���ߑ�QQ���Br�~Fw�j �!�:#P���2��X���R?%oQl�J$�o�hЦ�n������PW3�3����;Z���,�I�mH����R��l�AJ����q����[eʃ:�;��>��S���q`�ǻ!iY��,;U�~(^�����R~h�k��P���޷V�8��{B9�.�s�E�J@@�J����L7Ǆ�upF�!��푔��k_��X>�/��?bp�]�3i�?��١�:P���(��&�r�õ060�gi?�.������e���[�)!��1I�������?Z�N��Hi�7&�����YNWR��W�^JO/n���ǧ����|��/�̓!bHS����%�ųo�x~ķI"�`\��
sm�ם`>g]��}�F�J�&�e�Ał��-?69|L2��;c������ֺ\��e�W�3ӭx���5�IV�n�'��1W��J^�ݺ��v�s��m�м�[L�8��9��F��uT���`�^Jd9�����I%��Zk=ZZ�r�N��>��a����~0"}��^ѵB����Ç�����֑�qz �#�)�hb\�#���Q4�������#S��ݾ��z��F�J��O* ��֜�\�b15]8}��hY��wJ�2.�L��]a� `EgČ�9z�|�ff9z.n2�)��v����f�I�������̪|#�Ks���/t�=YM��׉�O�;���Sp�z_���p��~����}��;��{�v|�����鳵�x�	��[@N#p����I�ҟ�l�u�9],���o�ědyX���J�}#C���:���]~�¥'��$��G/4Y,��%�]�A�q,�n�fg;�_8@Z7�##tnE#�(ti(�W�z�.�ac�������M�e1�����`�q�(�n4q#SM��,��d�*�E������ʾ�j}Z����̶�#\�A��� �����P�/��n  ]�PВL��9!�{�S�F�s`�
Q�	�$v�}�D�*N���s��A$�P琰���tZC�\�Hp��#K�3!�+��8l镍���x�-��G�n3q<T�:�%�!��$��v]����J19�a���1�`���T�����y��>z�9h��}�y�&ʠ4Q[�ۯ��َ�,g����JC&�H����׻�f|�R��H�2b̗��9�O�_R�>m���J�_�.ҫmR����'�8\ĐxZ���S�C�L�ќ�5�+~x�Ҝ�&��頊?Σ�n����"'��j�� ��a�ZB��F�ܱ����J���A��ѡTBq��-����̮�(��h"��2Z��"��,�:�|����g�yKųЍ�WX��,wl� ����YI�?׫B~���<����x�0�j����]���c��øR��d1Հ|Ipv<��w�����y���=���Y%��d��<?Y��2�(���Τ�=hq�1��>��3����!����b`N�||irR� �L ���4G6p=tC�>�����
O�?�FWKv�ޜ�8��n���s��g��r�U�]�mH��$��_=e�|.�e�ԩ� �"�d��/'�[F�����8��iZme������\�ǖ6�@]�����K��Y�j��>o�{Db������47X%ҩ�=�LV���5��悲�Q������ԌI�"����^@������&�ϵ�oZ,>T-j��m�:[/�5����Ak��\e�,�%��#`=��0Ԓ�i4������K5�k�Ժ��\h�rW:���nbzX,Dw,�UJ�Z��~��q=��X,��7U�my�r�zj�7T=g�ܭQ2��.x	m!\E�e��Cu@�/�UEm;��u�#=����2(�st�+K�d�)���dz-�j?R3}D���^�;�:G�$���|!�X��Ni#P�`j���<hah�3�ϬA��G�8"1��d=��0O�|�|��$x�d�.���F����JDpv���Ѓ�i����2��w�k����,V�Yڏfl��4b��P(�&A��N��%�2�����g�-��@Xv��&\�Ȗ��½�N�;����ZZ�ۀ%�K���8��ށ�{~/��E���]s�c�2`m�ugM_K��:�R���!J_*6P�O���0$Qd��w^z,S�b�I�i��������=��MW�z; �p�[�Zm�/��z
"wT�����eQ���C?w8�l�ne��
�*>J�;����[���Fp{ݽ����1����#r� �R��d��� ���c# Fi�8tC��{������F�6��:	�5�k�P�B�'1Ї��^�R�u<+�/Ĩ2g�"PU?��w��i<��m*0-}�T���-�~�G����w�7���^P�,ГVH,��[�eßzn�2�7��M�э��<���n�C#4V#�[ �D��_SXpCW��hjJݝ�j�h�<�`�5Z�>�<�}��5|��TfL�M��69���
,3>WB��.�K!� ��(p��Qߜ45�8̱�͵����üN!�l��f��)���F�:���^���������O3k?,�7�`�v1u�)�Q�}Ֆ:�r��r�볊�;� MC/�@y�%3�8��w)���c��=r�?�
w�Y�Y6��i(�s�~o�,�	
���T�!�����u���=��*�og�"VgDQ'��E�I��\w�&bhFX�.�_4�8ܕXbi���4��cc{��4�~'[.ۆj��NHQD�;�Lͨ�M�A���Z��'�qt�h�����X�Df�`���A���Ƃ�ݓ���F,�]*r����Ug^�._]�-��z
���4v ��F�>)~��l�x��u-Q6�6-K�������Kqj2���~��w��[QQ�Ifo���B�_���HðIRU=�,JCY�����G�1�s�����������=C�d|\��s��I�r_��nc��z�\F�Ӓ��� ���d���Z+ʘb�#�	�(RRE�f�^K1����P�kJ�ֽ28�K���
�q��N`ߘ���|�Q��F���jv�+r%X<Sw��W'w;�N��^6���28,"��ب(������5��/�U��� (�8U�Mš@у��aV&%��/���H���}'m��e
�YrF�9�5lגU�~����>��!���R,���E%��t�ҥ=��J���/JQ��.��14y%KK�z��~N��xN)K���V��_y \�A�ΔP׌n`Q�"vڌ�MQT~�H����
(�X��6(�i|��`4����`:�b�����f�*�"�fľk��z����[�O�烡BJ�E�za�y���RJ6O�z_�Ø QQd	eCez��aĜ}-�X�0�3�l�%�O�e�U�����	��):lz����9�l���=�h�̻m�{��(��T��%�&�a}��<];[xa3��a�M�b�:����dN	�0#�E�����5�ҥ��f&)��:Az�/}�-}��_�^54U�����
#_�,ss�	2+�ض��M5�Aq�w��Q��DR(/5���J�]	6�J/'#�A�pK"��8��Xqs%�w�U�WG��#�ʸ���:�a+s��_��p�/[�AO~�W��YRwc��c�n��ג���Nw���9�n��f�9*�Zhq��b�+���Zè�h����&��F�R�{�c�O�Q�8�5�����.:pY���o��
%����ܳb�p� �9]S��7���!1�	���A)F������8ÖwJ1b�iw��qF�C�I���F1УOuz���jW]3� ��"�S  ���[]�=e&Ke�r���2�ƍ����w�77Y7��n��gB�(ÿ`-�o��ޝb1X�$�5�Y}��Z����Ρ^<��ΙE�%���"Y��M�0��uNgԐ�P���Cپ�[�+H��n���:��e��ϾC��*�d���~-b��~/�?�G""�hz!jw|��?�Q��	��1�9c�F�M�4]j�A��꿿��Lsı�9�I�u:a�n���5f�j���Z���-�;�,E����z����:�o?}|Cq��Y9�d�Ì�S���n-l�uzh&��a_�ߐ��]NT<f�v-�Ua�d�9Z�+�z&�Z��Մ6i���jS��$��ze2d��Uu�����.YhoF�P����gے5d��U�IS|�#��b���)����V�=���-�]=�e \�%��&��x��{�K�eR8N6��������{q��_�!1��:Ή��`� <c���^sa�Zp�\\8��T'c|�i�%{�W��Ɗ��`��CJ�(	⇐l�`�Z>NLh͑�n�i��ՊeZ�/�F���|���Ź�G"c����F��L�&s7�]�h���Q�Nb@��K|�z�a�Apt��B��/]��|?_��5�zCh�Qä$���V�5���0�F]�y�wp�t�y� 1*�ڰ8��J��)�@H�)����a�B���i�=5��j;�����n�@�+EN+����B��Tl���	�':�܉��p�����4s%fc����Um�̵o�,������S��� X�.M�`�V��p`Z�'�#�D��l�m���/i���dD�m3/���)�G-7��8�뵲�p����q ��?��Z�kP����L��y>�-�*JO�aE�P%�������.Mf�~�X��'̓�)`����n����@F�� 7�(�0��+/�x[����f$�:��Y"� ��P_���D�B��|PxK�>�[��ݰ�4�'Z}���.���$��>=�_�8GJ�
�
��<.��I3��d�1��w�H�D�_+�Q��IG9��~���s�/d�Z���ؘ�>Bu2Ka{$J!�r�~D:�M����1j�8vdY�b�K���r�B(8�,]��&�{���`:���Bq��������JS��|���v>c�E^���S�w�t��8�z�GZwy�G+�y�@���=9�\p�I��=&sd�>��1݌�®�C�x�;���sm	B",;V�����^��/����*p3F�@ =
�$�Bt��J������E�ܶ<	Y��{̋lX����]�
K�}�,F"(�n����4}q1��v�O�z�5xǌ=����㫡��r��Q��+ad@�9o�Z�>�Zb�b�+�!e�x��z�1v9��r#r7��%�
�"l����)� !�Z\j
�n�l��M�#�w��iy�GH��?���.�[�'�u�OT)7S{w ��5�im��z.�A����n��S���u�y�uCg���@1Ծ'ŰGȊ��T֍w���.�;G�g��1���VT�'��|{���UYn]!
�T�0��W�D�d� #����Q$��W��&C�ʇ��rSK���-��T_f�&��������p�q*]Û�Ɩr~�v�C�jB]0Ŷrg(aX��4�^h7dH��[��]4��4Ꭹ5բ������ ��5O�k�d��F/�P��*�~�F*�P���EO|�J=��8ŶD
�V*(�x����i]|�c��gZ1�/l$.���c	��,�k>��}W������Qg�J��=�}�D���_v�4��A�R:� 
C��.`�ǖ����4|/�"t���->i@+#>s��Ib*q��&��Kh�L3�'<�ISN>b�O�7�����8��D�*S�ZGcU:��`��r�
����BG������v#Nx i蹮�eId�x}�%�܆��i�����9�ObxEI*��/��R��8�d-7N։�~�$��Z	$�nXC���`P,���5��U�J4�Ԋ�t�>�:��t�V��I��!n��>u���aZ@VX�T�3�3B��mݥ��<YG~\�	!nq�J�S_iC�O5�St� ���	m�����%��<�'T����+�v�̲fK���#�d�'�̅�|���O�,w�
���t����3�X�-J���YǪ�N�5ص��]�!}�v��j���x<^�L7�H-�훯�&��V���G�4�Gɒr�yT����
��?>�Ui;uc[>Z��7s�C9"�ưt�)&Faj@ �Sg�1�n�4���^����死�
P��W�iL�,�t�y5]v`1�2�x��X|�?�_N��=.��Ϙ\а�4��)9-<�?�Y���u`A�Ρ7I�0hG*���!�����FЍ���Q7�w���]�-l��p��-�Q��6�k��η������$�2���z�S����u�zb����o���o���" ����5Ge4roBw�J�-md�)��)�Gժ�l�����C�P�����wF�i��7;��>�(0���|&�?>�_�7�F��`&�݋�&���A�1(y�5�w��m���u_x�3���~�bw��;�	��0N��U� ��r�����q?�zü���˺ P
�@��P^��p���k]ƜJ���!���"�0���� �ʡ&��{��.'�Ŀտ� ��ϫ��@]x:���+̕{�Ť
J���pq�p����k�zz"�H��޽71��Mi-�u=��o�z�]��)\��f������@�z?Y��c�b�8��ے��	0\�ﻕi�T�C�1斉�[�Q
���I���D�-�hJ���I���hH������2�� V�9�rq�ɒ�*A���~4�bCϋ�NB��ӆDPa./��U3g	TEV4�
`S�_OHV��l�8**,K��]�/E�,���
g�2����;�q�Q"��^����:�?��G����O�
q�����QQ`�\����TzN4d *�=��}�,oi=���#Q�<3��a'�UǱ��.RJ�x�[���m��5�Вo�{��}�i�Or�,�;���K
��G
o�_	�[B"��_\0Jv��MeA�|��ތ)n����Շ�`�j'f�����]���a��TN�np*��j}Du�hٌ��S�ªƣ��a�޹a�m��
ȇo���Y���L���LJ)����0	���[/�,��z����98#��[��#k����X��͖���4�́�kmE:@�S��Q�o�`"$e��H�$�X��lx���Cij'�+-�����@��4$��'?�vd'��#l'O�-
t۝Ѣ�����{c;@����Vj�3lvb�Ա�d�͗�|`ڋ!p��&r���m`��5�v�A��J||����i~T7����-Z���!�1Ln�ы@�|d�5FL��LlŦG�t{�0�>#���?"h�������E��|v�?�^r `/�ʧi���%�Uy���	1��;����e�bRV���U�a�J�,.��[L|7�E�%\����1�1O���a��m)�Љ4i�vG�$Ī�C>�nx�\�q����.��j�4�>u׬��\���	�w�Є����t����}�-��}3�C%?1�h����y��HLu!�T�ohlX2IQp����(1�H��No�S&�#_V���cd�������G{��1	����#=se���`�(���3E���]�G�L��ї�FF@?v ��n](N�VIC�k������OD,�r���r�X��u���Vmч������"]�������H/u,�%>��n���L�KD�;�r/%���b�,�E������aQP%�Rf��$hg�� ���|�����F�ݾ��]���D�:ك}�a}_�L�sQ�s�y��:\^'Y�?�� !К�z��C`��ﵛ�5|���ħ
���[{�I��+�/{�j�C�A+(�"� qp�G0}ɛ��=b8��г�S(��(�r��:�_]fXA��)��R�K1�a+Vv,慌\���1�v	�?J��L� H BÀY36�(M��t��#����-/�VY�r�{��Z���,�������^�'\C�� ,h���(������m%M;+��~�p,��s � r��o�ne��QN>�0Av�41����T�Ǯ�$�_B�F�ja��BU���Z��B^�k]�:1s�����%Ս�F+�~�*���Z��o�:��i�:�#B�E���abܼ��d<�[%V�Yz��V�s����lWB4��Ƌ�� TřTG�Q�Z�q��q3��gkLy�ŹsSz#��
��)�������a�v�K��1u~���صK��{�t���T��/�]i���l6g}~�J:���"{�o��.�S��{��sSK�ڽ�����7tH��	�NT��>1�9-WC���&հ�����X���Z�M���1 �S�>n��e2���/�[�n�O�P��.��¬�o�q�aW�3�f�����$�����@�I,���և����X�IY�@%|(�С��n�%��
�8"7U.��H��^{K<r>�)�gr������أC����C�#7|V{�2I�����F���L� ��'�+��h�?M/kE�Lf�Le^�r�)m�\L�I�뛐�eo�I��N6�՞�s�t�"I>���N�Sg���ل;�:r�x'�(Q<~������ ���>U��gy7(?$t᎛D�(���Z��6���`��A��/�X]~|N��9|0\O�n�G�ߧ �6�)�M�x-���Q��ߓC?(!�'�t��XHdj�S3�I��ɘ���dv��J��hOD��k4$����3,<r�3(�W�6MT���et�ӑMGz{A�������=�+��&uϿ����
�D��3��?�� (��&V�������$�[����ax��[I_�}�i��=����v�
>�Q���x��`~��d�}��@W�Uu4OA%-�`���#uvӇ6	`�϶�`s�=����K�j�c\��hQǴ�:�P�u�U�\'���bf����ܣ@�S�3M���V҃6�����[�W3ƨ��1	dT'�6���u��k�͟�R>9�x�kt�/��� ������{9?��T�|0M�J>��yBAs��/>����^u]0:Z��rR��������
�{M6�UTod �a��H���ڕ�-v��ʡ��I�����5��F��W6Cݝ�ZYIayK�3���A�X_k+�"�x�3�ޏ�slF	bq��ca&�Z��~����ޜ�g>&�z�����XĎ�N,ͯq��}D��I�6�P�!H/��0���Cr�F����&rg��O���,���0t��G	|�[���OMy����4iG�x9���ju�ت{N�b�Fcɏf���6R�R���U�.-�m�"-�$b�/"i��ZI9�!V˟Eu��wM%��}�j�>g�
��˳��[�Լ�=s@J��0m_f�~�?E�u`�9�O3��{ĳ��e��u�G��^͌0�,�d_�
�\u~��\���a���0qm 5�O�=���@���cf��НC��B'ߣ���,`�~�B��S�[�z�c�'v3���Щ_0��{��>�J���Y������f�i�Wi����i����)��<jN7s��Rf53��L�[>�U��Rh9 g*I-g���I��������u�,��4O�A���г�k�ae(�o5>�x�����۲6�=ˈ�9�l��=�)�yw�g1J��CY��Z��1�b�z,Xsp����J���N�87_~�&o�7��G+BEt�����̀/@P%����p�:��^l5%]�f�0���hXD.�pޮ�rD��7��ʽY (\(�r�ߋ���`_�N���
��H� //�ǳH:Rׂ�΋�ʡQ��4�O�z��GF��0�`W�������H�X����aDq�\|�o�M:;�_)_�޸0A�O���>N��E�g}:0W���u�=g���2�,�`ݴ�4 �����boȓ_7$v������"�	$�X�����j�$�3:=��; �Y ���s���9��b�젏Va��k5�Z�S(���bJZ2�5e��qN��>4�	?aʞ�Y���o ���/�w���k�<IP*4W��%���U|�fa��c��:y�^��0,m��O���|��}k#uk����D[��W+Ӈ�Q�L:�zf�.
�c1�"y5֒\����R �䤰�w�\gW�
��B�a��Q�m;���7B�輪�]��y)�q*�����;�Y���@+�!���v
�����B�x��\v����hM��zaw�R���J�����~|�Y�Ԃ'�ݑ���A����8>�  ��3R7�#�Ob4m%h� �Bʆ���~9@1N=�����+�;!���u艴�j������Veج���9�'WFy�Mhc���W��W}����pC�:X�4�C�6�8���!�J��=�(�����S�o���kF�� N�<+���Ki��s�8���
��hc�(��/���4 o���ن�Q�ߡ^ݠ��aѯ?���@S�ϘV�D2y����?摍�;}�?[���D�I��(r?��!�s�r[���1�1ջ�N���|B�S.�B��:���l��Rb�f�=��,����n�ג�$ї+y���6���-'L�{$%�l�9� ��]j^���ל�Ǝm�Bϊ]DH��[Q�rv�c��N�:��lb9�A�f�(F/�����.�Z��
n>h�#n�\gC�uH���1�C�_?�U���0_X��F�*��=ѹ�eē�p���k)#I����)5[�d�ͽ���ɼy|�ST��kU��H�,n�!��O(K-���i<��P_�։¢��M�K;���I�=as�m�}�U+E z�j���FVN���.��\I��z+]N=�}D<F�8[�r�E9ζ�a=(S�s޶<���0�`�&��!�[pw��{�`R�.�|lJ{N�2�
���KHUdl	�?U[J6� �\j`�.r�rӖMO�/��N8�QVf#��:�qm;�t����}��gKP��0�eM��<-<�>;O�f��C�4���X�y�`i7=���
�n^sngX#��ukmD2��uK�P��{Gޥ���9�����j͂���rD�0���m��x�}%KN��9\����?)�Κm"$��ݒ��]�>�_�y)�;|�4��A99.ѤHۮ���K��X!��G��2ۭ���4\4$��-���o��]��n��j���
<��v��S�-�Z���GV���*B7%��t�T��L�/|�߄*d��H��4Z�3^݋��CL�|���%�_.{ׯ�T/]�w�*�R��=>2�� e%�[j�e�y�єKV��bF�߃]b��h�{�V��^�0��!*���.�Pe�3#hfe?'fD�9��@�5=����7V�7�oDCo����s'v�a�,�i���т�8����L'x$���[X�Qd�l�]!����P��b�ȃ_��5�<�{��K�J�z3�H*�nl$f�&���q�{ 1�/�ڒJ\&�ン��yv��o�����?lo+஼[��?��m^���'��l������J�X4bj<78u,�BP�Y������j�����(��cU�ns?Ph%�7Տ�53u@2c�i��-�[��&�_{{y���-	�-��7�0����VEr5[��5+��q�3:��U{�~�o>:;��<,�9�#�0��.��P����[�E,��!ՄO?���{c@�.�^C��[X��t��;>��$]u3m�I7	�����㣃�$Z�"��ܝaj��s��۩aE\d�1�#M YX%So�=^na��'D�s����N}�@���G�gA_,ޝy�c�d���C����D\k���i@$�T��������;Wg�4�����\
;���c�t�nx΂�Ls��Hɀ��1[W�a�i���NH�F��x�Aˤ΋���"n)HZWF̄�@�Q>�Z��]�@J=f:u��Z[�^&�uQ?���w탛���ݙ��?���r=�g�/[B�(dQ��@�p7ʾ��rGߩ\m�?���2�8�f+2B�Ȭg}�Sc�ϐ���r�e�c���
�i��(�N�^ȷ�H�,��<O��xV�+��B�א�bo�E̎>�%��!�'�,Xk���p����<y�z���/� �w[h.������5�S�~����o��������2�5�����wx~4���4
�ͯz�n�s��Y�9�b�Nyh-�Z�\"�D��F@ �))
����.��uV?��P>�
��X��T�jK�2X?�S~����*����ED���x)fw���tS�]s�K��@�F�ӣ��,���N,r'm�ͤe�x\�)t��WpӾ�����'x���}��E��i�rO�ӌ�T0�f�H-��W���u\|�*�kٸ�,u�8k�:�U�>����W/���ąCw��3J��/� L%�џe+f8�J���k��W}�+t��:[��� �����+�����$���MhTW��^tu���уMj�����;P��`1���o�gq�t�Y���_8�����<�I�Mgl����q5�|�^���S�9\����}��6�!{*q~g�Ɛh2���N�K���?pJy7�F��J,�Eblw�48?Y���߂�#߆��(��hI�����2Wћ��U.l��ش6�2����bj��n�և�b�$�DNZCO	To"�!�5gQgpsWCލd)���)��x��3/�7bJ5 �*�ܾ)Dq&�&�zJ�h��}������1�D'*�A��*��vs@/��H��e~��O��xʮd2�N;7c�]_��^p�U|xt~N9Q��f�5≿��Z�lz�;Z���3���q��#������˗�Gie�mӤ-��S��ɒ���aŝ�x`�t���cocl(�Ь˔c����c08.kV[�	M�k��⭣�kCs��厘 �-΍�q�C}ִH���.�6[<m�n��.��b�L��ry(�!�c+DA ��	Kɣ���=K��7+�ki)�9L�S��:�����P	|N����oB���K���X��gdUf�܂E@�~�S,^-+C��_9�MJ	e��Y����O����(P�~0t���� � \��t����e[s�Xl�
�)fG��5ei"P������E�eT9����V2�i:� �F��&.��O�kQu:k��U������!��a~��ʞ��U��h��8��bJ��������;����g�Pԫm�e����v8����~�����2�`���(D�T���� �M6r��r��9?���4$U����b���V�6Nt�տ|��0������ؼt�?��0?����Ö�I�ր�ldq5�m��)e�a�l�ʵ�S��h��<s��T�RK�,h��m	{vI���3�j9����Qσ��:��+�|�������{�33^�-m��n���xw��;%��w�B�:�k0yJ��ux����t�c$E(E����`���8uM^��N��)��(�/���g0718u�5�H��ǚ�亂F�E�:Z��w,�T� y���SD�0n�(�uq��L�{A�@i[4�별������\ME�$�Ì��-F�R�����ne����66c�|�"��06S}��p֚1��sd�>Cw��Y	�܇k�s����Ƕ�f*�m�?(����h�"[�Ic/C����)Ĵ�n��O6�+��kR"U��n-��¦b��9�5�q^9k�Μ��F8��i+�
z0��xDe��~�3�����(>�I���rX�rm�5��y0^bi�y�ɍ>uN���.jJacV2��۟�l/��P��/2�s�}/��+�xڬ��9�A����헪��X����M�������?%�������*ޅDޯ�W]�1�rF|hK��ʔ���ʁ��`�x��8���Z��>}���j�L�#�0��3J`����d�����ť���:u #1��J^���7`�2�2�ۮ?��ݢ]bbRV�q��M;�����SGg��]ܖVR#�y�8q^��[xF,Qz.Ms�_�؉�w���5γ��Y,Tr�3�ĸ��hrL"�琥�S�.)���c�Zh��U�ńuQ��*a��q��;��1;|%��WWQJZ)PJO�:��wW$��<�A��qN��9.q�n@�gG�5�Uߡ��M���V�M��皐,�{����� �N�I�v��]w{@���ޟ�iD���+�@���JY�_tͬ�y� �7����{c�$u'�K��^?Wѹ7�������0M�z��
?S���k s6���J���z"����Vy��n��dS�G���k��X?��K*`��Z����.)O�$�-A!nǉ[�P:+���M��!�-�	l�Y�g��y3�bY�ް~��`L<p&�Q�܊\�����.$;ƭ)c;������T�/��0Ly��*t��Fg�d�9S��
׳����\v�	�Kh_�B|�D,����_�Q�����M�I���_��ǈ���~�s~��g��� \�w�L�(9�]i� "c�h�Yg��1�����|�p�2��K��yW���y�0p��� ���|<
:�1�M<��i��+�$�-vm��J�^��;G����+��(�p�<�gNs��`֐Ww+��o�	���*U��hq�s�v(��XD�Uce���Z�D#q�D1~SL��n��T�M�=�"�'�k bW����uϦxD�?
ĵY�ݩݢ�#i�1�Ll��8|��hm���-c�� 
܌��PR�C�bg�"ʟ�bg˳��4C��ƨ�f��Bz$�7�Џ����o+v�����8�0�%1��ʝs�d
Ӟ��I[�Ew���#��R[���b)kC��=aL#�\rPR��~����s/}樓"rڵ�z����s���OV5
�}�j�*�Ex��|�+�� ��Q���>P��ô�-$o1$Y-IشS���R_Y��@~լ��>;�G K8'��:��,�6S[q<�!���J��*��K��6�R�c1��˩=Em"$�iQ��4R.�%�UJ&���	`�ҋ�U �hb�L��1��XS�%���f��J�qc����YC?�������N�ar�v)�����`~u
�񉐎�F�E'���q"�?�Aw(!!�➮���1���<z�o��'����+�P�-��nc8� ��s�/���=�]}��A|�f����X�-����;����0���s�_]={��hBl[&���5si�aڼű�B�A�ۤak7"�}e�6D6��+�T`S�]"����RV��X�/s��=�U����N�!�Ԟ��o.v˼�b�3������UG�vO�1Dd���f�m�%�4�"�,I����P$�1�Gj�	�{T/��5�/�MdT�����L[p���N$���\��p�:�����0q6F"��9��M�W�S�_|;�q�YA��5�R�h�:'�2z;P�U>1�W��҂z&%\ɷ� �&U���h]�p���c[f|�mD+�_�:�$�Ƹ��R8�2�ez�sZ�O���E:�__4]�0��_Ylzݢ4��S������Ԣ��C"����;�"@�4	J��$�>�kU�����߂�;荺-;���2�w����S;F�5�C!0;Xe���{�����&,Q�E�68�;9G���
�u��|���4�"tE����h�D��9b&ղ�d�s��070�W��d�k2��_�Ԧ��6]�d�� ��[��\�2�|^�u��B���uH�lHt�̥l$�o�;7fj&&@*]B���'.(@w>N��
�]����4{}L��[��v�fJY�T��H#�}�Z��U�B]��'��zW'L�k>܎�.�5VQ�3��O�i�m��t���#�|i���Y&�7��a/�M��"g K���ڧ���l�Ī�Y�yz��Z5����K86�؈&���M�9�G�і޹�Ê�.z��������[������}�