��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aЫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A'xin�XO�v⨺��sZA�R4��g�psXdm"�d��Q� N��zS��|��[{��#�r���O���J!�M��2Rm��tu�%�n����}zP�M0��>���τվb�ч8�@_�e,]��ׄQ=K��*b;�� B�
��	]��kj7�D����ш(�����c��<�MVD�ŀyQ�g���G��(����~�3?٧Ɵ+�q_�/#�Lo'�1�A&5�����P���\��@�-=�r��a�q�����ah�^��!h/pS�L<��.��>��GD�����7AMA߷�VE*������&T;�+����^���UN8�V��>f��4ō_���e7��Fe΁�h�*X��3�S5\���嚶���4��v���x��kB����%(dŬ7��Sp����k���Ʒ�q��Â� I���`�fƢ2�7�\��^g*W����!y;?�v�����垤�f�!��e\�`˞���P�6�0���2�x���`v^�}��|�pcL�I��>;WK��0��^g���͏?���ĥ�W��qD�U
,���B_v.�hb {q�>$�O��� �A�����n�E�D];UM����H�x�o��-�xW���Ɓ�T��5����<�|@/�^o%oI�C^!�'�7���Iռ"�xE�}�酼B�J��M19���;�yH��ed�L�u�)����'݄x>�Q���.�X/�G / �8�THL+���
aD��T�	S�~`���T��꫺��9/��P�9�(e�X#�����e߰8e]`vg!�v(D��j�E����s,z���?8}ѡ<zm��@?�e*J���~���dD��O���e�[0��PK�\�x0�;���I�����<2��zW���_/����R�O`8(�	$�c�|���-�M���:�	������� fn�:в\D�F�/�C�K�����t�����Řg�.�S�>^]�}&�>
�Ȍ%
��%�;e��r���'��K"]�L�m��΁��EY/u%�dI;w&Y�퓦�M��l��H�r|�Ch|
�3�|򂼆?�/Q������SB�{��+5hdJCvL�<iO��
U��X�3�u�Ra��BK��~\͗�5LY?h4܎����=�3=��Kr��?Eb8�� IǺ�1�ʓ`�tܱ�;�/�̭u:�d���]t���ĩ��C�b��d*>-�)���]{������B�M�vqt���<-�����WkI�~���6�&ڄV���ë~�£�O��.�F��X�����az��T�@����u�W3m�o��]����DR�AQ�E�6N�:�Y}���,�X���ɞ�¸*Nv��C� �L��5����gz9�*~���Ԅ��ӈB�Hgz��c��B:L�'�?�/+T��
+�ٹlz	=(��~&�/�7ґ`��ab^8��[�{�(����xPu���ǬYŞ��x#r��]�{=�>w~�^�C�<�K�#�Jp�-�e �\Rp�������˓��iT�Hth�Ǥ�d����YV�y����^���^��� *$�����