��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ��N������N���^������A�&�et����tχ�Ј�cr����9vg�w����;+�.;�g���O�;ݪ&'5͆ �.$�é�N�c �)�f��{B�� ��J�=�LM*s^��p��	�����ê���C�K�(rk���7�p;��z�c�(Ap�*Pr��Qh��֏��;f5��A�e��[�o�sxʓ���Ԋ6�=ԫгH�g���?�Y
)�N'O�Kl�������mD�g���M��r��rꖄ�U��}����4)!��q��{��	�.4�Ð�aɓ����R����Eʳ���O/�����,bޜc��Ӭy�b� �s4b�iB��ِ.&�R�[�#[�n\Z��BP��ȶ��������
� �L���Cf�iȉ21��hp��6�����	��̻�q(u$��:y�ٯ�BfW����l诂0��'1���N��֣�">G]f���R�?��Ъcٱ��M��}q��W����,V6�a��?�=�lo)g��!��ď.���>N5)��{�9�_�ө)F
!Փ�b����<1<���4U��	$߁��W�E<	��2���J����$xD�m��B���8��i$Ǡ���A�����1᷂�^!��?6�`�Tzq(R��Ɨ+�,�҆"x�Zʉ�Z��s�J�@����Y�;�E.7�
Ѭ�>ژ\�|��R���	eG���斝��� �<�ܬ0�2<�^^i�JvC��	�NP8���#����p���=�
�V�������D���+ɉ�{I��?5H�]�s���X�{�x�ϔ�4>�H��o�T9�Wç]��{�t.A��WB:b�l�#�ѷ_�8�̬-y:�Id��/�;B��<q�
�ï�iS�]Oi!��#_�G�)<�(K��|AN�c���=6�٣��77��z��@O��V�����|�br"d}��R��1�yWV��Bxݶ�k;ҵ�ʔ���<6ꍊ��F6�� �:��o�G���&Å���v�a0��KH��3���M|�������ͣʧ�e+Y��`�mE�sݩI��^�/�Ί�Y��Ɲ�1]B�c8�J,�]΄��W+�Պ�K~��^!97�R�χ5I-���'��H3�Y_k�hl��2��>�?���)���e&I�!)�`_ZB�� ���b���
�w�3%������ �t���h���ew\f)ĕ�7o	$�t�W�Jo��B���g�w	�edW x�q�WU�
�º�׎�T���_[���j����ߥpf���F��o/��?�wDm���,5QW��ۨ��sh'��.ꇀ�|�w��PkZB�N��.YsA�%4*:�{c�X���t 6Ţ0]��L�������F��=��4����<�$Y�.�q�6���%����}�܆��J��~'N� �?JXI��v:���1�{�����g�xL�k�%(3�k�K��|�3=k���iss����3�/�<B����G�����!Ot����Rֆ��6�7저��$����4���V:UL�P�˷ךy==+0�L�H�4�~	��9�AS�+�~���@��r4��q�n'�j�<T��CX+���.7��}���P�*�Ɏ�%#fh�.݊��2F�^v̇��!B��j�F���/�PG��߶�!�+�u*�&04E�7:��8�ڿ�ɥ�E>�/�f�S&x�P��H��q�UQH����g�H!{���?���-�����Z����X�;b(oG�H����
Պ��Kذ��2%�)­�ͮ�^��	��7�#By�����!}����Q��j/���Å���H<�Πc���V뗘����M��<N-�J�P]�5UL+�ѱJ6��s(��[���w�����K8��t�@��:5m7�0�IFݳ�mՑ�s|�����8M�.�$1z�o'��M���{̏�d�H�h���	����sk�(!(iċ�!�y�IXnh�&�Q�o!ik@�Uy�4@o����Fk���Qd1#�h4������T���K({�U�����12�_�+�QP�%'ḋ�EƭU��XCrB���n	KA�6%	�w|.xo-U?��,Hs�兜\��4��=�t q�d��5�u`K��F�mc���3o��d�ȧ�-�Kvɾմj�?��W����!��;�cH/#z�ܸM���]1�E�ud7ݣN�f�N��2*r���eX�pa�+�����}��6�̟H��iQ�R� �90���o���l�$Y���L�Fɿ�질$Ѓ��J?ZΙ�;������f��0y�$���_�֑.9l5��T4�w,���(i�x*~�E����n�ms��v��b��n؛r�n�$�nXa����8q�!^$�6_��������{��H͢���6n�����#ȦOs�ʓ��k��x2��IrU	��=��d��5�7�]9�"ءA�WOJ�JJ��Q���.� ��;WIU����V#(��R�y ���1H��f9�0ݝU�lTa��>����=����l�9C�xqϓ��ٚk'��ͽ:�!�8�Mw����b�XQǂBv���T�l��VD��C{�����b�h� g��1b�2�o�9�P�WhPT�y͊�4�~7�ڑj������'�$�ے�����Z�Z!mЃh�����Ic�1�LsN8D��^hZ���>��[9/ �G1����v�^��,LP�?rb�B�ޚ��:��(X!���p1M ����+���6�K�+2�=D@p+�h�UM(Z�)3�)�1L�����aRY�}�<���疣1v}.�%���f14ޏ[3xap`�L!Ì��t�=g��@cz|�ŗ0���������?ZWc�^k`��(�j�����yu�����2�z҆9))�>��+/g��I��ב�Y/M�D\�'��J�:�^V����6IOx�,�Z�_���7�>���,�.�r�cU�}����h~�5g<\��+�ˉ.TE^>ds�h�:�m�RR�$�����:�/ɗ�K�B!�X�߷�+�ftND��[E�С�s����.��1���v\&:k�E�OFF1�JJCBO��w'��:�Ue�_�sEXُF�)�yy"�e�E�	�QhG�f�˷�VQH^�;T3͇��q9����%s'��ۧŠ��D�C����Z���������[A���LXi�o����N�´9�<�ޢh8TC"�ݙ�
�-i���"�ǩ�+_hv�s�P��U�����5֠<&`Z�+�z���A��Q����e�/X:˿�����`xd�<��,�P��,L_,Ci�y�Kb���|�<��ra4J��D�w�Dp�)KD8��Q^7�)r㩙�$�eL��T��L®��&� m;W;�5�>��+2����g��q�m�GA��B�m��3C�|�{�|F�u*���,�.�=2����V\��6�PZF٤�N��� B7zŃ7��l��d�Qe t^,n�L��:g$��^*Q�R=�I휇+���i�$ߵ�GE�\���N�_Ʋ�:�"��p�]M����R➮+�/p��x�R���d �34��������l�d$�{}�N�b�>�_��ڢm1��V�Qe���gv�*��@:;n��Iq,�vU���3$��_�MO}+��ߚ���{�@�E&�s������^�:a�5d��l�+�CdX�t��څ���N�I>�/���k,5q�2���>;��d�AX����u[*
>����L�Ѐ3�M4t�
#�����/�t����l9�Β%��_Sjм��=� A߄auf�S�*e�8��=�_ڻz���ћˈ	fGAWY��!�x�^���j[I�慮_�8X�|d�	Ώu�Y�\�wufp+�-U"�or��s�t�3��l9�H��Y=O���C�������ƴŷ>�럔���	�C?����>����1����w4'8�v��I}�,z�JK�Hh���e�؏����.�D�7e܁dy[ہ���(K�2����[E7�c��[���|����Ok�l�Ί�![j��#dx�^B4�R�V��$�F�j�D����)L�!0�8�����.
?c��f�),?���g���[����[@go`�bI�+��[}3���s��|�W��&��v�՟H����np.hc8����i�+��� ������lmȐ��^��#��E��x�a��6a0S�
���w�\��)��/��gU
�N.�SqPj|���LJA�X�x�l��m�q@@U��3�"T�r�>v�}ݥ��3 �����ح��PmKޞ�ʵ��Սo��f,	
���w�x�\�����:�`w�:J1�syJ�A[{���l1�(��u�(��z,���cHWb��j�`�HP�b�W�E|�Pj��4�d���cq��)�:5��4h��1�s�.C^����oJ~�c��ң�A���7�S�����?�Μ��˯��1���?��{�'�0�ar�A��;�`1MU؇�d�5ւ����0�'ad�\;W��h�-�0���Vla�N���P�w�ﯙa�C1Q���3�'����t�C\%ȵ�����qk-��D�Uqվ�#��r �5w#ۛQۦ�"6^��>B�f��A#����	ّ��I�uF`�e9�%�u�
�Y���b��-E2����C�~<���9G)���ʢ Z_,D8������D0(����|�Ƿ`����,B�wT�*v��Iާ��")Bn򈂇���7(��'�'��Xzx��U�U���y��R�@(�8[_��)t���&%z�h�,Ӌ�zP�W#vHF/�LW��e�6���������d�R4(Rn#D7�6�N�݈0Rr��h�Y�$Tn-(U�3�_�J%���蠸�=�߽_|��Ճ�۴�yj*2�^����u7+��2�n��rK;���!r�_��Q8!��QgˠN������8F8m��Ӱ��Q<2��X�5�[J��4�sߢ�'����$MG��hy����*r�m�R�\��Ѭ�����8>�˺��NV{-j��-��؁[WB�%�v	E�~5������#�܃�)E���k���n������hm�--����!��t�șqΊ̴�o�O�D]]�<���V?/���2Xj�S_�2�y�qk���M	��eH�O^PǷ��![lʲsyֻmY?����D(��Jg-A�6� �@&��b
�G��-���������H�[>@�2stW���Z9��3h�ս�]�Q���Tb�&c�q�@�m����H����g�q�S��DȜ��G��zO>)�9���Z���m�[���'�]k��+Ƅ�����z:LıҮH֥: O^��,Ŋ QfZ���i�Z�)h��R����t���3>�^DlQz6o���8s���5�����z,�n��\Ͼ�b�*By��XB╱�Z�d����˝�N��C#�>��O|i]W�$�	&��&����^�V�e��*E���d�A��%KX��(b�t�aZ�,aT_������mI�Pg��kLu�K�� ^�Ol�	����YHL��K0G�HH%f'�U�Cd���kgJ0k�T��F�@���djM��+���=�Ά&�X>=tU��hẂ�r@Æ�����~�?�g�x�?C0��p���Nm�ߡ��آ�L�ٻ�!�n�I�nYϺq7ohz�{O��������慺:���,���"��v��e?E^�^�^Xq��� >�q�g�N�l��IN�X��};�󱕯`g�Lw���)�5�����xmZ�y��`AgX���WE��vL��@�G��/ %*�K���Q;�*b?A1S�m.�3h�mKLz!��
|)̾1 ���_�7�gZ�!��*VYduF�߂۝�)7��bi��쨐]i�3��NʆQ���i���TAw���?FU�����N��J%�aW���&q~i�<
��Ɖ�����?Q�!/�Q���
�/���w����0�%�hd���H�k���:5;�$b���YI�@fP�:��5j��$/F�)?Z$�nѧ�B�B�xR��ۊ�6,Zȋ�mn"������m꒺���6����hvAQ�g���0W�N1:�k��Ht+<]n�GZm��h�X?W��#������8�Df �!��	KS!�0�7El�U�j�G��m̏c��=2�rݢ�*�:]1���-ڲ�GQ��ʪ*�gx��1�"J�y�_Y*K��׼�� <O�1��Q{w�oδ�]N��'l_��
Iz�vm�H�dkl�U�i��ȤD�SI�`ٸ�p���TL�I��6f4Ѿ�*Cц�x$� ���b1PI/F�ߢ��ll����	�p�i�n���>XB�m \1�L#����h�������Ԛ�t"7�=���HZ�(5��ڪ�N¸�<<����CNE�"_�0Q���I��}F��VU%E�_S��A.l�s/$l*��b�1�-M�SX��4n�1�*)_�D��d׈��s'�X�0d/	S����,�y��++���CZ��H��Iy�*�М?�]��L�!���z���=UReZm�L���!�xS�3��<TZ�g��~�."#�MS>¤�(�W�J��d^c�*Ǉ{̨S�����iffԓ���X���I���D�Q��|��X����Aq�v%�gV)��>j�(�HW召"x�����S�yg�3?�
�7��F��c��?%�H'N�8�dY�S�,+UtQA��m�j������K}ൺ~x�G�bC��h�9���Bj�0��LΘn���c���/�oT*����R�.a4o<��P�hN�����n�?ԝ��b����fm�tk:Y�⯶�p郤��F�?��i��ō���&Yp,T��t�"ş��J��h�'F�h6�������[��z4�k����KGֵ��+Sb�6��K�/��Cp�OZ���e �p�0F��Qt$��64$��dV��لF.�X�����U�H�7`{�R�rv�(�Áw-5�-,>u�|�������-w�R�M�3qBF�\Q��w�V6`(:�q�1)"�(쌼Ͻ1C�By쩣��+h�=�r!<:�~XMk� }��Ȍ�ۺ�<� o�d|��Bwb�+�#/�g���ci�2v�f��� S��;;��<�q[�y��ļM�o���"r���E�lT�uz�5�&��}�o�U�����z�O�91ƿR�VS����'�+�C̝�6{v���S;x�#/Nwa �x�������cm���;֩a�KT�*����-���C�gU�墭��hٽ���Y�Rn��[y��׊E&}���⡦�����~���Ҋ��4����81�{,�P.E�e���!UE�j�})�p��6��)t�·�uTl���tC�eJ��4T�#��������A�q99����!�{��@�bW�I%���W8؆^�m;^L�.M ����'�U����J��aI�=>W����	��+'^�4C��W@� bJ��t�7h�j�'*V��Lcng ��8�c�	{\3�`CJ��%���-�q����"�5�S�����G�ÚC"{t�S�*Y��k�}#)�, z8��#MD�M�8cY�\�Ol��̢4b�*@��8�F�'=!��������Vikn�[0gOW��N$�/�M���O/'�"�2aߟ��PX:�鄾]%���Y���zӐ\EN�� Y*Gf�C9���ll��$����?/�� Qy+�ۃ���^�}ސ�z|e��\�$`I^��gܵ&�	�1J��uM�x�Co����:8��Zu��¼�}#x��l��Ocb���PU$G�P��Syo��NK��(�Ax��q\��%I�;=�Fy��="���
1Sp�NH��NA��ј���A-u�]+���O�]d���t�XXw��os���ϐ��UD7ӂN3��;���#L	$s<U+���|�$���\+���8�h�����t�;@R�n�ڴki�hc�������+<(Z�y��4�������Y+ ]s���ia_�{�}+(fI(��J�z
l�DE������bh�s</=�t"I?�V_�����廒1(�Β�а�|�J��UnN�����m��U*v�!Y%�/�/ݰy���B���6;��=���@�^��M&�
�%�9+�ϑiY?J�npv4��9��LC �I�{���[N���$�.�;%��b*��`��pJ�6U%���
G��k`m�\.V��	O��l��b���O����ԋ��K�|�Q/`��v�C��:�U֣�^C��4�7��׫���gk��DlUɑuD�s��zM�b�g�b�2�L!��.ކ?0	�,���/t����8�oˏ�d/M�4|ߙ�.l�:�����{B2�Y�K��ϗ��s��nfĜMB����G
ge�3R�(���Q�V�P�[�J[�5B=�sR:��sܕb
�����f>ɽv���Pcq�$!�����)ک�i(!�UF���쒊�hf��n������ԏ�&/���F�M�7l���
��KX��1~ܻe�,g��:���"+p�����# d���oWP�W��
�m����l���c���f�طX��H��g�-j�ZQ7��8���V��,�7T��ƫʣӣ��s���4_p�P�-����B�6e�'0`֒�<�O��]��'l�ĉ�o��Zz2�.m���x�&I4@�N |�_�k�
ڕ�,���b��Y�	8zlMgB[>�<I����DR�N���`C�7)P������6h�[>A����4��<{7	�N\�0�2k�l(�L~��P��fiHCD���p)�Q�i��/_h�-�����b��k�4��Ms��b��8��6~-J}_aS����r9$�b+w�Ipq��`l7J���.����m�'{�-cH�GχV��m��J`������
J@h�0�
��N1��1�	��~K�7mr�~�r��K-wV8��[�?�n���CE�����~�Z� �y�ҝ�_7<��:t�n���(���1�D��KĚakF���3N����Ԯ��QH`���'�mZ�Ѡ4�1	�R���^My��C�	�Oty�ՙC	�h�����49�&Bn���\��g�O�u�s�z�no�<�W\�Z�[�tR>�nAg�b竫���6��!�W]zR�m�c=`{ ^+}KI���p�KS7��n��2A�,��."�;�xu�	k�ɽ�E')�Ia��v�L.���� �|�6އ�9Lp���;�sk�`Ú(��۵���_�i^��|��\g��l�0����k�$�r��CLt�� i;qCVH����J��1Fa�cd��o�ZPU�{}[�ʕQ���J�qtC�o�0O%@I �^)�g<J�y�z�$OYk7�������|���m}���c2����Y�%�<��9����!7��c�
	~� c�AP?F��H�i`�c>�?Јszo����d�3��0gc�53��O��ȲHG$H��z�g�Y�����9�=�N�z.��t�����!���V>a�L��''�*ߢW>������A�]\޿mĕ��-����S5/�`x�b�Ataa��-[L̩�~i�%	�1pa��̔�����2��<�����\��U��}�����SAP�X%�2b�0�Pž�Ȁ��6PU��45�8�����sDvr�y,�fR��ٷ
2QY��l9F%���g*J��d ��|.��DO}��I�wۚ(��'o^F�y1l�+��* }qg��$KO�f��+�D�ҼPA�7B����L64��� ̕����T�)�c\��:�$T OԘ=�+��������/�?�!j��}����Je��?q7쩟4��� ������UR��,�o��A�1��y��t��H0�g ��b��� 2T��HD@�M[y��v�g'�3���[uz���q~��ˑ�y��É��8�n��U��VA��2�ݝ$�����N�yCS��"� �a��X�x�?ޏ�Tx�1U���JȖ�v�~��e͖�!f0|�M���N���ZA��Y���/͗�A���4����;;�|�c�_���*��!G�M��~&퓟�g�����%�2J/Ҡ_�d��8�K�z��3_ ]���
��[^��W��16`WE<*|V.uLIA!٧��+��6'���$&��L�Ot�<u�#r����ϺG5� 
���
|lE�}�9i��0���>.�v`�e;N�A���A�2n[o��;�hJj"X��YAڄ��yO�*�o#���$z��� �fN��-ЍG����L�A�c�.���@ �G��[< P�h���7¸����JѻC���sژ���~��T�Ȟ�$�$�?���g~��0�ܹ҂`t�j f䁠1��ު�aq�c��ϺpcP^�92�,�K�i6}��]V΁dzW6s��ޛ��g�gan�YK�m�$g�PAgb,��9'���AR�BԿW�A�a�j�
�AP��ՠ#6ԑ�©�e+X��!��DB���]ƇbP�	&��S@�SD?�My~�<ٳ*dF,���I1�Ā��e]���:��|z׹�[��1i�H�]Bs�|�[Q��7n����t�>�TJ�Gt,�����M�Ug�	y��v�;F��W��i�?i�
.��@���k������:�!�L�]gD�_?7�i�	1~���d�1��Ķ|�5jk���o��t�������g�G!\`;2f��T&���4�_�=J��~`�	 ��z�
���\��!c�N(DVݻ��6�t�#�>쿐�w�H��[�o4����yvǰ�QE�o��߻��d��(z��d�&�]e;�b2�I��9g���_r�-�s�F+�ΝU�a����TDY�~���g}��?"��6߈���n�`[��kx�����T�Q��h�?k�d������DiS볚uS���]�f>�e�DL%E�<�-�Bid>&dt��+����p�!���5�p;���:�p�
#q�̢m�J} З���Tu�ю~ٕ{���e�^X�[�/o��SI%xJ�W���-����D�7�~/�ט��Pl��u#�_ɁLV���"�Ct��"�̴T�k�'F���HczZpZ��=�B�Z!��
�;�@���}�\��Q��8�2{�v���I��?����B�F9���+F�$
�Z�g�fMz|�JI�p� �o�s(����;5+4E�����,�?�I'�Q1�5�w�y�L���2d�}��s �ea�C��|� � ɇ(��;=p����5�p�ä��Ȫ��Q�]}���4�$�6�I�����	`���Jb�t��7�^
�{M��e��GL�c!�����E"d�؋u'd�]�dt�S��<ܕ�6!h�&&7PEѸܙ��Ҕ0��Ñ�YE���Ш��2��l�M w#sH�/��-1$Q(�^%#5,����>���Ո�����t��Z���5�U?,�B)�`�)���*��	��2i�]H�7���ݕ�7������b��>>�
�K�я@�3�ך��S`�
��Q�|��?q>�D��6׶Ֆ�M��M	��=(s�6�W�4��������)� (�$�،N�|_�w�t��Q�9t����b����?Jaw(�wz\K����q��B(�d:���	���:=+��U%���d�tʉj���]tO��{��F h&`�#t'Ǌa�<l24_8����d -��3�<��h������5��� ��-�����F ��ގ�;�anZ��l8�w�{��4�������Z����Ud�����n�G�hG�o4]_��߿>�L�u^$R�9��bX}��.�	iԸoU�5��\^ )�j���\�,��O�b0�1�/�a/���O���b4@oǛL!��A�.j��Q��.y�#}�ה��*�8�ڳ��Q��IS�,W\_%��%���|&��9݌$*"ʹX�(���!�ά]9��t������1A�0��Ȼ��v$"����y/�Mx&9���%�J
�s����7ʐ�5I�цH�n3�9��.����kD~w>��ѥ��=CP?;��p��D�9�Eȃ�$�F� n�v= 4��Z��}�ۉW���_�Kԭ���E*�[Q���5���:ja-��w�1�x=]���A�d����ʈy��1��L�m_tx;�]�Ѱ&��j-��Y�Q���杴U)�oE7�1�l_|�d�WѴH\�����D�Qz�l�Bi�߻/:�] Yd@턲�"ה��Λ�0���N�M�	=���:������/@����>{ĭ�ک}!�o7��R���g>�ҢDO(cc��.�Zr�n/]�-,�a�<�9Q�CG��뭐kl~�Z�R�Qz��=6|�c���=��-���[�����\�B��-hX�P�+�%|J�TP7c�K��>����v��<�cܒqvm�N;�ܩd�x/,6(�r~���G]zH���]t��|��^v(�/-���ŧފu�����`��	�P���.{Gi�Da᳖@���xU5���B��#1����<�V�K�\�R�l�m�ca^P0LB�%\�N[m��Q�D'�b]��2O�)�����K4�H��e�t^�D��&	q���jE)��s�4���բ0��_����CP7C��vy#s���n*��������\�G���sL@���N��]\գb�J�3��n��5q�Le58OC�P���b��0��ʑ#2;k;%�C�r�L�K����$GQв�����9���5�J�O�/�zE����D܎��h���ʴ;-�W�f�VR�{"͂pr8��*�-4��@Wxץ��_��lOO���M��}΅p9���������้��żW�fzu�y=�-�Th�ڐ��9p8�U1P��N`��8���yS�w�N�z�����DQ�?�]�F��sV��$ΎX�f�h�﹧��b���l�~�b�u�,o!��bm$4�W������ex�������^J������6�P�=?�%���+XzTϬ�f!_�J�����?�1i��u���'MBJt�p�-ni��dz����a���6�������i��J����7~���^�<>�2	��sd�o[P,I�(�fpE���P����鈃붸%��@���f�{�F CI�;<�eՄ#x1�����������s���d���W���ݽ�.̪�����������S㺢�l(2G���,I��:��nE�|�R�j���xc[Y.�V��:s�%��}5�̻�찬'���$Y���)F�@S�� y�)��Da���Rް���sBe��`�t+���ް�a�;A�,�yy?��}1z���&��=>hKS��a�J�Q ��0��:��(�#ژq@%o"�Qh�g���y�Y�0�������F�M������p�U�'Z;��F�꼶��Om�~9� -�u"|�ΣA�Dpi$�u��چ;w ���}Z����J����WüRp��}�!6U�#5P�=w|bN����/�����ɒj��V�K��E�W%��G	"\0�<Y�|v��|k�I;�{�3��F�9�16�f�������v�x�)nҥed��0�gx�l���F�-E="��Q�G?�=ü��Q�����9�Y+r4�$�U87�E=<�U-+���迈j��~�`��׋?x�EL�[�􇲊�r��Xp��~��Y"�>?#�����/�'Y���⵿`0�4�����O1�	���f���Q����S6az�
dʩ�]������D������Eֶ�@�z�x]'�vkC¢Fh[tϒ47��j�e��!�J�����~�Q��V�����Ǥ<f9Df!��*��YRx����� g���:���{n��%N������(E��d �^EuM��Q���b9�C���8_i�M�Y�k��9l�)�K�V}we�}��/8�]Jp�sZ�}��n��{�P�~����BM�d6�[�et�n]�x;�� �2�F�f@�>+�!�H�7麆8gN�Ϳ�M*|%�1Ԭ��jM�^$q�N:�R���c���%r�#-4h�Sc��oA�gq#�V?�m��{��D��؈����ܯ�n�!a��|�;Ca�i5`��'#���}4�/����{t�'�Fяl�X�2��-�b�b8u8�j5e�p���zDkm��;e)��1-f�>e�mޡ���W���Ĩ?�A����4i��J��J�j2Ђ`<tb�hI��XZ}" R����	d�Jp<��*���?�m�2��ӷ���V]���v�9��>�pA?ɻ�h�(}Ҋ������.�,���mNT&�Ylk��04�!��BԀ/x b5����1B_ 7'�8�u������(�6v�]���R}���$��lM�L�8E��-�<;�=�ؗƇ���O������ۇ=g�B�K��l$��Eӆ�?�Џ��,a�f�)l���~T#8w�T�\Z܈XkX��R���Jdּ��,�7;g���`P�� O��`H��a_m!`BH��D�ا�s��ŔL뙶%֌��ɗds)�Nue��8smFb�	i����k�5-��-�w��዗ւy��U�&9A���X���6G-�}$x�) <�| ��$ukc{�3�y��E����e��"����o�b�=�搛m�$_{[�ۿ��LQ		�`��^�N�����XI��48@UcRY3F�{���2>>�S�w��V�@���6r���40�ؖ�e�����_C�5�`�oN6.�{�gd?R�j�Ɗ�`$N.�0�a&�U�IE�ښӅP�o]�s8U�@�e�A��O�XB��k��?R��K�FGo��"��4��q���;e���|k�������a��/�$0ɘ���xU�_Y����Vr�veFH�9���nK#��x��n�,��<G-��Z�1��\9	/�dG�@Y(�G��&�� ����|8�֔���F%d7����Зv�PA�$s�o���7xQ��+� I��(/1O�H���wVu�3�s�>�b���Q*w��T}���S��?�g��_j`e���>��v�Ț �GMoZX��^�Ai�A���E�X\����G���<��&��8����?wa3:׶���o��X�G���;o*�5@0=�=�U�s��Lã��4�:�dϾ��S+�C>X`|�qe;O��y*'_c3G��*��h7�e�HC���<A#��?��;_��'�1�J�� m�|�2 ���g
>lM����vm�7��X�b�ܼ�nx��)d�-�c��~Zr�Epcks��� ���W���N�\�g�-;�MW���,�?M�O�M$���W��4�d��`
�o�=��B�2��%���$�B���AŔ�l�����O�V��C�]U*_G���T\�E����x�[Cv@I�b�ܫ4t��b��� lY�'��p������4�*��
��e<i���K�����" CR!�/��vǔ꓎%i.j<>���r.���������5q��9u������Zqآ��3� �}���0�n�ޯ���f+�ϻPbM�a^���Pk��Q��	d�T���;m�/��Y���n M(|�� �>:X����#�s�Kڌ>.�KZ?�,�PG��kQ���!��C��1��0�莝	����z�=�R2 ���(t_��4
�6̸�wX�#��݌�T@�S��h��s�z�'��
�4P8�d�#ÑwT����ʖ%��c�I�V�w����HU?�c��7�������1)Idw���_u����9������G�
��զ��ٍ�Rn����[sg5�1T�������v�� ���ј�)?����p�V�c�<{��B_���/e��el�G�v�K�`EZ��6h�c������D���f�*0^f���Z1Q�0&3(�=7�p�y�@4��2�~Z��%By*ee�) ʣ�����|X�w�$�	 �oLU�)���TG����p盛!�[Kը9�ݛjm=�������np�j,���F���P�~)�XYcC@�s�#z�R��8Z90A��6�yQܰ�����wA���K~�Q��� u�E�G��i�Y~�x���k�B� x �oNV�7C����=��Rr�hϔ�	�n���eV��=��d}�9{@w�>�(�>q���/?=c��;d!̌~���,�8 51�r	p�u�@9��+�Dy3��6/��*O�NO�QO�$����Dq���}]�.&e+�m~�5T�6���ޣ�#�d�ug����G�?��
Н�5;
������5�i�Eu������CՖ})`�����:��OJ㽶W@^j��`8�O
��;�U�u)��	\E'ۉ�3.~�?���w�n��]܃��<u��C�cMJ�UO��1%��D�յ�Z�阦]����p��*e�J�^%�+��Q�ڲ*��j�B�m��g;��������+*�n�1N�ߦ�n�,�2׺�5�1dI����h��~���	���5�B&�=���G��_��H��;�?Lв�S���.���Y���m	=�ѱ+�G��������+��q,�A��ηW%W��l���AV�}�y�섋ʵ��$ha��?/Y�B(���b*�%����)��|v�,�����0hˇ���.fr��~�s1ҝwd#r��yN%�[�i/�l�b�h��4�7x�.U���Jo��%\���� �v���l�K\{�"̫��p�0����ٟ��R!�{q��'�)�#u-7�n ����*�9t�"j܄���3���x>�=�l�����jW�/
�yk�����ö�	�����mS�e�� S�C�;���MY�a�X5j��Ƀ�7SdOޙ����q�H��ʨ��]2k������v�+Z^l���Υ�	�f���E`�U;�{����=!S4Wf�ҧ���hϦmxp�>r@K�lF�V�{���Zy�۴�Lﲗ���E�Meu!Bxz_6����Ź���h�q�����ꫩ�I&�k�{uz���;�cΪB�N3��*c����OG�I�9�B�uѝ������̀*��vM�QSAl���@����I�U�]l�� �'���6�����F��( G�� �hK1�I뗏�� �_��LFs4���ݍ!	��o��wT,�_(2>�>3�꺼N9�?�?W��������_�N� .�g{d��+ѽ�{��N)���6?�Čs�#�_�}����ŠJZя��9J�\:��ң��S�	��O�ֲ�R����`�D�.C;8V�d������2n`��J�`����3-MhYK!�|m#�r; Š�)��3�c�	'�~to�"�%1��E�X^���/�;�05ǟ���ߵ�bO�btԏ'������>ԥ�o�}�A�$�,�]�ȱ��LPHrp��y��n��;��;�E82c�c�3k�M��];58��6��+`@Z��rRPz �=����vDn���eA�A��yș�r_%`O���P�� ɧ��]����#Q���
 �
��
�ۢ��kx���?��\&x;9��t��
e�V�������@�cհ��'#���&��N�^mx4z잝$���H���@y�Q���?  ;uf�s��"��x�p���<>4t�OxH6�b9�e�3�K��k+�k��8K��%e�2�5j��,:�m��WP�[4��&��`k!�@���U��yL����v�k�MDf^)�mb��q"b��+yă'I�7zHP�0U��� nY�nu��f%�T`'ɥ���-Aq§��DH��$,�YXxm�C�T��J�6؆ގ(�`يY���̠	��Rހb�yM�L��� �d��rYR����3�KZ^/!��df�Rz�Gh)��^J�� ��\]�,��75��Oj��*Y�]��'��#�݁�_{�EJ��W)*��0��L�@Ս��|�x:�g5�5'���T�
���1�4�܊�oW�t6ߓ6�Q^�׮�e��o�2�ywpe�D�C�O��m��/E�֘ӹ0�m`P ��v�����y� �Q�@
|��{ؗ=Tr�������0�ֺ��r�%YŦ�F!]��t��R�*���,ܼK���R��?P�]G�j8�[`b��f0��[������
�Zi��j��?�<�������y��d;��#��9�na��I�J�ߐ������7Y�l�@��i�C�~9��9s�̷n�����N�.|�w
��ҍ��f!J�q�-�.7{,�]?���h�*����c��Wl/�{���帶�S�FX�g�)s=k'a�B�Bl\���qO�p���!G�R�x�Uj�Kk�i9��� 4�wa�3rh�}kSF�"�����6�����%��G	���m�S���u=��p�ݒ��B,\�YH|m*wm��ZT�:z箆����5W�͔Y����M��CUa+@&��:6�C�i"�"���h�ErBcg�8:/pe"^�f�g�2d	@9���kq��Y<yVc
w�%�A���K\����"�s�W/�?�)�aE&�E-A��3+Y�tC��{)P�"��;=�	O��x��:���^0����~�������`[ p�j9�mP���UTP��]/=%�g�M����@�t[|�r`]�W���FVAQ�e��[��|(��U1j�(CA1��۪w����`
�r�2��'PMͬAfM<)(oM#X����΢�n#�],���H��e��8z����6�����醰�� u��<�+p�	���ՠb�s�4[V���@Ǭ��1 �o`�3���[	�($�a]B�0+k�:�o.�=*vH8Kڀ	�]��B|�$�c��c�]�l舳"�赊M"�1JD棄E��ٴ*	HVBG�ݿ+���C*S..hZNŸ�L���0n�賜�"z�� Vh�o���]z�Iw�=cH�=��oS���v۩�3�J>�8��$�o��sq�	U>���c��N��7�Yr������aG�3�_�9�C]�r?��[K�:��t�Q؂�I8�t˹�.���h\�����S�>���E?7\���uS�	�`���J�m��3 �opw�7������������*��f�?D�>fdL�P4'��V��l����]�n�Ti��W� Ա�Z�f�-��4�n�Ѯ��´�B�%"/�D��w��:�I�&�'��N	�m�ކ��*ͦ(��h��	����I�^��8�Ds�` �Uv��
?��2����/!�L9��V�pf��Vo��97��b�#]�ٱeK><n5��,/���;�g��?D�3"���_~�m5�h&O�Y�9�51��A0Nd��{���~9��u�����s������'��g�CZDD����wqY
�b�Ds��N�����Ao�w�d\
�+�n��R��Z�5������`hTG_=�H5Y�Oe1�F2�4���?��ĥ4S��X�xKRyl[ �R;̧6����S��d1����(=I��A�ZVJ��\�YM0�/��k�D�
V�H>}��~�àNēثH%���w�s�+�Ygq��R3QyKc�dWE�����$�*C�#u(�@���Qj��Kȇ-8\�(������h_&٦'b'��xК�/H�����	dC�����f�ZGVTd�X�qWN����bu��*oN4'�B���S���`�Z�CjOy����	o�xz�,�YgH/�@��o�Xe�7�F�k��<��a��R7jpC�C�#K�����B&"K~R���F�j]H%��U�\w���9��e�@A;$��&�E3�um\f��b��I��<��,Q.a�U�c�Q@?w$�,�ʉw�ٴzVx�jZ����D��q��^��j$Ҭi�K���$�%�G�Py�� n�����[�T�2b,0���W�f�+fZ'v���B�JV�WQL�D\[��h-���ӧ�)���@R�z߉��>Q�Į�!�Sn
����r^�S��DB���y������޾�>� ���j)5V�X
$��0�Fچ
�+BK"9_�m�s��(d7��QcT�g<��wulM�$��w�٫�#�e֘�C�nɦ��������)��Y0}��?����.}���v�;o���������PWG�I"/��a`������p`��ax]����j���_}ZR�ݱ�$&n���<@adem.8�c:{i�RwI��+~�� �bc~�N���!���;�	���7�'i�d񱿷J��J��{�>��!�Đ��U� ���^��� qe��D(0���i8���CW��|+>��w2*�i �Q��?���Uϋ�v��t�y��[X2|�ԃgOA�+�Th��o�3.��������Qm�"�jMϫ�K"����̸|�Fp���z���x�k�;Z"+���ݸ:������z#�a��NG�lC��2�����Q\����D�Eˊ���Q�SA��"[
�k���^<7k״v���-�E��|Z��W�V?K���Ȯl~@Z�`�X%n�!�����[ۑ�l�T�9X��;x�E�w��R1Р��Ē���i	�:������4?ogӓ�V���;���dRjB�B�'P�%�VmÙO�$�<�k]+�������0��W��_����֠),R``|uM�FA�=�FQ�ؕ�|���|�q�4�=��FEC������*�\}2��� �eT$��c���>�C@���䆵���m���ǡCl�k'?��.2�n��ʹ@0���q�A�J_�DU*
Sx�0����m��\�亘lZ�Q�:��;�vT!� E����P�����z�a�,��I���AT-��N"�wr�Uᬽ�I�@���4z��q�a�.���F�]ߡ��t�H��7S��7f/Xdp��;�Un��4i��v��O������&?�Gq't'�l���58����n�ֱW��"1��q��G%��LS]<����%Jı�WA�g�T�v4Q�w6K����
*�k�>�\g�C��@_&������v���f��QӖ]��6,��M�W�aS��,����k/B,*� ��I2���j��s��9���k�\7�_�p�Z�[�k4�}տ���"�o�����?���X0�>Te4�1� ���׼W#�b��N�κ��f����zӫS�vөF�G/�Ρ�`���i�?�vx���b��a�͵ʮzÔ�%V�z�_���I�%�6#(�i�4���Y7B���w,����z�*��o��d� 
�:�4}��_�Gf�JrDC��r�4�m-��Ur�����ta����D����s�M3<��nS��m�MW���l���g+Y�(��
���=�J�����[Nr������Ȫ�_3ڤ$1�R#�:�rZ�o�*}2�s�@��]����C_����'Ҫ�Ť;���S�X;���MmK'_�NC�ĵ�����>���~���(��?�����˙ru�i�+"�bШ�SI���20��"J�x������1݀x�k$��I콬-%�L��Ӕ��e@�f�L{K<ŅN�<ۡ]�E=l0�\B �? ����*(��r�d��]����B
%y�2�9����~s��VG3�Gd�@M�@��6�)�]�;��ܜ`EDr�/n�F�E {�u���KAV��.Rr�����@SlQ�J�9��4+�Z��%e���r�=���K��ҝ�m��f�kx���gfFA�[���n(pI�E���P�Ԯ'������cxo�(ŝ��i��/�`H�Q6��9��t��������".�"7����i�j�KLeÄ	���A�ʊ���o�a��t
����ފE'���0�1a�K��*����ꍽb|-K��.��6�ڕ�Ԕ�3P�j.��v՟���g�}�aWi\��$5�[���N�����T�~�?^����C()��u'��Q�^1'&��E��h%$	��W�HҮ�>sVS�G�r!lڞ�Z�H��9P]jiw�?S� ��#D�����hvǫ<�*���&qѧ�@�p��������Q��+]�`�g.�rO�+z�tʖ$�Q?��3��Qc�M�n�*��������7X# �^IQ�Q�lk��I�C� 9�({�w�T4j/f�N�% �}��O;բ�ņ��?��GN;R/�c�s�K]�O6���-eb_���D`TT��#��k�nn��z'A�C�-U���Bg�����O
#6��nv�_R?�b����f^�o�������	~��X998��0���e8]z���N�U����ae�&�n�g�.	� �����5�)�~i�	n(�Y��m����I\�[���� ������(M��]�v�'5�K�Jvf�KH���v�k��p�S�G@�h�s�
��V�X��S�>
B�x�E���c+�����J��&���a��Y&-��6Q�����m<�r�씣��rV�hFŗ^!�*e&.sm]���hL��_}����s�D�Ĵ�P��5J�j��b��QUR��Xkb�D�%��J͠��g��T÷)bD ݲ�$�����i�K�M��?��IĻ-F�/�q`S������e�?O��� �T��h��iI_��!&�2���8�����۲�B\��Ge���P��kQ��u�'�/偟��yS���K���~)1`���e$�s�;���ETs	��#�za���2BR<���i�&��oo'�N�9��+�m ��#��J��e�cav����v����2��z|e9A����]9)�'�`�)�����L�u�e��k����:�I����1��SvQ@�d��s�����+�@C}K�U��}tH���h=��I�˞��3H!<�;��8�%�P`t��h7��=k�<����i�Vgǯ��c2 ��Y�)Lߺ�^&;����˨�!�1����;@�r��Ms�� �����$��ʩ��ڋ��M�X�ݎv$׽
1`��I?kƽôc�H/�*� �R��t�=����7t�(r7]մV5M#��O��,4����N�{�=i*7�C΄�+�DI����E5ʗO��k<�����e�����7��_j��H��ɉI�۱�?�G�M� �6�_�_��P�|�!��C�*�U��۝)�^�fYdBY�e��˴�1Wt
�^������N#��aQg�O���K���@fHOoЃ=C_-s�,�Bv^�����O�T+A�v�/�`SrI�W��0�����,���[I��9Ɋ��6��H�b �d� �t�kϿ-]�
�P����9L��@u`u�'MyĬ�M_�dk8tdY*�8�.�/\P��@�H�o�ERc��Eϥ��g��ے"���tl_�������8��}�y(*U�n���"����V�K���<�X�S��n'��a*�����9�dƟ�<���Su��	h��N�;�d�ۅA'��|���S
o����� �^E��i�5A������5$-5���r�T�t�^�c�ӵ���L�����P�)�g6-��] �K��!SD�Jv�;b��|dZr�l�����EY�Q��n����_��ڌ������Eo�%�����v.��l�ʞ��	�ú�r���.:����8[O�,� J�b݀�V,�<M᛬#�����R�F$� �40ʋ�vD?-ϧ��{��oC���+y���`رbVJ*l+�y�%$G��N��I���e����#`]S	D�9Y�����>��T�ea/�
�����I;���<��7*ߝ��'t�J_�x�k;���s��K
²K���kX�*��	?�q��6֘x�� �o���!��%��
NxS�,"�޴��X�;`J;&V,������Ɣ��k��EX"�ec��I���4S��-��������`C%�t��'U��escb�xc�1h')�pq���"T���0#㋸h@y$z�R���Z-ڥ���R�}�\HX���n�#�l̰^�A#Pgl}��5�sA�ǿ��G��Dy}%�H_0��W3���6��U��-���X�A,��.W����~��S�!�"��afq���\S��)i���c�#�4��;������Jh��QZj}(�������ia�8t�B�;�v�������49%M�T��0���.�5<R�^�ȧ�p����,d�P78�~�X�I�f$�du��S�A�H�A�����wI�]e��a:���g��&��zMG��*�!v��U���6�K-��G)���1oi�m�7�@Ks��@�[zY�!�c�4�Y������e���*��2,,�ñ���|̠
m$븘��NQ�lG?����g\ $���҄a�=q0�#&��j�;� �7�o�L�\���M��E��U"d���V�y���{��Q�i�2DC.Le= �{5#���)	u��d���soZ�[���G��\�p�Q�'H����X��++9�!�T��.��M�K�h16�+�3�]��gQ*�
d{���&����&H�EYi��:�jm�A�9}l'�&�:'�ƻ�?�f�*͒N��xm���;��og�ޝl���wv-ϏG]�����X��Xx��^/�K*X�x	����ʴ��ֲ]]�ͤ͛oe�|">�rh�Ņ0Lm$�1�w�L~g�O3����q`���ն��M�7 ��Ȭ�j-=@���-��ó�M�YW�^0� f�M�"�hy�q�,XT�U^S���[�HE��s�[��]���餗��0� 7��9Q�Q��j'�x������2�Q;=�_���B�C|}��h~@7��Fi,FS�Cljx�Iڹ�	��IO.0$���s�� h#Aw�$Q��l��?��G�YT��h��J�ے$	��a�R���[n&��Ч���s_���P<�������H]���C\"���m�C|s���ê;d�m��@CC�&�XR��M��h�e�G����n���a(�`%��L�� 26�7G������|e�O���,�l�x��ӔT�T	��M��<84��LjqY�r��H��fW���ra�MI�+~�0=�.(�~�A^g�x�;���G��;���`��q(�M�6S�\�}�5�g�C��q|Ϩ%�5���Cv���bQx{66�� g�C(1a��^H�eB6���E�C�(=N�;��.ޟ����S��9O��/���*ٜ2��K�>m����%�M}�|
���wy
M9�ޭ�G�`��jz��"��E�6�n���5��Z�����/<�$��=���n��Q�T��GR�`�?�K��i���;�{��f.k�	�r+�I\tJ�^1� O���;����atql���ٿ��s�#��	���j�q~l$��~E�F��M��Z;g]*<9�֋�%)�:��\�W��������A*����A��@����ێd�@_i�Q�bQ'��G#�&:}��k���Vƍz�p�H_�DMG���QG#@~��/9y׿�h�SmYI��mJ���ϟH�N�,�;�B�y���E="�L����g9����O�ۭW�9_Z,qS�-~q���(b�u4���E��cY�^e�0�7QOU&�E�(�{�z/�.w8��Zd.��J8���绬�B����`ՙTj���N��L%k���=��ĳ�e�:�������ꌘ_��<�.1n��(�����7g�r{͂l$��Y[	�@j9�Y��̓_9��&���#�� �4�h��ۭ֯̕����Һ8�t9�bV��b.�|�b4
l� �~<�Dz��(��l]�q[���y�w�w1h�KJ_�uh+gl����5��޹�KF�3�hb�@���F�&���)yE�3��:p�I⻢��0��Ax)W����R%����"�Y�)L���t�?�j�B����µ���I] 6�٩�'�-�"<�3�`�}��l /hZ��˷�g���v_�uU�)�QT��I��C��t;�%�ϵ{:v�ap�9X�m9!��{�>=�.2-�����^`Q$��\.,�Wh޵���c� B��_g�-�TU;J���8�w�\�(R�,�Z�j�����mU�1�J20fp��^r�}�Dy\3��/3*|�ewy-��5���p.(-�d�W��FՑ0�P�j�+잒6�k�$X�5�����[��Y�����������b��0��7���[�����~�r�/�qӖ��a�-��w9�� ��8��h~Ě=�Dv�L�U�ԗ����o������#�����H���%��h����#k��v��.s�S;N�R�E��Iy~?�^n�������N@N�p���v�+�H����G�@��	��1�D'	�m�t�;�l�p�vs
���AU���'�_�Zo����g�-��+��/X��V�<z0��9���2�;�g՝��b^�Q��.��{ds�����?܄�,ls<i�ǁoҜ�z��9Tˌ)!b,��^�M����l�OB��[��>ظKhtsW Gq�)VP��#Xvu26�JW��|�$$�õ	.���Љ$kV^�`VR���Ӄ�}�T����$\�������J��rda���Og��u	ȓ�,�s��z�|t�e*MBL�֋["j)��nPջ��a�����J�"dm��[�Mi\�d�V�����]N^F�ޚ�G�@Z)�{*�����M"�����\��"�{�8%-������H����I/g����R��x��p.�R�;��C#�%��ĥO<+��#�u�{D�}y�.,'ճ�{��W���I�?���A�C'����|��Ms�E���?%эC���ꆩ�2*:$���.]mp=�F��?x�l��GI�o���&�$�y=,�����[�#�6zOC���_��1�X� F5Ȕ��H{���G6����V�2V�2�cu�~���>��X�bj�� N��v� �Ɇ�Ʋ4Г{����6̇F�����O�a���p�e�
'���g/W��3v���	�;Tr� ��������D��_��;H����V"c�2PkIO��<^{�ٮ,�vTI�Y�g^�J=�X���Ʊ��9�E�&��HW	���+�`�B���[G� �Y��"�s�^ԂL}b��u��w$6U��kbڞ�-΁����c�4�FD(�q>�,�M�e谩���R�!��u�˃�넣-�Km_\ll�VO��y]b�!����^�H��(��%7���G$j�(�$��4��x�<�C�\��1g�葆��F��P� w�Q@%U"��{��d��g�uj��@����h�3����h��2+[��*m�H(�w��]�"��P�a���O?�[�-�v;4w?��t1	�p&���CBO�&������먕T岏��ĶI]z���B��F��9����x�-�d��gU�.j�{�t�d��0qǫ��C���f�I`́Bp�ę�ro����]$(�v������l��8�O����_ԯ�9�t�r�i�y��$N+�S&�K�mR7�K���t������A���Gj$o(�eZ��8]�Y�{�Wx[��Sԟ��j0��I�@�*���Y��AZ�A��.?��O��Ľ����O�zhsWt���H`�[��Q�/�� LA����&ݢ9H��j�6'�b����FZ��e�D�/I4��Hb-���V�Mk�g}�}�f��X�w4,�s�$<�K,��	��x�׀��=��Χ����H"�����yH��%�<h۾*����{����b`��ظ(�{�t��W�'��y���$F(�kG�u��x�d��� �]՜�KclB��� tN�*����R �dNE0ѩiߘ��f+�{ͬ��G�����֙,��ݐ��B��G�Q��@+���Ə�ǯ��8�9�}�b7�+BM��
���nf�3W[��$;י˵+U�(o��U�/g�ݓNq�4
{�Zi�����t��kj���!��5'o�~��G8����X2����tLt2�ӱ��lޙ��僤:=�灙�~�a�-��@712Х
��_1u1���Pmzc���{ud=߄t�s�����d�/�-w�g	vu�^%�}=x�P���e2l���[�aȴd�8*a�r��?�$fM���D+�A��Y��ڥ�6�rj{�g�>�I���q�cW%צ{<>���Zz�G������$Q�"���o@ӏ`tO3�q03"�g���U�\qLWP-ߴ�Z�S�{��ym/�V2�a�W��6.̵,����J)
31��peO�;q ���|�N��p�����W9o�3nZV�6Xr�yW/�p/k��?}���?Y<<��J���#0+�!�s#`f�S�hT��'��Ϡ.g�R��d���W?0��hVV��7 U�y'1�hۆ��n�&������i���c�j�w�Z��ˆJ��٠�Z	<�;G�l�����8�[g��q��fxC�!�e����S��u�9�\��^���~��>�Q�4ǭl���CT�����~���o�_4��O��!λ�#ӭ�|i-w�ۭ�B][�2vc�b�Z��U	�?�ܻ,�2)��ZM-<r��4 ����2�A�����dw0�M�������-	�[�3|Y={s��W�+^��*�0��!K�����ś���pu�.��)(~m�}��<��t�V3)�o���I�T�(��Y-{�eg3��<ˤW�!���h�  ���I��DK#��i�"�Lo ��	K�6�t�	�r�/����LX��Sl٬�����9��ŀ�v
���L��}��t�	SQ���v��s)�/: �/Ue�Էʗ7�l,�?�6��y�%�lҒ��t�ԆA�v�9��M���II�L�r��{i��?ቆ�"����yGr�V19(��<Ny���rrR̴K�Fne�����Mc("o�	�m�s�h�$$\#`�(��
�W�����6z�у�t��O�6���]'ֻyӺ{��nV����?�R>A��~{_Fcd���V^�e'� R�!�/�xo�Hg��\;�!���j�4��@��^�L/:�ˡ��,ݎF�[n�F�8����3��K{7� Ȏl�'�%D�g��|2s���Qg��}�3_��]m����>\��iLk�G�[to��NR4)�ޟ�)��䨿4#ۀ"�:���s,����j���|@�M�x��^sZ�a_��4�rh����QV9��WIIUWKB����$d��KO0�'���ֳ�5�z>�hr�P�#�vx�9V5F�]����T~epx����}��/� ����qL��z:�#'�b���~��=�z���D%:^+U�z�&@K;X��yv�n�R��ӌ ���)/�đ%�չ1�ʰ����\�-{��%�������V�*0Η�\�\��fA;���с�C�#8����i�t<Q����1Y�~� ��K���b�Uwzs$I�M�����)�'Z"Z��s�ȻZ�`�� \X�9��e�z��_Ij�m�T�b҉dj(w	�~K��IM;�Vg_g�E��/K�f�}�8���D�G%��7�9W��d������'K)�a���23��*������{��ރH�,�V���^H�K�~X��xTq�a����^N���?�����g?AF�J�2���!t[��,.	�댨1πc�!����d���H�)m$�Ə�#� G��s��Ń� ��b+u�&l�|3�5p�B)�J���n~ZX8)oհ���w	k4x&����xc�Ǯ���ʸ�E���2��훐&�@HQ�����*�.C��+�U�~ͤ��Zr�JB�]�xCoܬd� �P^�òQE���9?$r Dcـr�����Z���Y9�~�p�e���ֻȮ̝j�PC����=ቝ'3qoC㌍x�@��ػ��KU߭͗���9�W����f����DYfw��x����#�=��y�y7;$j�$���6i%Ys�k���/��{�h�)7��������kT����޺c�?/�*U*W�s���l�}S5�A*��F����P�X�Cpk xq���SL��1��J�G���d/_;ᄤ��r�G��o*�#5�S�E�?|>��_�E���I�[��@k�?���6�
=ޛέ�v�ԃe$Mo�C����a�p�J��Ŋ"�dy(��.��Ƹjl�����Q���T�>7Y#�^]������<�$4����gV���r���a�1�>��T��*���@��Ⱦ]�T�������fz J�|�7�g>]s�^o�R�4�)��{�b�aL �˳zNPsf�!jf�E=�~���ʌӌ��jӎ���X&������B�*5F]y832q����=u�2��6q�r�����VY�I�,��bv���s��{	��Ლl��M[�͹r��Y���i�JZ�
 <m�j%2�:U�x��lT5ls�����ؽ7���5�)'��G�����x)n�Mx�	~��9">�NF̾�A��8�,FL���'<�CO �k��՟:���R_)�$���A�/����/������p��Hp��e0&���_`� 5y�d���N����;������_%GaK��gE>ei� �H��x���	I�\Md
�Y�A�rOS	��]L�R0S�%lѠ�'Mfaꦖ�nپ�}��p|n�!f"\����(�k�t�_������`�K�Sj�6�FO�|{9��"��7�{��<�k����- 7��S���}MFO��f�`��Kd���}+Yyg������@��Drҏm%�Ŋ�`��{㱕����[�wI�l�@j�6a�sh�ʽ����'��v�)7{Dj*;�@��̖W>�4���y
 ���6r���Ec3�/GH�&���ڐ����\��T!���_������H�}�����@`w&$����5�����_�	���;�.���ɪ
X��C��Y_�ɀ^1��^ơ�����#KGtԄ��k�+_���!�t�"6�`����;鐱�g2��]�����LW�v�&e�,�O����.²>o3�.��^���V{����cD�b�*j�?��/��RRa��Gb�$C,w���+�b���>���34X5|���	B�,�mF�2�44�|�k,�o�(,���A�vmB#�L��N��;#�D.q��m�;<XitbpY���Wkw�w�\�^-���-��C��{J�g�[��ٸ�Q~R��LZ�Y�|�&�3<Y��~4��S�"-c��:h;�e��y؇l���f'c�z7���cvZA��}E �E؄ˍ�Q3.��i5��(�4���䪥��Z����)���ن)�,D��{��ɱ�3����J±���9�'4Ma�"H�C^�ڣ�����.���T�ו�f��p"��"ѨcV���M�"�C���=���ZH����ih����^�/@�:��	P�G2w�!~zµ�7rg��"�.ͅ>��'0�=p�8Z*�P��C7(����i� �2���`[�[|/i$��:��w^"�e�hx�E�
�,��_%��j$Κ�-�g���Q���Dh]�u,4,��LNv.�n��\M;��%A���
���7��Xx6e�\%k>��>2��LL�(*�qg�k�4Z���c�0�i�#��;r�s���T���  7�)c�r
F>[_���3�Kx^Z�t5`��9����X7�L��2�Qn⼘7�Lh�3�� �,5�0���I;��7�ڌzt�k3�� �=��o;�ԧ֌����✗{�����l�i�;�!�P��ı�����0MX�\�;����k�20mP�Շc8z~/~����bbAS[�(�ɸ@�^���v#&�	ԉ�u%�N@���
R/����������nb=jz�1�Kћ��&�'�9�<K`�B��Q:�Ro� �.�Y"���~�(�2�hm�m��i��mc�6x�f�` �9Ա�?��n)��^�����yR���m���+�[l��M��Z�˃��&T/Gz��04+�@��-����>�z�[S�m���l���m���\4�|T L�M25E�]��W�x�f���03I��x1�]����k��v��W��t[��75�v�Õ�̀T�O�`�ܾc��e�r��ٰk�ߋĔy�.��o��µ	�R"S(Qf?�A�� 8?r6�p�-�>=�4�q&��Ƙ;R5/)��R�2�J�]yJ��2�������/�D���w`�e߉�d���v>��dվMc��g��"���]��
7aʫ�`i����7-D�Xd�xz�����#�hr�:	/K���������?: �(Nu6�O���D4\��(B�ͧD�w�F� ��r��^�/y�D�@�!J�t_$Q|�h�+�}oX���ٖç�\[��8����m5!��"`�����Qk)U��D��i$��)��`-�Im���i;^�� 9#�W&#U`�1�t��HU�+ʄ���o:s�#w�Vզ���ˇ�ڐ(�0�����t��bK� ���U�����Q�]'Y��k<5���M����5�>z7�O'+Ʈ_��nq�K�w.r��)���9"�5\)�����7S5My_A.a��{��Մ���z��?�՗B��<�p�S��`�5�j�r�T���Rb�;9$	�1��s��Ѭ1�7NLչ��hZ��� �����*_U�@�?8zG!V��������J�b���Z�3f��{���3��Z\���6c�x㣝��w[��X��u�R����m�2�,7*0P�����eVX.2}�
�'�9�<����3�w
�����O�:�i'��(�bH��8�VV�/{��蘒z]�j�/��_,*.a���� B�Ť��՝��.G��Q�E�]dV#r�R��y �FM�E57Y��B���2�9������.�����:�����$HÏ�c8�F.!(�N��ʵ��.ɫ^�a�X�N�IR�]��e=!!L%���ga�>cp��'c�/=_���Х���n&|,��k1�� C����K6x�ND1���)�ԥx�јdw�S	,�2��7���r�ի��[
��}�R�CT��m�|�GK�����0�[��G�%��6�~��,��,6��;A=.�>���$�����l�;+� h��3e����	������٘��9��h�bp�����j�rfΆKv/���H�� ��#YKb��f�(0cſ`i#�4&�co�S�wܩ�(|`�@����a��J~y��������b�;����6�U"M`?��>��2�<[;������te��%Aw�����~�i��ˬĴw�G�k�r0�.
�"ӷ�i��jmU��Sd�l��p��cչ��c�Z����13�E�W��k�ñǡ]��=�U�%r���{�4b# մ�{ah$ҋ0�UPX�6�-��CU�i�Ts�f��è���}\�<0�}m�="���(o�|>u���4mI�*��r�$&�J�I�^� 9F�~5��^G���G\ҍ�ǣp1t�� �ܷ�3�~��v�T���<Wc%��KM�B=[)y�u@�hʹ�	��^Ý�쩥�tgG��.�}<������{ǔ��D#��8G<n�o@.��$W9�A0V���<�4��d�(&?L���.{-��	#eJ�}E���2Q�޳�����Pm�:����a�.)-�	�u%yf����ƞW��2)���Cq�ӯ{��ڣ�w��9�t��F=���y��k lú���`wk�px
��5)oR��Bc	��$/�K�#�!ǫ>(��N9_���ŕ�'�8����\��'�ʷlO٢z^��yH�{xS�FO��
1h��Ʃ�r��-�?Y�h�eݞ	�V�#mT�d�{��o���q�D�5��bl�5�/���9���>�Ѳ<pi®������Ü8�Q)@���إBK8\|�8���"�tA��[��O�����yu���G�+~����p���b�Oi�/��]�1G��v$�r��L�X����Xs�T���@�9S^i���9�Y)�q)2� 4h�ж��ǲ.�Q 4n%t6C�G��X�?b�x�]����[^�r�]ݚ�0P�|\�H�p:�Ұ����г�'+�O�|�P:y��@�M�@BE��k�f]V���F��Bm��d�"J���C�1E�Ug@ԧ�4�Mڡ��x�e�������b�#�i�f�.D�`�M�ff���tf���S�$f1,�m�e�ݒ��(��.��J���=����N;�+A% ��"Ԛ�������mR�ŧګ��	���u|�5=%/�Ձ���h��hZX#B�^gq=���Ja{e�=*�P�f���ma�p�WZ�M-e�g�z!rב/����Lo��k��Ȭ�Y�����gOǶ�(#^�$�P�7P2�@�D�O�?����&����D�y%��|��n���<(p�σ�r|n��ڒ���WNYs��F�CD�9k��l�*΋Pܚס���Ǐ�9塑�NYJ���x����a�Ҋ>����:t�\?��-�٦s]�I9F��C	l��a����,+��7��gFH�z ^\�@ʌ�N�4��wY�'�K�ݱD��:K@J�|�Z��'%QD��h���<��m<m��ߣ��T���7)���sK3���dR�R�gR��z<kQ�{�7�ޮ`FP>���P���?F��`�؄� on�OW��{~i���? NͲz�+��q��L�����D����k���ھ�A���1j�3X�]7���	7��ժ����`��obF,��}r�����=�B�[��n:��#A��o �E2b���T'J�]�Z����y�/��$��d�I�5����?�r�k�2�]f����}���4�����R�бD�������t!?�m2��?'��Ĩ�r��?��t`��AJ���m�d�a���@�.v)�� K���âf�//�n����Ul��z:Q��n�7�T������+�X����M�?]�u`~���o�gca;��,=�����In�r�m�ܤ�[𪜉0�s�#��k�����9W���Mo�#A_B��v|^����ȍF\���"՚;�x��=&��Q��$�{��"NzrTI!�Ş�iK�?��u��ġ�^V�@.�-�����K �9�s%&�w��P��ߕ�[�/�y�S�@Z�������s�"��f���(�&�� ����nΞ�-o���#�{qH�7�n��s��ː�\�S��)�W��)(%Ȼ3�S#�.���kV�3eǨ���-p�����p�!P=�����~���]��:�8�^W�,C�D|�DZ�أ��~u�"y�^a��7�p;�;��.�~��� yB�|���y���/�Fm����%[��]�1Q�V��#�\Q��=N�J[���I�h��V�ќ�@{[�sJ���-穇���i���F�����5S���>��� ]*�Q.�pq�I&Abg[~�	%���t�Mq��d(�Dm#[ԝ�Š�p*�"��^7tXE�O\�ſV��)H�W1��g8u���7A0y��(���x�̬GJC�����샼
#o�|g�?�F:crO�
s�����$�j��#�q��uR�A��B�����ѭ���zxar���XR�}ϖ@f��(5�4
1�I֏�i2cA�st�3ر[0�a�/����`L���X�Y����Pm� �z�!wK���-��\6 &+o֫?t�F�xq�o���re��f�F9|�S��?)��;$��l�ל8ٜ$�����>�y�^�B�xk��o\��X=�ڌT�]@[[0%\��Ǿ�5�y����[�����5����c(QD��R��R����"j�n���~����Ì�r�{����*�T���9�N���鍨W�(HS9=h��@߷���2 D�B@��8h�?0�e���jv��E���!��]�(Z����x��'�`�l�&,8R��q�:���nD�d�Di���t�gpU� �G�輗t�doiJ�O��]�O���v��3	��ws+���Jq{�,����!�XHJb��(^m��ޱ-̥�B�TF\IqA[��u-��$�C�����A�W�Y�iP!��l�x<;X�2Ԍ*J{C�<%��Ƈ���aDJ6ѡ����뷖|pXŢdW)��x��.��}�;m�4`����>��&	��6y�Q[���dH���6Uňr���Y>^|��ҥ��#d�c"/ܓ����+^4�%�и�7��BԽsxXf�W��9↵t��;�����$�+���U�Մ���~=f��I7��a"uXN#K�K�]c��V�1h/��?0"��VmQ�`$0��N�0�v�"]�?��k�C�W�]}��A�(*����G�dk8w�+���X\�?�n?=hD�Y�&G�,��/�v���SQ| 
m#9��:�B�C��L���`բ3��.����E�w���M%�:h������?����c�9��K����YV�R8������usWU�<<¶����5p
��MQx��zW�W�$�Dj��J�w�!6e�����kXVE5;��@����c��V��/�\�=���+F1�9��TB��>L��@��^d�A��{���__��g��E��z],��޴Vy�������&�]�>I��c�D^ʻ
�1�_s#B��X�阨~�<wX�r�Q�S�O��Ȗ����3*�����[�f&��m�r�ظjp�
|��y�ǜ�ͪ��{�r���f Gp�Wi������a�e\���4��-_��!��2��yU�wx���.O6�,:��ʉ���ȹ5�
gJ}Y�r����bl�\F8Q%�-7xx�g�+�nx�5D�WB��"����W�Ӏ���v�]�d�X����'�J_�T����\u=���U�TM��b.C� �F�!.�w�>Q�,��M�a�/�Gʬ~j@��+,��v) TQ����Aw��l���-� 'ik`��My�&��k9�Q&a%�W@��=����B��w�z6Z��I�F�M�݅�#Q�Ȱn^�ջ�\ȭ+:(��_פ�a��� ��W��4�Hrڼ9���H60�Bt-��q�9;"�	Ak��t�zK��2u-��#�Z�������ӫΥv�K��1l���#Bh軭E(g�8�^�#5�k�#�~���wu!����ĵO���b��!� ���E��}(;����V	٨L]�q�t�'\l��ɿ��˱҂|M��2���g�F�N�otR�?�o?z�/��?�~��2�c�'U�b�Ɨb��F�a	b��5�9��s/rуIO��k��8!�~�&v.�^6  oP��K����[8$�J�0S�V���9��u ����{;�7SZ���a����:T�IM@2h�`��n��L��L�Q4U���Q�ot��� s���Ę�yN�D�ĠL}�
@8�]+`�HkTg�0���7��Z�{c;���c����,&K�t�Q��9��K�±s�0��k���p`�;Sf�a������TL�}*��I%��(���f��
�ǵ��XrK3+8��Ř@��Jw�>�\-R���I5�ǖ��C�R�咥O�X�mf:���Դ~��e�p�F?*�H����nm�l�U�g�X�+�� �Sbcە���$���h��i�5������co�uy
s ��C�����ָU0�|xx���5+C+3�����V�D��8򐏗)U� �:�M��O$�z~p�Stgs��~=�K՚��v]ژ�]��{����z�a����Bz��w�+�TP��lx��bOhɟ.����͍�Bc ��%͡����L�ط�-�x�|A�%~�@�&0"Y8����z�DpW�즐*��J�N��$����Ƿ&�w'$�W������>���T�h�0THN�Pw����EĆ��[\fA��^*�i����e��Hș5��ˢ����v#O��2�X!~Vcc�A����i� B���c�b8��ey��r����,7|��70����C���dMM.{FO4��"��];޵/��&A�)R�A T�.���G��ۯQ��#��^��.��o$r�� ���zC٫�?��=��3
zC�8¹�lhi�U�iݠ�,+e9�i}���A圏{kY� �a��XI�P�BbQ��G�M��V�O��^�����X�$��USD�C�����rnc�^Cn��9v�BoxǼ���ys�O����x�/Zp��M��	����R��^dޔ/����9ܢ[G�؇�S��C`xE"*S�EI�V�_���L��ۙ��L��ECz�`�p�1�����IᏒ�0�l��6s�l7*�)���c��*:#��Cqpg����S�o�Tѧ�����9K �]�]O�d'�t�3�"ST�ܶD� ���-�đ	��~�b[޴ְM:v��:}�e&��KN,$�̫}�g��ٮ�l	v��kLP�`�����	��mu&�ֹ�n�(�M?�7�(0V�I��]�,���	\[c��ctl�Rp�+��)�t��}�G ��@�_�t��^�r�ʸ��I��=GIp��m�Z;�v���_Ò��)1S�DD��z��z�B_�[��<J�&��2<��ʙ:�AU���x����5�6J�= �������g�/H ('W\�ȁ�w�	"��p�k�#U��cC�A7�ɠK�E��D�L�5��I�$y�D\cЭ����o\�͙z��d���Kµ�1�����(� ��sR���!�mc8Y�too*j
s��
��ZN������hM,��\ ��UR�f�4�;�9N%\�� ���yM�<5�Ts�7���S��} �b�8��<?�6Z	�L����/�\�����]o?�������q-b��8���vr��]i+�x�a-���?��T�P�C����}�Y�
�}�De�]�)VΡ��	bG��u� r������:���-h��qZ9=੊�����[��ow����L$0���q��&V����P��]b�؞���.7=P���{ud��qq��W(�Z5��J]��-zT>gg���m�r���1!W�vY(/D��w��&�֪�X��g�q�K?/Дb���2��&���?�'5R�;s���K��;�2�]����Ph�C�������!��8�p�S2�c��5��RY�2�ʒ/8-�Nu�i-�ϋ�(���N_�';?�\ן����q����>p~�U����Ӄ���Cj���6Qj �� �����]�s$qw�1����z�{"���˼��^t�dt.�=��L Uǆ��x�Ƭ�8���y�4[=a�aΩU��@&}	��4�\������T��
&[�uM�q��V�g�8A䤆���H$���U	8��:*����Y>��=�ax���u3竞Hp�:@�!^�-��e�8�� p�,)t�=K�V�F�"��x���Lp� �DFj&/|�m���RsV��� ��HZk��2)?Ȕ�vG���+��+/�X">�D QY}r�e���\?Ji��.B���x|�j�+��j-��U�]�Lk�(����v�cb��+���Qp \a��-u��P?��X(��Zy�.N����@��$;I��%[N}KP��̉�.a��r���"��ޖo�}�+��`�������`Ɩ�T�q:i�y����sh�Ͽ�@���U��p�J-�!|;!|&�O��.'|��!������Ƽ�~ǽ6*�	
1��=!��8������WIpD� ����ݯ7����3�"���gf5qэ�=�<�q���^@+n�:�
��dcC}~�i��% �&IڕP��'��fs�%��cti�zHְ!�P��x���B�7m�VP�m-M}(�
]do���9�kH�3��n�,��Eu�-#�� @)Mu�P����iva0�8�(���Ѓ�gQ&�UH'j-a��l+��kY���
8S;2z��ҍ���]oy�Y���u�%�������0�X����3*ԟQ�,�u�`�ȃ���W������Ҏ���&�]�6�9pKi1��u�;Y�7�9g`f�^8���H����w�j��HCp�<��B����Df���&�� �V�ֻ8t��"��ʄ؄n�c��Æ�p�<v�8�0�1V�X�y�I[��v(#��fʈ�?�p�z�J�k�Ec�����V٬���m�5h���xt�����Lϊ���nh�F��Ve�x1߈��nR�d����x`��衳�<��ߨ��������`G!���V�L ��2F��_����߲��R�Ę0c5tkU �  !�G�A�AY'��A�U�Ø< 眅[��!m����Z�q~�?Jh5P|���lC_v�Y�01?����o���EV(I�>��ӻ^������LUF�$ s�wWl�K!�2R�u���ԕk��}�d>���M�k;~Ab(��r,xe�VP���Y��S�o��N�c�{@p�ׂ����̎�2����*0����e��*�)���Jy��ea�rv�a�_ȹ�bU#�8����|�K�M�.�ۢ|�w����p���H�A)��Ia:���=굽Xj��[�K�����E��ɌIG夅�x��$}�*ſ�x����d�p��2謔F���$���*Q�ur���X�N(�.q��nE��gwiR�Q��H��'��W��e�qbـ%h$�dF0ր��b���N<�n��Sa0�ݬ��tخvO�1��L�2��,�I�B��ӆ-�7�L���3�n:�x"��d�QR�x�}Y�QN '��^ ͇�KN�qۻ��Ab�H2h. ��u��Y_�$���]D�9Tcv�w���ndb�PU~W�T�'���4�E�����l�6oi�CZ��(�[��K�`K����P'�tt�͸?X`"^t���h]�Ft�WOv��0"���Gw���j�s��4�m<��w����rt�n0CE����D2�&�@J�Y~b�t鈂A���_۔���6 �n�w��!�T8枞G���Yپ�Gcwf�P�C$3N���h�P��ij(��4�i14d�Hѱ�#�����'�.=�=^�v1��r��9]te� �������mC��Cn�j5َ�8Z)MD}�o�b_k*�1��IҠ;H�?�M�|Q�r�ǛԶ�=7]��Ư��C�/�U�����E�/nb���x�۵�+����y�8N��m���)�N�`�6|o�]�DELmD���4d{��ހ�O��:#�SV�+kD�H�U��Q7ɰ2�Z�t>7Vwb���[5� >
�u:c�ݦt	�@�5@ކ��%'���C���%K*��l�}a.Ft�C-�%�zK�,�-yq�F�'__������j jG���[����f�c�$��ؽn ��:�!����0"�:��q�n_k,W�6������s���O�5c�iR��MH8]6B����'s�`%*���,����q�J3�Cڭd�j���^@9���Ƈ�l=�\G���a�VK.�g���wf�!N��./���,�[�P9a�Ql	d�$��
�y�s��!�O��	{�Q���;g8HpN
?e�*�q$@�*��<�#9���y=��ӣ,��h;䋾���X��'z{/��g�.U�H�t�G�67g���Ƹ�7����P�!�* �+:xƽ��.g%]؞��F}eSFP�L�o����u[��2�\�zs�i�6*N���<z��f����j=�`d�d�����|�y&oZ2����K��Ռ�?d�5,��Amk�'�M�{����G ��}\U���><��#��?F��Mhr=��9A��h��\	@s>.\A��d�OQ�u�dI0!T䁅����'T	W`�gF��( ��P�~V��iP������ޫG�y֍�>6��'�wO8�>����c�"C���cÃ�'����N7� |�W������ޭpёs�['H�p.��:��{w_����~�-�[���҈������1s't��̗o�܄	�sLWܦ��
��R˹e�32�6���[~�|�V;��j�{�x��r�x5L���1��$c̾��U�$ݓ�3��C:8t��>��iba6�%�
�T��{��A�ѓ���6�IF�'����h�r�zlc�3��f c����z��y����S��߼k\i����~F���Nw��x�mj�H!�a�G�nÒ9�pt�?	�\�hG���-�?�o��|֩,��O��.���9��Tb��E _�T�" ����65y�k(s�=8�@ƻ�y����o&DS������e� Fd}��Q��|a-��"�&S�ߏš�ӎ�#�--]�8����c��Jܥd(���\#�m��Rg���W4�*�\`�����Be[C�y�J*�l��g�K�x
���ns~a�L0���h���t�*t��x�6"�1�,'#��ҽb���g���+�]���k{M[��3��n��s��#ۥo�e�ֿ��f�`˂�L�ը]���W2��N^F���}U�دU��
!zDsS�*��U�?�@0���� �Ug����1u�����]3_�ر�80����V�y��`��좹��ک���#����Y��c��%{��O��g��ђx�
���(� �.d��1�����}���aJdY�J���!�)F"�|N�S9�����"�� 	J-�j�ZA��~�Lf����O����܀���y�*���ߜyV#��O:�_%�h�d��	֘�v��8�2@��}ź��d�wD'w%�ܪP��kq:w����&��&0�����',� ��_��^�_cL�V��)9؃M_����;����C-^R`�dd���O�)2�2��
M,:��pA,�,k�5�΁\ s���U�&��'!��5�1��yU���� D�~ɡ%uU���bH�6�'��$Z�}g�v,��G���f|��pm����h�=O,�s'�R������އ�ꖈ}Y�[#��J��݇�O ݔ5,���4�^���4���nz��7 /��'��H�o�3l�C��"�%��O�Ē��n�_�Z_bw=�6���`w���23�cE5��V/�>��P�3�~�woǦ�k��&�zr=qk�Y��[��2���e�k\G՘򐨟0�6M�36�������N��J%8�(3b�=|=U@c�
��r�����Q��ԣ�.)�?�N+��K� aMk����1��Zv��q�Z'����Vt#���*Ǘ���$%wɾ���O����xʱZ�Шw֪t�RAV*�ٔ=릧������pi��a[w�t�{���2wp�^�V�k�
��b�?�39�d
��-q��3u�;3X�T�*��L���|>�Ǳ� �ExJVkR��o�@ɲ^#3���1��U��}s����"���Q�tF��,�6��?Uj�@���B�{?�Y�?�[� ��娼}�2gTԖ�eE���#n�jo,y���<g��:.b	S+��U̙�V��B�Rv���P��)sa�Ԏ��u�}p�%
�, JU��gL�&`ij��a�ǝ�9�7A
mݜ���$����:�L9���hJ3O0*���`���"'8�clD�*��S�;	I&}c�.������sb˞��6����٘q;�fG�st]ԑ���޸���F�����MX���t���ۢv��?��%zr��Y��EU`�3(<Q�~�T6t�4�5��zy���YE ]�ز����	�Ǧ�^�U�Z��Y��I�O9*�κf{�(Nɩr��?a��G���N?G����pՄ�e��t��>�˴2��BǾˊ�r���M�˦���d�D?�SdUtC:�a�����[�E��Zng�U���Bt�Uj:C�ﹹLS�'P6��ZR�k��罧��LyK���%����ŔӢ����ɣ�t<9�;Q(�D�_G��Q�7P#S竝`�u5X���ziO�#�J��7�}�!�M>���������e"�co^'vt�Nf -+dd,b����ÝbСp��b�h/*�^���<�Sܱ�Y�K!;��1�2�`���5&�E���"�q)�o�Uʿ\2Mm���1A��Z�{v�r5�KC�o(�Aw��(
�D� �P
�HYU�v�+"Ϲ��,�D��'Q�AO�b��nTO���L.=��ٖ6���6�
�*�o�ܯ�V��@hl������4q!wܶ=���[-�f�����J�0{WY �<��|$�������eH�A5�l�����kک�j�>��U�S�&�%A��h���h���z7ؒ��KʫIa$����X���b�(��C��k�|��ǘ__���B�7��b�D;��z�`ģ�G�'�&�����qRP������ht��s0X�LR��I�	����UBD��*��IA.Xn鮹(ٶNKU�w��Zo��] �?�q[�K��S�Pod�Ht+au�����+�U�r(q%�����ν�z���%:������6����(��}����<�#�,�R(�}��%hf����%�}�8�����B$��
���AW�P���Ա4_�n�E�����Rխ�͍��_��(�qFr�OM�@���Jh(�:(	�O�L�N��b�!/��=��@-҈k'���e�\���(��=������v���5����T@QO7ۘK���)�����Ǧ��}�ہ(2$����|�	��ɚ���G��	��u%���%~qS�x����x'�����z�z0�v�R���hGb�0R��K�V��1��T��Jh��xo����$��ɬ�Y�'H���&�?RX@��7s�@Rx������������������5Y_�{��b�7��a��9ɼ�d���8b�}T�lL��! ����x�芵
�%�a��6�#G��^��媱/\������)j�~�Mh�pn(	���r�:q����Jȡ���w��V>���hP3ߕF��2���!L:(��oQ�|��G�#���ҡp� ��N��p���M���XQ�;ʷٓ, �]u��u�a����J^d羁�hR
9��ܦ�Q^ZE�^����F
7�t,�P�k�t2l��C01�G��>Ԅ|n���3�P�d���U����C�#"xKEӆ�� �`+P9�r� �ڒ!葸�l�(�n��@Q�BW����!�1^��Dܰ�����/�:�U��p=�P�`��RGi����č^TW���%���D @���U�{vd�O{��L�u-���OJ��)V�=_���F>y0I�T��Mp�B��8@�>Q�ꈟ��w��p�z�4{��n 駵��F2���U(W���xE� �|I0 "Z:�{;�E�Ұv���ྐྵ�����������6�� 6���(�������+�-I7刊��z�����Y�n�P3Uvq:�Ug��6���,.�2&@M��+xƽ���&�PL'�Fu�dR���L��A�b��Ւ�h�����Q����?��JW��C>��T���/�lJ��{�-#/Ly"��kԅpZ T(`s�v��M��P)K�!�'�Z��\���/q��pɘKQ9�4`��h�'���g8�A�����ۓ��x7o���臬���&du���Xo,�9Ѷ*���_�GK�K+��w.<�C)F��6oG��v�Nt� ��̃/�����0O�5�ڪx��GL�2O�����U�&��W��f8�r��x�c�E����Z�>�Z�!:�C��NZ�ې��1�_P|����79Ttτ��J��?���t
���WU������]&����{1��e&�R���"�l[�8�:��k��ʪ�]����lDղKa�t��-�1R��S�ü���:�c��[pc�|�ƃv��aE�5M�6Z98��NMj�G��L{��;�dB��R���E�n���{��?��VЖ�.��U����bgR�q���ł��dx:=
3
���O��q�q�S\�KR�y/e+z:d�5N�$I�\i�����D�b�	��캦sx�Nc�F=���]INgjEcA|��X�.�xpML��%i,�2�]��1�s���a{�̎�Ԛ�/GL8�0ɚ�$��4�Y���������U�NL�W��N~A8�fAoJ�E� 5涉�2���I��6��̎ʑIj�)]C��|8�WׁIdc��b������g����ޘ;K����ˑ���yBם�3��R"�U3{�վ#��kPdb4�8zc�d��	��-><9�����l��S T0 v.r�R�l��=�B��UO�,�?�i�	~)�.�g*G��/[��1��t�o��i�T'��@<��G�Q�R��7	�I�&$G�ĪrIx=W&�0˼��ě���Y����TD&TY~	��<��x����2��*���V%A���j���QE+-��hx RԢ�7N���s�4��ά����‒��m�����΄��*�>�m���}�S
=V<���Z���=���L�XmȺ\�
U����&�����r�#֌�(�k��.���W&r��E�,#_(F�u�	Jyr	��Q円�c�w�Avա&8g4��E��<��9�uF3�k`��v�5����L<�Sv6JrT�o	���Hf�)��>�:�h_�����^sk�Z ���;���l'�M���RǇVrj���Z|z_^0��i;=�+��PԈ6�3>�vpG��ff�K�yPK���&tE��НU�ٝV��7i��-@l#�'����p�ci)'�}�$���1�YV���'�%�X��T[`ݼ�7s��v�*���͆�瘱[��{��"CTJ3�	~v+Fk���{8��s#�h�ٝQf���Y-��c�^�6ݍ!�mJ/T�e�q�N��dcj!>E� վ�\�do��P�V��9�D�<�n��k$>�	;�.�*���Y��������`�N7���p-;���"�-GƎ��b��K��6�u��uk=;�Ѹ--��B��2�Ǉ��d�FqpW /9��h�P�(M��ꦢ�� q֧ؓ�O��l��um�9��m,Q�4,�����3�X��o
 h�(�'�U�J~��Փ厸7�C{*�^[+�Fc���
�T�5K'��rh��]E�%��Mj��[�V���Y��Kěk.��`��1̳Qը�J{��X��DI"8'�2�:܍3���i� #��'Ƽ��L�,�Ph��de��ȃf���!p��wo����1u��6�D�
Y�w�$1�O�r5%S��������M�Bz@2�= *ŷ�Įgj�%n)����ߴ��U>��i�>��P�ݼ���,b�1.��2���� ߿�@X�b(I:+ƙ���
Pk9kæ��e�u��l��BdT�[�.��KH�cښG?w��M7�^@	&=(��'�(G�Ֆ�3� ��*!��[�ƅ:Ԃ�)d?]���`����x�X�d�5��nlV��;���i}�y���7T�WH��^&��UXO�I�wF�����{����ep>�=�X|�� (�j��_`F(~ĽM����3>hQ�W�ֹ"ż;m�RE�H ��q�gy���9#�jP�^���_\>�~�	���6@�OP�Ea��(q%�Ϡ��̞�2��8������ �6+Yd𝭠�*���8_pd��=g�Q�y����m%)��~nt�^�����940�4~�އ�˽M:�? �m��r9�U�:�!�HYfn`ݞ��k���^(�`����0���[�CtX���eC��Ld�:@�������	�:�����R؄ ���N-��� y���[��D	|WE��n��ʂJ���&�,�A'��MU��L��1����Z�Qn=��k!�:1�F�-�L)�}��o�B�ިqQa������٩n
�����$4�\	a�+��Gj}�C'��j���~T���7mu���/E�K���SF,F1Dy���4�z�$�z�f� ��{�,���=�wFy�fF�Ʉ�A�{�1�!�>5�cW�c)�0�lR�����3w�!������/���'�F�\��(rU �p�K�@ �P��!s˴�.�������Gn�>���h��&k�t�N�2�$��9j��������%'J��^&��V��g���\��a{u;�1��i+��lo^��q�4U��v�=�I���5��b ,W40�]r�
��	�Vp\`u!࢙��P��9���4��w6���g	�S6�9�����	��T�ʚ�E�ӷ��L��%GMͫdX��0�"�����"������+J��=����ZQ����Dit�T��'O#��%��ٮQ���.S�W��j��\�-��@�%����S��h��ի�H��"�"���,�C5�t�H*4�	:W0��̛�)h�s|�p�����[� ؜�\.�h�e]�p�_���U�3�M�J��ߥ�,,LR$~�*N��������sUP��Օ[�c ��r��vl@6��0�֬�y9�=�փYx�v.o�Gnc��O��r�u}L BZ�H��a�A�?$� O<�AM^�iQ$�k�[,
ң���F���y�\��#B��+� ��:�_/���ʤ�_�Nh!$��$x5jR1H�� ���:�aJ�0Q�ڤ#$��`X�N���d���AAx#7�!�A,>ӌI ��R�C������bG( �B9> ���"
��-(�}�G����n)|��N�dJ����|ֈ&�}�Q�߳@D��'�{->�C�'�Rq6�����r�$`��&�p�X=]hEZdv�~�}rJmh�Udw�ϛ�^�x5r��4�������'�\�{tM}X:�C>����H��#���L�6?'Mw���2���k�2�m�Ď���J�3t�a#�~sw��������19�}�CS����z�G�S��%��Ѡc����-��7?��f��\VE��꒞��F�J;��j=&���q���t"��g�3�2����9\z�`)
��u&<��zW	-��6E������=V[5���yH�?��-���H?:/��?�eZ�<J]�w까��ة[k7G^7cuβ������9��]�h�%Q�rg��Ͽ�>�c'�'Q��N�3� �Ly��Ÿ��=��eY4�F�~�>�\�S��X+J�_�� L��fnj<@��<�����s!����F�P�5���DƤ �=��4�:�x��]f��f�Dے���Ho���F5v:�S�.����e5� �Ͼudq�3פe8��qYY��x���!�/ʶ�Q��4���Z�%ڌ��&s��L�G��sd_A���y��v���ݽ9Y���:]�s#[�{�>KȈ��L<�0������9�����c����0�q]�Y.[�%k��7u����#Uq����?m���f���<�H3���TA�O;Y� ��T�����6A\�=�_�|�S5�!P���m�l��oп�л�á>�z�2M���?�=���b�U��Co(�������j�Agw�@C��՜�|������/3�_.ˢ��-4ꓱ�Q�ik�k�wuu�A8!�����e�@Y�SA.qA	���*�x2c��0&���J�i
�|N�^%�w $(�oO2�⣲a�HO�-oùW���>�@qCe�t"�=��f�A��I�p�S�¨���߯��u=}�v
��tE�z1:a��K�3�ڻ4�u�hT�?����ΖY�n3b�7s����n�r<]P\�E%hF:������X`�1{��T0�xE`lO�ew٣Hפˡ�`�Q�x:�=J�ѭ�C=>-�,���[?�������gDHX�RC.ئ�����݆QH�n�ˉ�,��2"�s������zbN��u��c�X~��_���P�#GV/�`$e>p,��-�Mȸ��M��r�a���y� x��8�Y�Q�_�F,7g!�I<��R�.* @��tsl�[w�TA(#������lKrgn�.���zs�(��'��q��Ŷ��@d�1A�<O���C�f;"��Y׃�ʚ�z�!���*��4�!`�Y5�l��7��e�9����:��yX��yu��M�dh�b3Q2K�YP=N�<ṟ�p�Qpa���l,�JԄӊY�C{4����s�