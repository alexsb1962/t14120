��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P:� Z` ��DJMS���Z{��N���^�=�C�;�H�P����h�<�V�Dqe?�'#��:�.�d�~\Rnd��~i*޸�!јe�h�Gca9��YX����B���#�V�,��<P�u�j��e�5�p$3���`�1)%LsӼ��ڌ��y�3�J���0��"����"�O���"GD�A�s�`�a�ۺ��#�!H餈�?zӘX�M������V�}��3"S6FJzͱB3�%�8�YC"�h�����_��̴;����M�q4���g4z ��Ko�t�M���[�A��_9�+�?KS�����%*ߤcՔ�wp-l��N��t�����S4W��2�Y�v���4����P�e3���b�����+iAqȖ����榒X��T��[�;U,0Q�u0����?��wL���|��$ij f�M��ЩdK�.�R�>1��Q��N>��^�÷�a[h3a�̙Ⱦ �:3��0����s$��7��fN�Y2����k���~F\pmw<f|�Fjg-��S�i/�����s��?"+z�CiTs�0��1�aQ���Pe����A#@� ���a��ݚF�l����+|��.�}�,(i�eԹPk~r�	�隕+��=Q�#6J輆��X�@������:J�v�.����$$�� !���S&%C8ͤ0�|�ͷ�������"#0n�����{Oe�;��lKa�`A�ٓ?A#�Nq��RCW��	M���p�4��|3i&�7��k�M�\��O��|fS/��<��v�?Hy��d�*�]����~3E�����9��F��P�x���C���YVMby��˜iK�6b��庲y�b�I@Q�C���Z|��AJ'�e��IS���7߼מ]�7,���"^kzl�;����\�K��qe�/�Ȟ{�f�D���u{��X 1�A#Q���
���P�C�X�M;\��Z_v����Nj�G��+�!�v«=!�giow*a����|�@�K(�$����"���pll�RO1b�Dp�[,}	����t��\S
$�C-an�:A�?4�/�E�5^m��ӷ��,��?TT���R _/3�v��):,�Y)�`����Ã�9b u� �R�Z�JO50�d�S�AN����-��x�{��t
/{J�/MXx�*�߳v�Y֍���	3���vTwWr�2��V>�k�B����5(���5*u���#�G7
�>��׋��[��B��N�Փx�*n����E�s���n�3~,+bLf�TK/M���O\7i,������R��w�ü� ��]T�j���U�=]�é,-�.'����M�OS�,Z"�B'^?���OҶN��F?���rw]0;,�6\�P�*��}�\�}��|Ns"���-N66���%�J��b�NO��?���ppVG@�X��R;أ�w+B�F�'uB�-#�%����{��K���1\�7��43��j7�rF���-�t�'(k��y_~V|�>)�����8�G�|��]f���"�A7D���ː\�Fi���C��F����ǚT
^�����E��swǷ�r��ܫ$��~6�ZR'3"�޻�^Cl�;$�}����t�t��u��}A��9���ùxe�����|**�z�p�`(i[��Dr���=�ɖ�����zyԷj�̬=�KFt%)}��x�n$a�?�W��h�=��AQ���=
��a *;���ݦD��!�U%W�������<���|4���2�T�=�Q�b�3����-���ǫ����\_�_��j��T��U�א6 ��xw�	%<JV�Q0"�i�)�A�K��׆�Nɜ�Vk�-�W��I���@�VG�v�4����.��'wְok�"��b}~Qō�p���5��|46�
���_��Z9��a�����	_�_�� ^�$u�_��w֜�t�J��7���9���V�כ�=�����\�п\��[�n�D�j��o��GS��'�x������"4Oh1�&�TS�)���/���9����� ��ܢ��޴��N$xQ��Z}�ey��)���
�B@ �l<zT��BF�:�c��	��������(^}у>�[�rJ}ū'2�cZ��]whX�e�@?���?��@!\��iJv\���u�5�0�����;A�W�<�m\v˿I�
�V��T��.g�L*������f����Ϫ	�ts2��gnI�F���](_x�y�\z*�%�l�!�9 UA�ps�O;_��#��������=&OGs>ZW�\0N�p��Ciγ"!Ef��Fcu$)Xm��O�[��3�JM�\"������l(���r{j��	u(��`W	��<���|>�1$�Eg&�51��}��Z@�g\oG�F��nw��'v��/M7.l��R1޷�Tн�=H@3Q��y�N���q��˒Ǒu<�U'Ȇ�8��]�0y8^��u�fo��拒��`+w�#iPY����N!T1[P%u�T����E���
��Ԁk]F42���,�u�z�p����1��jJ������`j��PY9�@B���ta�R<l獵��к���̫-zЌ�������	5�7�}��飠�[���zg�nqnq���	,WM�U�p�d�_)o���U���� ���D�9�1��@�Qf�x�GK�����!Hn! �z"E�(�L��=�4L�G���d7�5�e�FN���ϴ��)%9D^)buܵ����w�*�Mv:_7L� W3�ĹҎRl�"��?W�.����=)�����ȍ�/���80���nC*I�����ר���]]�ʨ#�N���{F�؊[�]{��oUjx�V��6[�W��xj�Ϗ��7��Z�h;��)�����r��XM�L�����r���"���Q=��K#�S_h�Z�)a/Y�]�ul!�;�����ϫH�5(�*���xIߨav��RB�"i��LR�y5���*�<�{�y�-�d�,��թI[�T��X����e?��<�r�(|�S_��j�}�`2�������	���-:�j��M�gRt�P]�"�dxm([���P.�	�e@�%�"oJH��(�1����C<�tw�c�����k6xN�*P��%����C��ruW&�bJRX;@�o�'�Kg������m�\�K+u�~���H�,C�xh �:.���LA��Ǳ��@s�L7�Jl������f�C8�kb��R��Q
3c�e:{�W���4���*����y=�Bu
DeѨ�8���˫��"ړRy�
���:��cu�{0��+��ԾB����|-����p���`Cw��_�}j�	��;�X���#rGc5��0� @Cq�;$�o�"Ӯ=u;�ҹ`J�$�lkY/2S
_�x!�ܝ��S��!͕*])H�����k�ue~�pM����Ȑ�kaȈ�.���+g��q��/:p�vZ&;;��nx\��v���_wR;��Y�;�&o�(��V��*Q�5W��4�B�[���U@��;-�*�Q�����6Qr�?���|6���/�k�� c[�c��OU��[��"�p)�E�
&FC���p5��R�ˣ�^v�y�y��&���A��kQ�Bʖﵴ0W�R$4_��d2�.iG�alf���ޠ�Ε���զeԚhyAP��ul��ua������2P�,�z��&G��*��c��JaC�i፰�J�аC�1���R�Y���l�5w^�[�q�[��!����Ž�;Ұp?)��!�c�dH٢9�)VQ����1�����WIŸK�nb��=�H��&��N����t����`i;Wb�_��*Q�q�������+�^L��E��y��J������nYZNƢ�<$��M�Q���>.��A�[����?�1T%��Q���2�E��x��C�2��6�U��Q��evO�	1��f\>�C4�-����	�ᑍk}���������g��7���������f�`]�s+�u�.Dk�f�͵���H��u?Ԗf�A/n9hq�]`|��S���X]�<V��Qm/���C��;�"-G��^4#��)|�5������s)�IL��hG~�i��7�g��sZ/n����A�ܽ�Y�b���0�[Q%�Q���˱e�0Y/���6E���t��^��o����m��e�L�j�]���@��	-�K�i1z%t�N![=�O+n��nn�o~���qi�c���lv��~�iL�k�j,�r֙��9�/���ֶΏ_�v+�/��H�*���m���ET���2��̵K�"�7xz��yb兒h3'd,�s���@������ؚN���h �^-�v�Tr|/5R>��\��m��@ATE��{馶�hF<]��ŝ���x���x���`q��o�j5�W��%�Í��y�2�猎F��9g &�~s̱�}r�~m�Ҁl�H��W��(t�mW���eY���'��t���U$�e���VZxt�@/"�X�
TU~a��kȻ�ݘ����h�ˬ2����3�j��D��aY)�i('_(���T��Zb�Zv����ΰ�*��J*��A�ju�x1�&2c k��z.�_ݳ�
���B�8��"��is�~�%� ��eϧ�{>�k��&��
(�á��,��{��~��L���2n`�&�����0�Z06�eɟ!�pF�	7h�|9��E$:�i_�F?���0n���IV	n����4m!�G����R�  ^i4\�0��S��-�+�qQټ��K�e7O����T�4%~Ot���J��G0�!���&�Ù��Y)��LI0!��P6c�8�Z��@`���Pq���rA �����I�4�(��¶���e@1� r�`��yM?�37��k	!#���tݡ�mvX�7���<��\��ô���?^�����#���p�+�+rj��jB���&'`[a�U�p#f6�q*��!n g�P����˨��d��W'V�HxG��������rŉ�ۖ;�Zz��Q!]^��«��hFf��@�D`/c�h(�8��ȥ�1?����U?E�4�泒mYWj��B-f�fp�O*`|�U��Lhr�B�,S�M��,񴣰��������n!�ٍ��u�[D�P~No��գT�����Y�4�ņ�
���k��5�,���S+�T��:%�8��M�|�J-is�xo}[�!�a����3p�v�1^7*}�3W�������3�a*z31���?��v���+��p��b��Y���#&8�>k�����F���\�2�Ǚ��Y�z��E�
�tW������,��z��M���� ������.�4����r6���'�����M�>�Ӱ"vA^��}���ֵ6N��f;�'����F���{��|�z�'#���c�B*�s�m����#t�m".Ԁ+H���,������J����֤ҕ�M5������)�?��	�aW�9@��-��4�&�.HU��K���K�8�J>N%<8�&?:E��ן����D�g���T�H���h䥠�Y��(X�oE�{���ZH��Wh���e�Am�}b�LO�C�}XX�w���]�K�U��E<G�h���`nYR��y�eS������^z[\���P��`�Zh���ݹ?A|���`��ۋ������ ��CV2hT>;c���T�d8k��7�"�&�8�y�����}!kF�۹ʲ΃/�����Q�.u��o\=�5�����E�:x�U��c�d��TD.ԋ��!{���x��~Z����"x�����ǼL7�A�@t�ud�t_&A��%�h�x�d&����	y�g2�� ��M�j=rxw��SQ=�9��f,!��x�ϽtW��>�3�=�0"���R|�L�Ia�|Lh ��Y*�f��aP���C�[�{�\Z4���?�=�NP�}"�?��[pw���9���@V���ڛ]���#���|����IEᝪ�����^N�����X��M�g�x��s�n��$l
f&�&��v���ڑ\1�+T�<薽sb�؂.��Dg�������e���*v��w�o�|us�Sk<ju����OŮ��;�Dp,/;hW��E&��)�����Zˣ��ήs��/�Sx�z"t���T*8O�� �%1���?XO��.8�[�^/�b�і�2��"&K�7>�i��~o�'�Z�M]�ٙ�g���`\��|��s�H�ޙ�O�+$��Ū��E���_/5�t�@���;r�e��&���j�vU1c�� �̌��,�[��U���#b	�EHY6��9����J��ő����/��$R��޽������f���dV���xu�bcM��c6�z�C���@Ew�*�����	��j��e�