��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� f
���O�Q�h� 1[o���zp[ �c�p �2q�:�W�9)�t�(�����1�B�ps�n�ri�s�R�ng~r�t.��:���\�d�@������P�R�;^��42��i�i�h���71���e�9��9��X���z�]-��a�g�g���w�4��i	�p��� g���؎m/�/�1��~�8V�;�$�5��V�xo%Di�%J��� rA��/h�}�	&�+��;��+�����hs.��,��ӌ�*�:6 9N'{������+�q���a��6�hszx�ݒ}�����_��9���*C��x���P��r�*�C���¶"�[fJ�c�.M� �3�ls	^�I�i~_G�X,쳳�V�U>h������.`e+/�|i��U��=��dF+n�I{V�Y�����azڬ���_�r��7�}P;�}{��+��,��AN��'avVhO����V}����[�����.�*���Q4�VB��q߻$�	��
V���y��35>~~��9Ƹmn"��)yA׵X���~�TO*�ad�m^�J��
O��f�o���sM��?��@��] (9έ���.�Fr���	6D/���e�L��Z���t�k�'�`xK4���ܛ3�/�d-Ny����Z#ŧ��:%�Z"�R���U���^4r?��4��Z
s�	Ȼ�#��x�O��F�-�⋀��a��\�S�����*���̨������j$��ʨ�)��i
Uݳ
k�i�?]'+��I��hk��� b��=�qy�Ok)���&>W�Q��ˇ�͑�/��es~�;%֫S� �f_�n~f?���Ӏ&\��ؿ�`�3z4tϴ�L*��O�%ȵ��H�z�aa�d~q$�Y=Z�iW��Ⱥ͒����>Xܲ�95��P��UU��ܲ��և>uh���� d��<N3:
t���O�t���C�>��UJN �3͢� �Җ����ezf8��Y��&����Q9���w�n ���'>�|#�W |�P��XW.����R8yhC��Qg
� f}+(%������$9s��5��-��@�Aj����Įz�ZI�K�����K����jCx__��Kr ���f�J΃���Bc�������Co�x<3��Tr;T���9T�eM�Gb���i�$�̢�2k� hqW9���V�6�����y�K�bch��ԕ��1�4e�U}��wf|�M�@
�R˃��m ����.6�������}���(L�*$�٦Y���1	��!z��s�F�7�C#r�ҪX+��i?t�4";�s���A�w��y���}��2��Ff����\��w�wAm��Iԧ1\���I���$٦���L,6L�Y���[��^<��+pƀ�7�h;>6ax��l�~���y��P�H�$��q�k����31aT��z��?��6j��oc��"w�'����/���Q��y��jr��������Z����dg�8i�{��P�U�O:�����ܐ;�]m�3�����݈�����߫�"	�f�uc^���O�~���YD!��0�ƵQT�gů��]�2��%��J������Q����c]sC
��Ji�N,6�;P��.�gS�EE�0��dP'�nl@>[�&�Ll����h�6�]/��i#(��]��gg�[l���ͷ^���� �c�� 
	6�� ��iOb�^ ��ɍ�"J(��F��8�f����$��3Am#�D���@�-6!�؆�y�T�~�������.�mL���)HJĬ�R^2v�xbR������F����������xFq0̛���_���C�h��;������~��8�+iV��O�Z̞���Q�p���	տ��d\���~O�S�d:�"v@�"@�w-ܴQ'+u�HVs#��k�IT����8�OX�K��� K�v�5L�H��-���Nb�]��[f��(���֚���v����H7*����r�@oW���#}m���%�I�k�X�ҁ�K�e�=�����]L����w�=.���e� J��l)�i�SP�=\��fiE��1Q��|m\2��u
��|�;wI�1:��	���(tY��s�߲ly6�5\z�ڽF�:<9�����C�?o�a�݃5���E�`k�����3
xJ-�Ӷ��g���nƐ�o�r1Z�_�+�o��.1�S'q��ߙ	��&^f(~)��}����D�ߝ�u��ȎT�jXW��n���փTx.��~)h=��Cb���Ǟ����'���I���C���ڞ���jJ�UK~@Z]�L���}��f�k�-Y��P��k�X�D��J#��c,��c���CR����m����ߖ��Q��b�'V�CW�r/���I��82�&#��4����T�^�!�pz�3sΧv��&�B�R�:���h����.�Gw��Xp�(���P�`���D�H��n^XX���`!�g���Y��������H��u�L^6�����A����cb��|�Y.���-�ìTc�-��$����S" 3c#)l�'�ؓ`��J�Jy�r#�9i�|�O�@���.Zi��⺮K�:�6D�μl��[��ߣ@n��F�h�n��^`�l���#�C�&r�Z�'N�z�)�b6��S�E+͎CD�?e�!�Aw��ܿݩ/_r�^���C���T��.M���][6D�����`K=��M*�����
�lo0�)}���O�:.��i����A�\>���}����m�Wx��D���e����}愝�?6��ob��$P��𩎗�M�Sվ'�r�G�x߲Ĭ!]^��S(�f	$���?՘nZ��쏳��a�չ ��|�Lل�`��`F��iT6jݍƟ�[�������^�ٝ���[�h/~��k �-O�B��Y��Z�f����z�֧-{Hl�e�Gm��}�X�2D�I��I��E"���o ֐O�_^py[�<�b#n�!��}n���ƓlF��y�z@G������?e9d՝��} l� "5�_��� J'_�� ��� OZ s4�p��w�p��P����,@�%/$����N�Yy9�4���V�l��۽4	g�����*�R���Ŝ������}�D��;m0�>�w;�q�x_ʂ�E �[.ܑ��Z,����g0�.]�!�9vS�K�ԕ�ŒtT���Ů�U��Y�sJp��i��[�i�_~&�svvR�{}8�32H����'��=�G8Q�8��q��JF��K��!�,�E�r&{�\������d�u��G藆mAZ�_����@��W���|P��dz��g(���!�{W.�漑0�ޢt;�=X�rR@��)�!���c���*�W9��:�
W�3)f��j|��;�Rp���������Jogp��������o+U��[�:;�D�����"m_�Z�֒�^���Mң�{���A)�<���A���d ��L_֣C���$�����1VQ�q���k
��Wz�� ���nB�{�]zL+l�49��z���(=a�
��r-��>�t# Ɇ�����h��9�BJ�8���_�kg�p��!�,���һb��%Uu�^��E&�&������   ��L�C*��骁-���(��lz/u���ߍI�7��c���W�	n8��+������Գ�
�qx&Q6��������������ѻ��cf��L�28M3�հ
8��#�'�?f`
'h#@5XS1�0�Z{�����^y��=���n/{�}�S�x0���B��h!�q�0K4u���}�ѧ��뗹���5��B�֤p/V���c��+�T�E���v��%��C�/��U�5G4s4TZ�QΨ����am��:�:`��j@�'�8�f�9ZL+�x1k�׭%�SS��Aw�Gb �EM{_�ϝ:b��7t�Tҏ�j����lp�S\��	��CC���7���C��[1�x}=���p�V�.�D#���+7�Ѝ�ǅ��4��TF�m�&V-g�s�*h���K�>W-�#���8����.���@;y����)P�P[Q;��}�`�
�FU���� ���Y����:J��:��t-�2���=���4h>T)���ut7r24_p�!rd1}Ѥ*D�	����爞Qu�C� ���,<	��v��K�g�U�V���h�%
ܧh�����`�X�銍��9(0!�	�����۶5���,➙�r�X'8�|��GkD�@��1U!�w3�M�S����e�RP?:�2����%k9�K�f�M������6&���ڝ�(��y!#0�9V׼4N����{�K����8ep�h#Ac���=�> �!X��%*Ylv�\�_��НC����mӑ�$�&��j����L���X1��]����t��Ԍ�xY	�!x9TɅ����0:���죙��A�Sg�ΐ��(�&��7�U�C��^�[�~��V.���<����#j�R���#�w��j0{߬�7x�KAc���cZ��Zڛ�<ϐm84Cc�I+eǠ���
*3c?�&n�&�S����f	������-DF>��h)Q��B�	�K�-�ͣ�,�k�p1��|3�ݦAV�M�8��k�޽T3V��d��Ѻx�Jw$Մ�OXFs�����V��=K��c'*���`�4�ىE.��7߇��B����uƱ����c� "(�ݺ\
���F�B�dB&r�W���Ed|���@��U�+���ZU&��9���X:�C��@Z��:���k�1K��{�ܿ� �������M��_��ciCmrڕ��Q'��,�������w������h��Vȷ1�Pg�Y-��d.gL��Ppp+(�r�2
��k���vU�P��6zM�=ڃx��2�abj_h���0�-v#;�rH��U�G[�BVF�3o��^y�����z��p���;<��K�q��+l|���w�kDx�4�Ejp����:(����;7M0QA\�g���b�6[��������0�I�_�C_�&�q��-E�8���z�������F���\;]i�j�ȸ����3^�~�"��Do�zbΪ9"߂�1��QZs]p&K��Z��t�� �tD�}�l��x�-�;��x�U��L�ܴ�P�1�to����Gcܓ��uȠ��R���@~pƷ<�Od�Q�zbM9�"�/�*��&�LV����ɹFB�4�.�R@��;�Z?�4��~y��gA-~d�|鰘�	�Pt�����`=����W��Z�Y�$�tԌ���0.��<�fP���*A�%�G����z�o�� ���zA�������+,ո�=9�k�>��E�	C�NT�5��,��3�J��7�t�8u�#�Rr���
.����0g���rEۈ��~��*��T�@��$<�n/lH�[�F ��?�"��LC���qE6}to�6���SD�����2ü{�^�nA�u{q���!9�[�A�Uxk�ð|�0���K�Oc��t�Z/�O�NW�T/%"��U�r�e:�GJu��w/�l����h��b���2C�����v��rDR:�O�;�+YWZ�>�ߴ�50r��s2oU'�L�u�3�Q��A�>ji����G�]T�4���񱟵��b�pݶB/y���N⇃,�C�T<E_��e��k�+����R��6;��\��w)A��Y�8z*��X4� ��opF�s/�Ŀ����n�
�\�BϞlRBE=k�Y��"��������
�Tf�C�+��a-ġ�I�43!�e2���|�=�L�.r������b�Q='жr��qu!�<U�d���|��R���M���:�F��������/�fI	ސ��+�A�]bK��NH���%�D�����5�vW|���R/Z+�����a1��0D���ҁ��G�6�ck 5�����NM���,s�>�rl���;�� HV ɓ�{#Q�������3rUN��AI.)�j@)dp)�� <k��J�L�?c�هsh�d<�
G�-�C�de1u�4���4�d?�NSX�=�ĥ#��('�'�0�����jͽ ���A1�N�}J��ܹh���2�?�6�	@$�m�9���T	���_c�/��6ƈ��F��ngMG�cR>ūA�i���@�rO�L��%��y�><��ش�|�������ì��|�"Y�]�$l.Q����0_d�;O��c_;���R�in�.�]ˋ�9��P����$<1;�>��*	{�ʲ��p����:�%���=ф<���9OMw��I%[��ۣ��ڃ��8�ߋCHR{nZ��6�dLI�l ���A���Jl�G@�9��Uی��=x@�3��eΏ��鵅и�T��'�Q�ݦh�W�u3�L�������8ob��фg�@������)�M�Evb�j�ZzF0V$Ixgj�U�x��C�d�� �����TE{j�k7��F�"��Sʁ��X�@��� p�,���C�s��=���@F����uw���*�2>(UZP�
٫\�N��L v����q2ժ��{��,5n#�,
�Bx�M�c�f=X�y�48�K��PA](C |BJ����X�,O�~[���^��Zy�&��~��:��1�6��Ƞx�.��Cy��|x��;^�(��e�X��ܡ�F�^Y~�N�t�V <�2N2�%o�o�_�N���,�؄?";/iʗ'�Ҋ�׋΁�g���O��K����>0e?G��g	��gG$�Թ�{}���m�`��QuVG�sV����*%������yH�@��9ŋE�3���y�]�>f�!Rǚ�$�U�m���,ٍ����)�<�4��}岹e�Z�{���v����_���#���N /�E�
1u����Ƕ"`ee�� v�)ݓ1 ����L'�U�R���T���2h�'�]!��@d���@+�s�j	�:��+��O/�I�;<g��z©1���~p�T�����40�*�9�KVa�Π�.[�ģ���PKMZB��h8��1��9<�Uy��Q�3#g#�&w(c
r�.5���h��9��H]�%�dHm��FY�j�I���(*��l��� �w6�m�|�T��ڑ��g3W[T��i�l��֬�,����&���(#]�}�-��T��0�ʔ�	�v�ԛO�B���oGK
�ٕ��P��'"-���\3r�����.�h�&Y4��;n��9�њ�]7����=����¾Q�Հ$֮�8��8�,�%?$��i�5B�ڶs��*^��5����^�2���_��V�ϨO\Q.[� �k������6�'� �W�XR�?�����*$��a��YT��T�L�6���@[�*�p����0 |S��%�j(�|�����rZ[W�~(, i�L�a��~�W?;E� �x��ǟ��sׯ*�յ��0h�ҭWj
XC�����7tJ���-�=ǋ�Q�����R\��/*�g������Ca�*G������,ZfĦì�˲�����P��ط��O��g��v0�w	�2\���Fp�x���܋�$��$Y��8$QT"g��\5��]yE��k[e�����i�S=��u$��~D\�z�//���+u�jEQ�~�%��	��ӥo!������4�Ht8B����I�/佌H;F?����[Nq��3%��#���0��%��J�t)����R���	��X��h>i��LDp)�M/�5�j����I�6�R#�_h5�>�}��Q'�Vtk���z�����&x�"����K����SU`H��0�K�ttLxIgLՌ"Р����쾼�q_�5g� �Q�n�&nL��rH��Oi����A�������٨��P{P��wypL�j`oBl9�0M'�S�qW�����h����P��g��a?�q��̖�|/Ja��GTO�ݘ@����vg�z`n��D@��r�"���U���U0O@�<��V�z����[�V��fM?ߙ�WtC�TS��ݳ�0���S�6w[Sᷳ7��E�^�d��~���^D���;�~_e/7�^�LI�b�j�>Hj��8`1預�Kv�{|>d�y�@�8yk`{z_k�!7W�c����8w#�e)	�}\� g
^�{3����`]����N�/z_��  4A���s�J\��z�,��.&�x6�<�2x�ᦢ!�
��u%g[/���D�����ʙ%�h����҉0C��Nً�Oj�g����2�#���CP[7�}��n�#p�1��f{7�j�Ӿ�ۮ��	u�����̳JԁѮ��]��e*�$�*UZ6ս�3��m*�������m��"��+1���; oJh??��]�J�	L�w��x��z�B0��U~�R_�[��i�	r�'���o�a`n|I�q�b��ֺ�����w��h�o9԰��6�4�0�u��j>8ؑ������E����J̙��?���i�eN����;"���"!�z�Nc����@�u�[�1���W��-FV9|�]�I��>Q6�%�٠�v���É�5ΉԖfhw�ݳw&4\����
_�GXm�:�'_���FF�r�m-|St&�[GM,��QN��1���o�1�V�8Vi7<�>v��$cOD���O��1����<�ͬ����ubYO��AѺ��m[p��dga�]\x��V$�Y}�F��(������ �6&�M��8 
{9���T�c�4��m�s��F���쬡2�TJB�B��U[��L^�ѱ�:�#uLR`�K������E�{��V4��R��B����L	�:����+T�	!֟�c�&�6K���
���bXc�	
��7��r[W:�p=0�.q��ad���b&J�`������ߴ�߮L��s}G�Mpp6Y��#��'� k=�KxU�&�8˯��bJ��b�0\�o_,�%�*	�f�q�/"�Cl>��L̟{9[�VSëc�u������\sN-�%�ōTţ�G]F�����]vu��� �S���6�<����{��U�@Z������(� �MV���;l�%M�됎#x��f�����{#4:�o����j�̔�\f���.�����\�#�nʖ��榚(����hڹ���&�'䜼�K�����l��I���Jb�� GlI��&��_�>�դ��}�*ȗ�ւ�फP�,�_PF|E�Ζ7d�$j\px����%A��R���y��;����&���ҫ��^1ً�Y��#t�>i���T�̑���b�("/�ĝτ�i_9��R��KJ��!�����YjGի )£��<�q�ц�S�e��
qq���IG=M��n�suJ	�p{0d�$�n�U3��nX�@�X��8R4hEPQw����B,��r��5]�e�o��&����G�$d|��fJ���qI(-�ϼ6���27ʞ{Z�P�>�9�Yǁ��]Ow:P��DkO��H��G#9G,��s�f�!#F�z�w^a���S���L��e d���B��'o�OKm� ,2��Q>�#h�{|�u.m߽P����U�[��a��A�R�]���A��i,É�=`�|��MzZ� x��[��4�+34�r���t|�0Ť������Vy�"�ä� �4�K��pH\�;��Ώ���!�u���1s�,T����޻l~����X����r�C�^�x��k:)sEA�����Ap\��d{7+����
�H�g�X;J�Fq��2���bh���+�S�$��ƴ9	-�B�S�R�V�z�/ ���G6<��t�U�����v�[���Uu�mN���#�ˁȴF�	z�x ��#U��T���DB�| 'K[�D��Z.�3��	|��~BJ@��m
H�q3L��#�7�2�O�M�auZ�9f���z"����+s���R��DFUw�kRY�V�e:�e��:���f���cᬟ��zq_H&q��i��^r�]�M"k%q�U�����?��'�!kV�Ș�����htt�k��i��;�{7�;�p^cS��&~����ʃ���{�	��=�r��n��1k�o"�hm�&-�I�7��������ze�J!=�i,r�$Hǰ�PQ���8N�e�׻�q1���#\�%�;�rsQA׋7��f�(D8�2p��׻����h� NM�I���U���&_�����1������#���N����2
94���r�Y����ʈ|�s��t�ȉ�Fȵ��DE�-������W��~e�#Wɑ(�8U�+�ء� �MAj��Rk�e��I\�
��I��"_sI��y�~���ҡ��%�e�{wU��V�{���J�	��>�C2K��V�KKD�����[�V��x��L����0
�O����pr�X쿩N��u?H���\1��������vK_oje���kV��V�o�:��ܜJ�G>�=�>��V!�*�߲)�%^ފ3�� ��?�+������;��s��ɬi�C�����]9�p+�'�{���H��R+_�DǴPX#�����JU�4⧢b��'1W���OV��O���e6ƍo�V��Ǒ��&��L��<e�xPFc��N���G4���`��W��6��Npͱ�F�0U�����]���Y���L�ϰ���2~�2�:	UG�b�"��4�%//�+`���41���5��/�]�`�_�Y,�Y���W�4�md%x�3J7�!���^��t�꫔M�Qfy��ϴ.�1�.�؄9�o��6��5��v�[�}�Nc�Ƭ�d��#"����sb��<JQW�{���F���#%�G)RSĵl�`��ӯ�Œ���E5������� �E1�.ð�(�����>q�Y� (�3 <O��]π `{��
Z�\WQ���0���ڷ�8�-��U[�����	
q	əlpj)�����n�aE�x�������f/b*�e�{�Ҩ���+-���1�Վ�O��(ٿ��,K������s4�d�`#�FW���/V�Ć��V�Fӕx��ɗ��g̟νu��t\�nj�[r���%y;�o�_""�.~O��s ���t.�6���I'��de�(�y`N��&�O���p�z0y�dv�$.�ֵ��bx�	[ݞ���4�pr2K[<�Ց-?I_�� 7���B��Wp��*���˸�9�U(:��i�%7�ogof�?��!,�6����{�������lFZ.��Y�]x����c�扏�����N����"Y�~�0��K��=��gU4��ں�P�(�0-��g	g��ig��M_��e�tK��Ս+�)#�Y�,�3f��2��*a��#Z��.K:|�"��s�W����vߒ$J���'	��>����[p�y�Oz<I�����SR��&�ƹ�Q��U4��
�%*/���,?�ζ��р��%���VN�Ԏ0a�޾㣲�U�\��E�Gp�����5������:�*�d��!�Q�8��G<�мR�#��LO�q�j����Et���|���p���0�m��{i�s��B���xOO��~��e�7�뫩
݅w�xslHOn,�W`�id���B���#�_�����\Fuv�x(��g{1��N��0	Ԩ�vo뫜�Ӏb�5�����I�+�<��h���D�23��KK{����3���"��Yܩ�J"
@*gǷ������=�����+[���M�
���fnVP��A�Z�#%\�*oaN����'���lD/����&U�����T,�U��v�L������Q,��1Y`O=������g�g\_;�y�@��%��9�6yM�-��7��e^dHc��4 �����ԣ�y~�҃�}w%D�58={&˻��W��ÝM�y!~7�r�zx� �!n"u��C�qLI[%���t�����{�!	7��t>�/�Y}}�7���&���%Aϫ�6"=X=pU�Ȯ���v�3��7@�m�����B+������e��&H���A���!?�>ʑ��c4*�)M�U<�Y	�C���0�׼[�����lK��zC7�#�|,ۥ쏩u3����y�y[�$vO
�9��U��E�#�H�kě�#p����B?��w;g?����F*���2�;�9����p���Ǹ�((�[ӊ�׺H�x� E�Z쏀�.�4��\OL��p�Gn��J���R,��;p�{�2����>~#�o�}����臔R��0��G�
�>{�d��ͣI����Y*��K�!;<Z1�H����
��;}����mvAC��CB��NO�� �����1����{����+�)#����tpaC
	@m_*��}�,�<�l"���qk��������#�#���޿7�GX�z����F�(��T�U�u)k8&X��*�K������4�/�P�]B�EHI�%��]<�Yz8A�%�9���F�ٵF�ʥ��p��W����n�9�r�޶��3b���.����N㱓O�T�'��I*7�"��.OT��3��6�M�ѷ��V$��kݸ�sϖt���O*#o�f~�a�ơo��=)���3yYm��<���f0��/�Ycb^��<�Í8P�[�ե6�m�y+�K�Q�0����A�S�m¸Ü�j(�!n��Џ�Mes�zK����h�3��I�_��QFRr+=o���.d״�J�b�I'��[��`D�t�_�і�?酶X�1!�[Az�N	���˨�թ�`o#����	��@��?{s��-�(Ҭ��n@=%@��;�aSZ��CɊ�X����qc�M���ӝ�9A`�5���6�<򒏻�����&G�$b&'>p�!����2�!8�H�-X1C�%�Z��'�����u�./�YJ:��(>�d}	��_6�*v�!"1O[a/�wR ��͔`���OT��Ü�ٙ�˷�5�5�k�c{���_3�z˕f�Aǀ��1Yh@�^/9���O��4W�J2 �SF�#ٸ��4,�� H.�<�����]N�+��H7� ��ؽi��Zr7�C�uUǳ� �L"��g��ɔ�	��<����G�+��Y��L ߢ�ٲl�|L�oŹ�W?�ѽ��D���������Kh��m����$���s�т�e���-�ɋj3�4>44��V�3��>�j��(�	���8矍��(���F6E��y�T��Ezt�KJEcCSXe���P2�K��4e�aĒ4��⃆fӝ1�����!��#���ܿ�i/����k�����d`$h�����
�'�R6"���X����X>��0�[�v�׹�W�PGZ�f�Nu�'�������u��
~hQ-�\0��6��k{��4r�*��������܌Vk����?č���Jraj�v?M/�>�d�)�P��j"�?S���a�JY�*���D�l���N�4&���;��Vph�Byб��a�c+�,qs�9�
絳���0�=���rk�n��dU�.Rkb�re��?&���"d�Ω(x�(�qw�#�)~�S����N��� J�Y� ��U�LT�5[z]�VrE�kU�;��J��<h�V�syÖ���;�$C24�#���-3��1���a�P4[V�;�j�@��9?K@[�r����
_� q/����Sj���{,pZ����/� ���hL$.'�q0Y�)�O�/�b|�)�_`_u  ��@2hM�i�C�zoW����I���A[\Q�l��8��<7�z���I����b�LD���{	�iA���l�{��4Q�9]n��hH��|#�(�+swUt\S�kj���}�y�@�5���|>'�۟��|�M�dd� X���v��x"ޜ���:*�d�%�@ZU�\I��V���|2i�H��}�&��s.p�8x���lr��Z�7̼�� �c��a�!�6_����u�enf��q�W����!A�G���\�&>�95de�8��bx(��.`{S_�����u�i���f�ԙS����zD?� �ԏ����&&w㧛��g��EI��W�u�M��3����1���x��+�Ϟ/f��ݴ(� �l��bc�h�>���gm��V5 +��<�R�q�xI�`ڮˍ���v����vA���*\pW�-E�1/��ąQ���O�/��wp���O.�u�i�@p�m� �h�QW���o4�L��r�3H���kF���TJ�E�{��z�W�x������&�0}�3a��#�+�c=��4@A�7���Tr)A��Љ�!kɧ�3�S��h1�������H=�>�'
b%x抰R�N���k��4I0ɮ���d��B_����5���t�.���gO�;�+(��>�P�ǲL�ۺa��tK-�oſ!>x$��j��-�k�l�q��@J��m(;U������|����u
:>���"��ot��s-ψ$`�x���7.�3/�?&?�����F��C6	���v'���xy���m2[Ij�o����nN��+����9^�b,1v{Nt�*m"ݡ�����W=2`���q���������Ƴ����h��ig�s�&6MUe`И�7�F̓?D��^Р �%V����
Q�#9��4���C7��gw|�-<T���z���ac�L������mz�v�6�L����>���w���uQ.9˨3��$��]X^���ۄ�^g�8��-�[4��s��'i��%���u�!h���\#���;��p���vѷ/��
� �f��p8�/J:y3���=[��0=�X��XHw��	�ԙ��H������]ڲ�ːg�h�{�e���Rg�c,���S��e=9�|/{�]�����^�<�~"�A'�Ѥ"��-MЀΠӠ��A��u�����M�n��W�<L���E �����Y�B��a�sht����TZ�3fe>�/�X���������èJ��
B~�N���Q�����=�gfa J'�-�	��j�Nڥ�J�"{�96Lk�Ă��E�a���o7� NAo�i�o0���W%eg:+~w�,���:�i�e5>�S��˅@���nb�;���1hԭ��Rd$߾�n�v�ZS����8��-����� � �T��W;_>��[MF��E0��<m&�� Ύv�� �4	���Mъ]L(�wC��n�L\����Y�|����Hky�M�P�S5
�x|��v�5�_��%�����ъS(��*��-GЉpq�qr��M�A���9{Y�M���޹Vu����"i*F�#�h JM�-@�֝�w�m.�����+�.Ã�B��h�_ĵL� ����]%�-��+6W�!���:R���;}��8?+'A���u�0�ԑ`=�S͛ϯ����o��	��hS-�yVae�2��]j���z�F������:�W�\���p�mX�P$�����(g1�Rd��dyGpc��Yy���Z�,�HǓ|���bn4U-��ږ �5'���鏿�#*c���	"�>��k*ld&L�r�6�+��j�㋑`���7[+�5$O��k�p���� ]��7��MJ�C"M7�߫n�J�Q��aj{����%�Z<䀪Ҷcd7����bé���{?c �;��	%ʒ�J�kK�]YWb���\^Z���	JC!���`׭���6�wn}�{-.x7��3c��be�OD�>�Dd��5=�&=�۠A(�}~����o;��1Ճ��mX|��\�J�x�=h�fS;t����4q�����Dz��;�s�/q����My�9<|��(�:Y�9;��û�*m����I���9ͳ��N|X��!'�E$Ѵv�H�lG��R/Y�B�D�Ƽ!�o��/��G|�(�藣�7a�Cb;��Ҥ:sh�^3�D��	�\-��)�>�����F�W��^����R:��â�G.��R}�}Z��y���Ο�%�j�t��>P�]P���[��f�w)#�Evj�<��SLqHtO�`�h���n�<��G���4�WH�n$�F��i
t˿���)��Z�'h���6�pr$���-t�9��4V�#C��d��B�\[xo5P�|���9� �MHxP�c+[U�#��X���J�6�U���'����۲�ڠ<�jϩ��j��Gbv����_�Ǟ�XV?�'�o9������-��ރ�<�a)�H���0�����ﴸmR�ٙ������0��!uO�]��L�|�j�q� �N���� �P���;d_� ��+��"�cq��<� �$�+��Z��V�J�=�ֺ��:�BTp{�5Y&�p:��іL��ݚq�Oc���AA7�����s�H��<����-��*~)���tw���f��zAo�{��q+=o¯�
Q�����i縍b��[�q��3�yy�#�FM%���6�,]�_J��6*J����្Ǔ�qa(Tw��
�`���SN�xr	�m��>d�xx��N�����yن���\蚯��hqK�B)���+L��"�!�zO}�&B��\�����XxNqi`��1d��l�Ņ����v���ш�ϵ����{�[{��j�|�`^/?)�j�*���Ng���k�m`c��+~�=n�E�i��݅�/�fP��s��Q�j�����<�4�'��F�K{:?M����l�+��1�S�S��g��l�'�l\��Q(?|���H���w�y
J�n��zA�	_���{t�M�g�N���D'>�� Ǧ%��	���v��y���#dC�ٮ���G7��b��Wӽ E-�Uĕ>�i��;S\��u��F;	pR��}�n��	�~HC.ol��{t�9����}�IF�&��B�wjG	z|D)�p������#���+����@�c:��(t�+��l:,��it�h���<���[��ˌN`�t<�~m�ޝ���ܕ��-���Tf����K`�K]�1��&̖ѓ̏~�J�	��5�a>Ҷ3��Q�������'�G�=3�ea�>�4nU�1/?�΄à��P��c����{���ov����p��5���7�𕸛�j�m����75CٝF��h�e*��,��G�]~�X9@�N�n/u��Tt��ӝ��U� F����(D4�58�ƽP�>�'�CHJh{pI���y���[�������3���EH0Q��H���__�2����fI�?��Ffֿ�9"��Ã��^\�^� YH��N�=g�8����KƸ����#bh����Q�l�i�(��\>3-"���$w����5�f�w��T�Ԍ���uT�s�g9�C,�#����.֮D%�_?qbzUWz���\u�E�Ś-��i�A��?�~��K3���X��bdS���Q/[{��U^%����V��0DFǀ�q��p�g:�.%�vT��D���iA�Q�͘:�:�	F8�1L����~����r��3��L>��[�l��ORD�g��m��a�E1����ʓ}hڊ$���CDK�@��Ztτ��ipTW�.�`�V�HEU[A#��}ڲ���H%��W"އ���<�ª0%�9��"H�} o��Q#���i�)�SܳP���nȀ��b�������2i-���r�ӄ�-���S���p~-ҽ�DF���
����2��S����dy�Ոy��<���qo 1����2��H�h�q� S�k@0�,0X2��4WBq
�4?D��@Mwc�u�#��~���R�a./9� �6y���!Y�"��a��,l4���K�Ci �bEKmBVd�A����Ilr?]�U�r�('��4���H	� y=�(K�$�~ �,�]ͭ*9ۖ��Ƣ�2e*0�닎$-��N&G;k���3ibb���O�7���A��jTU�cE\���yPqG緒/k�<�Eǩ��L�Eܩ¢w������ܡ��H����\�aиV<��^������p .Q��Z#9D}��2�z�-���q9��Q���4�Rn;s�<���m;3����K�� Q����P�����R:�UK��-�A�¹ws�j�`�M�,���^UPժҶ��f����鱁��抣���B���K�JR�D���v=������K�Ю�0����<IC�O�9M*h�}��(����1#���Ǭ��^�b�1V�o��`#�j����F_��G���}������>_yF`L�پD*�(Rii�F6�)�/ac-�C�#�g�ؐ���ꟲ6��v��F��4{c&�;8�z��Z����s���=��I�YCN՛���D]��/�xpL��5�vѧs՜���p�k�[n��:K,@
����C��  Z�g
-1�`�x���j\$�?w�<� �HL��S�m	���=�}���@29Śzއ�*��c�X� ~n@_�U���I`����E����֤m⢸���/ ��_;�6�1���a��3Gp�Ɉq�=�Eȭ�Zum: U�����[AO��>�vN��$�eo�T�p�����=4�7�|�w޾>����� n�o���)(���4�>~�f����ٹ�oD�/CM���[�	ui����@�"����"��F1p�����������2��	u��@B�ϰo�'tY<��m���L�-Gy,+9y_C�~����ڔ��d�k�'�vGf+��F��?�m�kì�)-�&��`��Ⱥ�Gb�V����]��8Eh9��N��ZgWL�M H·lS�]������}[gv����"bq���&uh.S��~�� z�׵�����=xQ�Yv�N74�J��5��Uh�y�?&��5�R����}J�f���N�&�_���{��EcLX��.��L��"�,����;�)�37�D�6F@�p������%�拯Qҩ�l�KΕ��/�{v-~
����Q��7	J��W��6�g{m]��c4TP@KE�O|{�������Dfѝ�@Dą;�2� ����-
�TD��:;�y �Z���%߈C�z�����Gbe@Gv��	e83K9ĺHb)���R�r�������_����Qu��c������;�I���$^�%ja&��D|=������QR<�}�k&�����R�[��C��Ԧ#��)�ln�e�a7�:��\Cޝ�Bj=�R�W�� �3rX:�I��3M_e�rt�Z
����K}5W܌b��"cXi�(��@)��ߟ�J���h��C���}{��;c���
@2�AANݵ�Kz����:�U���3K{� �߹���k��tPIF+��߸v�c7P��_K�c�*˜��Bw՜@���-s��c�γt�%K��3�DRr��x�ޅ"�$
� �ujϛz�o};��Z�{= ������Gu��뗨�X�`��d�B����|�~�`E�F<�:m'����ݵ��