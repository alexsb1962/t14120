��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��<��T�@d�Gu�!�h�����j~���C��P�Rc���FfxXs�� PC��԰�O����p32iXA�t�"�Q��&?,P#̓�*eA�9T�x��0�8nVHAG8A��J	��c���G܂y��S7AC����&� �?�,�	�B�Ũ��aU�P�̧Θ꾸^�����\�(+��F�I�j�z	�Ϩ��y�g�8!�2���%Q���_�m�$�x���b3,B�6����9�@fZ{�G?֔H���R ���o�;��Hd�����������O��3�m.��]k<�B��I_"Z�L2��:*p:߶����aȈuJ�L�_&�݋�w�����j3�����:6���Ɋ=�����e������0|)
m�N�|[d�)��H���ڵE��Jq�)Tꗓ&�^`kC��O bC������h�j<��+�E�v�)��G�i�SN�p��x��Ǔ,�z1��@��t�ܕ돹S��Iເ��8�^x�)�=��V�fE�s��a�3c�e �ɢ5xE�'�fr&��W`��r�E�m�_R�W�(�|1��hR�%�O��p�ʼvkn��I���T;6�<���d�Gt����d��qkcR��H�5=�E�zD�YX�k���B��&+8�w�}��3V��Cbk�9G��3�����h���7�#���J���j���d�]�O�x�kk�J�1�A_��,�&�:�C����+S+�p�R�^4fN���U81�{^��_!�R�q�Da\��p��{��Ox�o��,ȕ����
J��wܡ�V �p~�P�l�}8���KP��שX���B֬ȼ���_�R_�?Pٷ�x��4TZU
�4E[vS���J(R�v��3��C
�)�2B���a��+]+�Qjm������{��]��֘7L�D�,@�so1K����7& H��k$%U Oh�v��`�(̟�\�*�Yw��dg8�I#qs��t��YR���"���K�`������D�PF?L�%A>�,��l�4R��;��8�����E"�*t&<�(S%�Ѱl���m5�k�%vq��\��V��-��-��ڲ~5 ^���8��q#=�tCnI�Y�ٔw3Һh�cn��vi<ƶ�W@1�I�=��i%/sY�y1(�E4��0��|w��ha3P�n��ߜ��=��,�����m�U��x\���1�sq�4B���A�͈�o�Lq���x���A΀#��7�m��@HO��{z�ٱD�����:���%�PH�l*	|�	I}\��	i�!$%���AN/���ֱ� t�����nZ'A2?58A��CR�S�Z�� M_{�jd� �yB���,&�妡���r���Т�r�nl���қ؟U�F1�4����Xb\\��I� A�g �mFŒL��66۹٢G>�4�j&k͹���`I�k]�&y�8Z,W@�g��z� �GV����l�2��'�����2�>���
��3�헶~�7�א�k����O�LM�B�S��jq�7��������v��lz�m ����;O/���g�ǌ��u��7?��X�!�g�Cq��&���o�3�`��G_�|��T���D�lǦ8��6K:iC�=6x����Ȏ�=���w1A�n��j:{q�5��yh�ktB{Z��0,��Y��&,�t���lT��1ؚT�ĺ��e���e�A�sʡ�z��O�C��E��g��b}C�5� ��x��A��>�)uU�k m��tpO]$�tT�W5�Z��z��,�6$k��[���%۽ym����+��}Rqq��nF�6�8C_�ʌ���� #�W�k�G��5������^q��fS�bb;��s$��X1٬d�T�1:���{|���|�+���U̗i��4<R)ͯH����5�W���z����|�@��!��}~�lEo��>%F}=�^�
����$��t7�	Q30İ���o�:�X�Ak[�6u��P*�O�+����%x��zpf�%��
>�&·�K��8J�_e��!��RX�ަ��Ԛ��w
�M��vU}-u2(�Z��/q��}.���D�LՏF4�&Ҁp���}��E�Ih�ʪ0�� <S+9���C��'��<�}<j�����4�ps�LS�*!�����	7%�aU���>k�Զh��:���˥��{˲3�<`�w�'���8z�I��nu) �Q��^ސ�\��6Dz���WBv��k���=�ǆ�Զ<�O�e��=E!�@H���	w١iڗ��d�� P7��3��0���dجEU�\Q� ?��Y�v\��]9I$*�����A����)H\h��N\�?�*�3� OI�9�? [u��y�&i���#I���ٴ��<��j�G�u{�i����!cf<�PI��Z�9΁��0�LzC�����1ܞ�?#sQx"�4�	�j-u��F�?�J$4yJh����!�!��!�3a����;p f��jU&���x|^�u�-����Ӛ2��7�2d�&�d-',�ɔ�d� ��Es^Ň{���D�O�b4��H�]�Rs�%��.[ǆ�q8)8�:2p�gh)�1�ٳ�!G��^2��K��P�j �S��!D��-8K�.3�0�G�-���=��*�ځ������/Mb���U2qد�1����)r=�����]ԵKO��ڮ�'h�0}?0&��"��[���G O��B�(��0�L� ?���$�G�� 6Wc�Lajj�rjX!�kyhP�eZh��&
%읊�R���O;����_��Q�{��r�,
��CCc���S��e}�	ӗh�Q�f�K�f��|E�n\BdAAX��c!�y�0�c���$=	\gqbAQ!0B�e��jTUlOw��L�xY�.Ոk��DF�E�¶��C�#�E]��Z���X�</���g�[�-�8��h�;����H�n���\���*��7G��1��:�?5�����]E������á�i��
�B�ANy{A�j�fdU��.�a�Kշ�y�Ki튞�\�Ϳ�ڼ!Բ����sN�/��Ґ���(�_3 "4\���U2e�ƒ����/�C�qP�R2[�8hfY?T.L�hRu�c��b��1��.[ݛ��3I��V�۟�Xc�[zֹ�2'd���ņ۶b�K��@1Ћۼ�J�Nh�ih>�Q��ۇ�?�i ��PZ���WA�?���C�B�9G��Ճki�5U0S�<���͡�F`�����#��*�-��և`�S��?Si�-s�V'Ehp����4�#���C�|ݮ����C��!}"F��=D�U���ÚМ��	�����`>�+Fd�/���B*+�"�t���"���Nr44�b۱��y$r�z�F��	M�`[H�(�9}�eJYr��y���̇ѡr��o���\��+�i�SY�(&1��%��{\&]
4<��;u�����x'8�����ia�0�{�ρ��WZt��U c����Qm����;PO������네ߋ$u��0�{H?>]�J����X���S�U�}(���+���a1"4�7�%�H�n/L���0��������yvo�A	7����B���~��+���Ƣ,5.�ԯ��Z'+G�Uh��֍V��uQp	�"	0���d*����I����j�Ü|�{�x,	��ƆpU�!>F�㗌�e넙썊GxV3�Z5C�/��ٲ7�z���t�РW�r[~G"�%�|0)�L1 \8,
z��xɶԙ�S�7��2s2�I��h��y0�� ;uxO�^��3�[p�@�65���܌�8��Ы6N�ѣ�S4�����GA���j�[SVa��h�����NbR�Y��Z�Qۜ+���*�!���w������B�%�o��I�"84Rb�٥4�r�J�3p�͂뇂��G՞��	��$<Z��U�%ȭ�ի$��G�n���'��95���U� ��h;�5d�UC�e8N�j{�������Lf��z��\JrU@Km>�Ӏ+J�d\��7%@}�T*_���
3#��b�*r%l�� �F���^j�����l6��4�ݍ�c�C��H�1us�������/1A�|N��y+(PW%�&f����*��a� �E�fm N*,��Z�����&�$!z��fo���5�gP����6l�lڪ�P�Ji! �B}�$[>��w�T
X��i�*���4]
	��'\����A��z�qۮ<�csw�;M�-�5��
��=Y���$[��8ێa�UvI��[Q�C�^�W�t"��\��] Y��,��F%D��*/���'��Βp�P��c�G���}��3~�/�$����G)8�q�;;��;�N����x;XԄOt�������)�S{�y�z�qO�{Mϊ�&=�T{�ʟ��~�_m�7�9�I����}�FY8��!�%�P`����k�ӘZ-0'"��Ͱ'�ɼ��/��R�Jư_�Ng����4�C���Q����~�U N:%i�q��*}F%�-Fn��HU�  �OQS�NwLի8M����N,P�DB�m��;�QԆ��x��3�&�hH��!&;�)�.�5�b���?����bӌ��Cy��<o[�SE���s�*���E�p`;/��׏U�3[�q�����[���= ����DeCD�7��/�M����lW��޴g�9�g����F[:'�=��P�l�fㆥ���{�L�q�#/U�e>끢B�>q������e�s��=Ѻ�~gXlٜ4������)H}p5�)~�,v u����ύj�N�$n!Ѹ)������5��>��~5f�J�'��Ҋ�!���#9hl;�ی��K��0K�l�)Q�|�RP����X�|d�e�;�����������N���A�-�
�ۇнC`ttg��6O�ʷ�!	�D�sX�T5S��\�/�c��xJ�ϴ��ߋ�*�z�잞���(��L�E���s���:7�{J?���^�N(��9���M+��g�\�L�Z{/7��/Q � ��;`�5��T-N�r�!a�ȭ��4^<X��Rq(�_�Xo��:y|�NR/�jo&gB�y7��|^#�E34nUZ5�m���W�w���������jS=ٜ��k�%���	�/���+^[�Δ��
�뮿��������,q}[,��E��:Guض�&��G�|Rgo�T�@�Y�A��aI���6&X��tdə�S=�t� j��VӦ��@;�Ve_��2���ep�p��P��MWƭ�I����i8��t�R�j��zRO�8�K:F8��M�2ۥұЩN�^կ�r���[=�QDe	&Aa����{������<y��
K�W�H,�D��n&v���ӭx[]�`n���U��`�7�Q:�j����B�)��7��������"��������� ��܀�W��iP�Q�E��-��r�b\�w����Hi\O���4�Գ>�P�}7��՘�	f��w��GL�Z�/t�����?a��f��`�p%��*�� ��?��?�g�H$�ٵ}W�m\��\�
9C3n-ܫBe�M������Am[�k�&�B�@[>��/���j�9�CxM���a��\�":*����?�9K���I���T�5&H �cg�hN}�-�����du��ş]����[��Y��"ዳ���չsA��-z(���n!�思¾���hP|*�݈L��=����8'ƲX� �\"	;YL��Ws/����G�0`���a;a�՞�L,`�?A�N�E��"�Z讱ȑ7@Lfg�IX՟�de��I�7 �*ȏ [Ұ���G� ĩw�S�05� Bߡ�n�qv_QVz�>x�0`��|�oV�c�1*Vg%���2�x��IRYXƤ�U3�'X�D���$��@��w�+��d0�?�k��ZK=���&������L����V������$u���;/m7|p�ٝ�zR���	pF�!�����[�1j8���r�^
2Q{3!.gJ��,حA���.(G�=s!�d�-�Z�f>3Hq�lZ�KL��`D�w'/��U\B���c�Y
���a��Bz���oa�Q.�xL4�گ玲��Ձ�o���>�zD24��S^��G-H;���dyn_�c����8e�y��9}�5MN��]��d̘O��F�\-��+
��8C�ݗ���9�?�w��� Eja����0̂�m�,bߐ"T�ĕ��㝥��q���M�.��Sh��=!��pt�5_0|_��{�1l���Y�s� Nqe&�A5%����9�2��˕��y��r���3N4��;���(c�nRrc�����pfb�$W�m��u�J<��;�Dh�6��>¨�d�ۘ$Y�=��ʲg !&�ٲ��J�Fʪ���%��3g���ǃ�pH:v\�=���d!��f�l���'��}������\��<�� ��;�z	ϡ�;��5ruvw)����p쨦��|���i�b�3�����0�R=]Z�L�O�7]f�B#�����tE�으�z�1���m�(g�C2��|ԢA��<�hxC<y���-3O�U����0�O&�W3X�����~ܣ�#I�%TH�͝��������]������M��''�8�+@�� �b��( N_�Ӷ��n/���<�uίM��2%2`T�NV3Lr�(WI.@#AZ$(}F��ק��S�m4I���U�nl�=�Zlz3�������'�����##S��d�I��{c��c�5���sB��z������*�k=2,�y�-$����W�Bw�ht�BPl	�2ig�4l2���7m��%O��'p��u��
�"�p�65⎤Ȳ{�M��"	�x����MiG��X�F���d����=����ߡ�x���Ƨ>�h8Wk��vW&5i_O��Î=�;SB�����T㋃�Q�6��7�T��Cڍ��Z�Sd��٣�����59���Z�;̓f8 )\{F;���x�|-�)���>��k����3#��L��.�7��V�����,�(7[�,�& �D�P'I�G�S��c�"�k�K}�!z4h�����"�$2��rZ�k��
��v32wQ#����q�o񳳀���q�Uͽ���M"g��i��v���s�Cnt]a@C �	ACz�S�`a	lh�CR���sS}�q�]
}��f/F���pw��3����J��s��a;�K��.�?���>7�*��%f铜�o��S{`IS�%�0�#�4#Sw�wi	_�K��j��@,� |oJ�q���An����эҵ��:*
�\"�,�1�x��w�͝w�1�.�����x<�Ac�����g\㱅�J�3�V�rL�	4�9w؛����Ԡ�w�և�/��Wi�;�������{޾�'���؋+�zi^U��Ё�n�?Lg�kJ��U�b�S���#c#�4�W�Rzs
4%�c���,E���#�\�.�:��x"0[��Y�#��j���fN�8�U�&썒j�*6W�p��F�5[1ߧ���u�����bh��(���8Rqf�C���H3��r���D��=�QT��Op������Q>�����v͛z�g0ݿ����^�<���f��h?�����yC�u��6P�������!\�ANiZ��F�G���\��w�n<������%��]�qJ��B��K>�� LK zޔ�	�?�f ��~Kn�<�d0�FX&1��wE/�G�s�ߋ��[1�\�Ϗ��ej�	��vK�4�$,�hB�������p�W��fFFT}���tHj����%�t��cy+n�_X���z�����B��Cs����*1���Y]�=?`����i�����>�F~S�u������ߞwd�H���Aw$���i,h�������^����:n ��`Z%/"[�*���cLGo�j�s׈d��Qz*V�Q��Hܖ�[�
NMS=&]-��}� 颤i,�H�dlݴ��4�S�:/��~bPq�<>�xO@[`� J��3��� ڴf�@�._#N�P�O�S��1�����1&����y���%�u�������>՚�:�,݅P��y��=>Z� ��ENH-���U�c����a�n"�&O¡��~6A��X����WSMIs�)��$��^P����G�a�S3�F��DI��z4A�G�TZȡX�V>�Smɣ��ܳ�I6��ּ�W,S��j�sѲ��uW	;���V�)�E����?M��8�#�� e����#�;���<��D�	��l�(~���>��έ�� �B��W�s��k�����I���-����厽����U3N���X�4�l�bs�&�Cc�lǇF��.��"�h���)�� ���TG�-��˲�:R]}m�=���db�f&k�v��Zцs,Hj~�*R$m��� �K"�}x95^�6^����x�K21M�x�5[4AxG����OO`s2^n��a�5	�ɩ_{;[��ݙq�C����/H~����3�΁�Pq;��N���\(���C�߽���Ǆ�@F���C��]�iw��ܟEb祧Q���uAt*��5�z�a��h
�Q��\���
R�`��Ѕg�ԼR��O��^����0�U ����.��O�u|��6W��b���{��!!��׽�)��q}���Z�Swƪ��2_��\OF�g�E�z�@���\�NΌ�h�D�sS��K�	��D�����+�(u��K0PN�ԑ!c�&[#��i3ˉ���b��u����ӽ�W��.���@�[3��o*�Y$��,�Y;�nL2n��Y	�f)���G�s�\>6�5�$�0�!NǹAU�aNbP���Q) l���8$��Dv��YD� �z�S4#mF�������sܼ ��@Ӛ�<���[�(B���v���P>�Jf��ę���R�@���j��Rz3������&�!�n�ӿ��%�V���˒@��1��f�%�p\�;,�U) ��Z�(�l�%@!ǖѓS��v��}�Z/�z���fVx��~����7=�kI<����na]
�teN"��F�c9{����D��H�izp���m�j~蒑;��$�#ňm>��\�2�0����w�m�N�?���9�
p�\������J�%����&<KB7A�bIf��M%ٲW���ްUaڄ]��d���=����)��E!N��ꊄ!������}H��y�&W��a0�Om�y��4d]�EO.��zZ�J���b��a=L<bZ8��}�81aB9�,鮄_��μ��Pr��6�AaR��9i�bE�iw��ݗ�n�PD9}�igj2iig$ ��MCVU�&pW�f�^�K��8��)b�Zef�Vq&��Od,���c̨�P�m�2�M(dţ�MR&Mׄ=�U���T�s���2Fr�._a<������v1_�}��׿B��V�Js˂�h�G#u3��rK왃 ��%�=�VmH��vMJx�@�ͽ"�[�G�M�$TFS[9�NcS����$��Ψ�jr�8݃|�xțJ̖��	/];��w�f���TX(�i,݆�P�\Y��ȳ�:N�=Nw�1?N��o�k�׸$EE'R2+�{�P�|W�n�yv��ዓOq
�\'��B��v~3�醙�<�Ģ�Ÿ��mԼ��M���VO�-�H�N������h'4��k}�-( ��?3�)�N/���VU�i
�6��-l.�!'e�: U�WQ��xmg!�<�{e�%�� ���P�F���ܨQ@�jKQ�w6@��]ڧ\ܷ�'��L�ѱ� ��w2W����{�3۽	�ob�4A���$��2|>�pQ{�Ko���~V�ޒ��C�ʇO�ױ�Feu!SUf���lx]���7��d˥��	;wV^@����r��c&N�Mv�itr��ҁ)+�U��P�1u{��q��Ls#��;;9����^�!��Ǘ~��A�O<�z8J��ō����	qJ�rsw�DTSN�k���6x?��NM�\Ĳ�b���k��l;���,��][��QP{mV�al3#U�Î�|�a�"ހ�0k��@-��X�_�`���Ro�����w�m^���<)K�k\}@�xz8�!�\9aw{�c`�t�7[9(��8�Lbs!~�4�Q�������pcL�e�N"~�KO��*p
��KD��i�	Pouk�A�����ef�&������~��iO#%E��v�9f6",�Tr]u�EE�kf�C&��Y��"||Y���V���yq�B�[�	j��y��<�!�Y0��µ��H{Dx%���Z�q��}YB��G��wù=�^�k�w����q�,xЗ�@����{�,�ˠ?'��F�V���y�|'�F?� 4����^�f�wZ���\8̧�1l��u/C��	�5h�/��>`1��ΦF%K���w�!��Eg��!��6C5&����,��
D��v<Ű׸�ݨ���cp{uX7X��F:�m��ܖ�H���F�}�{0��u�����F�p�˶��� *����B�A�Wb<fQ�g�o_�b�Ue�l���2f&�x����:��sP� 0�O<EV��PI>u����(z�ǎ��x94>Α�oHY�#s���[�ֿFfgG��,����a���>�2=��;b\�4�r�K�^���ӭ^�eD��x]r��(_�m�;�x#a�m��>�^���<i�Y�E��^L�!j��onF�5�-�9��Ns���Ք�U���)X�\����m��5��R��j�+�M�zg2�cN��V�N�+r���"oЌ���h�V\w��� ��<��N9�c�U3��Z�+6��,�ރ��Q�JV`nH�I���Y��$P�@�-����5A��hZ�;�$.�N�53�se�
�C(96����/. gQb3��D�X$������`f!_/�o�A���i�̞���}� #��P?������Հ�YJz��P)�=�
pVo>�s����+�:��9�yhQ;��������Y���w��zuԬL���Q�]�YF��7�6p��tOLh�����k�?o/y/ӄNl�`����DPW��wF�]$u��KzZ��4���$��%�ʈe�S?o��E�#}E�D���$T�h�1l(���>r��_�+p-��V,�Gl�|�eF��wK�$#,�����U>�}�0�4�oH�J����7#�>n@�1V�W}�w��1l����{큕t����R%�+Fu�X2�F[�yғ���,�^�o����D讙�,Gl @.c,v���w���5|��l��ig,�Дm�\bu"QCe��S���kGW;->��ư�J����ζ7�|
��
�����}�(�e�+�$�$�Q�Ғ|�:@I%�Z�a�r� ��z�C�+�BJH:ڠ�s\0IA�nh����#
�2��@�zh{\�c:�]�c�vgQ4i�R)��jObX�Ƕ�"3yH��P_z�u^���-:%�˭j�9�C#r�߽H�B�D�[�7p���[d �%��j��g!���ߐdİ4��x�Ҳmw.��C?���L]$�1�`��j�e�S�"�n���G��u5,��]#�X��n��ON�K�����[Z\<��E�ѳFS �y�lUH)@�S����w���v��=L�SB������F�V�{�
�z�z �φ�WnX�9�l�l�����y��@�^��]�Wj%e�ߛD�Uas?�P���Ө���y/j��9�LP*8F!�C�-��8:/]h-4�̯�k!l��p͵�5�.�Me�nǙ���(7���i��xe��9�+5������N��Ɗ�jv����(?��٣�`���=��S5��1P|M���A��|�d��u�\Ҝ�t B�?�׮3�B���l:(ws,��lI��=��
�DI@��윪�)B�E.�Mx@�Y�mV�0I�VҁUi������?�'�à`���#�v%�����+RuO*h�VL��Ojh����8ĈNj�/|��G�+&��Oc��K������R�d鈫|b���	���hb�~�-_�Ҿ)�3��ڑbB�j��zi@�m��z����kbْMO�� �0��o՞JVR����g�_��0HP�&��Ej��:�����b���|��So&*��͊��E>t��Bn���r�pn�xY�E�-����-&#���x�2���ɇ}����'�OE5�=��t�gjݛnn%�:W��ˁݍ0[r|sI���P+KjW����;��Oh�v��DOJ�JQ{+u� �]�'}�NQ��Q0�DV5����DN���J��
�����/�,�e)ee$)jC�[4�'Q9��k�1;N�F�X���G)ko���:G�]N���eD�$ \7�� ��l��s�ۋ ���ݟk�x[]��n��U�D���[��C�n�S>�c�<�����ԯ�1�h��\f�I?�q�Z��]�����ۄN�e9�5ȣT�p��`���xE����k\�8_lPCj�vDI%/��Y��(P�I5���-��6O�#U��T�w�W��!� [��v����`4Z�7l�y������t��*�O�n�	~j�MK7 W�{C�'��O�GO⒲jԇ�R���'Q�l����ׯ��R|��5v���Y�V�l��9��)��Q�P��+ss�-�<����ry6�s�iC$?d�*g�F�#K{��JTy.Գ��km2�V��l��ww�Y#�Yv�J�R-B��`%�ޤ�o@]A���Ts�n-M
h#�t�[IY�ĉF��J(:٤�[I_3@�]�[�"{s�6�VPv��h:��7؇�ڻ	b��گwy)�Y���^����[��N├����ـ�A4Oʹ^����zԧ�ˑ�"x��0���k��	y�5�Ȟ�z^�`�]�a
�$}��Ut��M�4"$�P��q�#���0��qKJ����k���lks�J�����&n.���-��ٮ20���g�������Ň�2���7z&	�W���0�I&�wZ4�[Tl��n�9�Q[W���I �D��pl&-DD��m^/[�����ZȰ��峎5Y����sZ��8��x��w�\�N�/�k��C�L����P�-♝㆝�Lߛ���ʤ�v	|~�������a&V�Y��/��x�VC�e�UY�|axb#����*���E�~$�%�b�=/b3��_�Q`����2��e�?.����F��v��H�r!J�s��?
zx���۸��Ir�r?*O:�7胛OȪ�M������x�/�R6�+䡻���
�b�s��m��$O��&
�$�U�97f����!d����W��	�ܘ�ƕ�s ���_�-G��#���tw潃Ʉ�+�Б���żO��#�`�4�Z;�]C{�?�3�D�a;� &���<�uQa&�^�z�8ޕr6��^���&2`��l��˜5��)��l�e2� e�m 9�����:\`�/��|���~���і��O��0��vu�����nsO�6���n��F	��oW�*s�&�n��>!����VQ^�b��+f����bx� �;�(�Հ3w�����t�U ���[Uo��;�?½;#zӗ9X��2�D���G�qjj�go>�����-~!�q�é��`a�OA��΂�Z����0�>?)�,J���=z���=��xe��ſ�d���ө��E&��� c��a?��%*l����;�eaS��ne&#��H\*���?D���a h��2���i�Y�Q6{��39�H�r�r^�_9��}�����l0~�2S�{@��~BT�ϒ$Uc���
DM+�¥O�ˇ��o�!�C�����p:��N�����3-A�Z$�QF�W���K�k�#"��m�������y��[���+���w����!�aڌ��@Vb<�s��(89w-ʒ�)��r��:p���<�x�__ �y��Rǒ�-p���h�;�J(0I��P�
deKU��_f�P�mm��r:��E[x��{�L�E|.3Ԑ���B�C^"I�{��S�q�Z�e�R��J�KW��-45�r���h?p����<=�ܴG�%.��H�BqTSFP���6(�p'ɰWY�-2���;�ށ$����vYZ�i �C?3eѓCU�1�d9Н)�����ń�ۜ��6��Һ��!�fr�������Awg ?@M���g�p�Ύ�s�j�C��6b,/��Ec烡��n�g��N�H�جƂl"��h��`p��Qj��717<<{�b�5;!66ޡ�'%@���rQ(LHkX�|0�g�"ϕE���5=%�n��~R�z�`�#�"��?rMR�$}�q4�;���� ĝ�QfcE�ѼFllsPI�W�L>�u��Y��h@
_���x�P_��[��$���Cc�H�9o5N�Ԉ�Mb,��C���*�=ElfcW+pP�}%���ܳ]�pt��H9u���,�,�D��
�2�ro[@��.�Qmj�b#2˫��Ցo�f ��C.G"�>;���NsY�7�S�ԅ��]�j�F��L� Ȳ�Iؽ]�� Y���89����:�5��Z�6ZX1��S+B���F�-����D�5x\�Nd%�/�f��������'�\e�m��D)�ON�޾��zW٥#1�y� |��լ��I�M�.����n�9� �� 6�V��߷�?G�F���u�BU/�֏��ao����>K�*@��f>[F��t�����kh`�g*����������wt��j�����m; �!�1D)+X*�\u�K�.`�
��b4�%]����-�9��d�Ԡ*<޷�n*���A��C�}0�*�&Z�]��Q]
m��Ϛ/T�'d#熿q��g+-�$d17�;8�G����o�.2ʏ�=ƍ��҄g���-�ʷT�z��.aZ�`���:���J���m\�\o�1��6�,W�`S��{G��>��S��r�wTw���{W�@����ŮY��I|I�6UPy�7S��G%c{(H�l#Ή�~l�˛ir�w�X�pw���=�$ړ!o�kj�V�q^#�Q��Hr|�(e��* !����K���q�Č��7Լ�Ej��//�5��g���D&�Z�t:K}*''�h��p����Y��>�S5�ozCi����M"ԧ��������g���Z7�n�)�@=1��}W5	�Җ��rɖ���A��̔:@R��̸�]x=��a�����=��m,��
^qjAf�x(Ih��#��(�,�m�q�0���+�il`�u5'6�rb~r:��,�W�ʡO����_�����+S�$ȝJ��듌q�mzM:�����y7�g:v�����zL�&5���(����il�;C ���K@`�����=�f埨γ�43�zvM�8�z�޲�!L�]/D��N8Ej�(�On���J91���
��;�W��4�aK�|e;MV�G��l��^2n����[����=U��w�ށ`U�ɢo䅦���+����� �}��j����!;h�����ڹm��`���{��J�~X�N�L��  �ے$'
�QV�z�F/��a�;O[;��|E��'.��5�u�w�k��c�*�)�@��%y�L]I ���,>�9��a�}���N0p͎v}�����ўV1}���o�t��̑��$��4����X(�W�R�C��b��cB{t�0�r\�)���˱!,�5��M�p�3����_��0��+F��eoqB�e���5�te�<t�z=����c��	(�7��.�ņi8�A��h{vK�@Sn(���p�������ˏ��hS]%*N4���d��\�#�at�8N8%@G��z)��~��hM0`��{<�x��:��-�T��\�UA��1.�]��3y�o�@�ޜ�~a�nvh�Ћ�$��L�L���9E�����%��O�Q-�:��'�*���������^~�B\w�Fu�D���
�G�+��@��Le�)��C��I�p��s�[�玮,��`z�ke�ܰp�;�pC�`�/�grEjO(r庖>��S[�c�:4��"�xu�~����E2�nJ�-8�Ć���5V�S͋�� .N�w=��$��L�0��)�M1L}c��Www'ʼ����@�SnR��Q)>����=�C�Y!Z`/��"Ǐ��1��B*��0eKR��)'���z.�ّ��8]���h�uM2u<���/��Yf��aX�PЊ���p�.�U�_ow�@�-�)ZA���d�б��,��Ƚ�f��R��'S��#>���р�u�nw:04���Io�rD�;0ʍ���I�����n���>�.�SY'��@�"��%�ʒ����,x�+��b�:d7�X�O�HI{y:���M/��d�ˠiO�
��B�ue���V�e��6!1\9���ER���SL��a�W��C��{˓I����%�֠��7}�Y&��k4>^�#3��S�������������w	ӱ���E��WWc�0տ$�Dt�/=�Ò�_̸��Y�_�����83�څD�@0�m#>�8
\�I��J�p��>��X��ߖ	T՟��z�P+�Q���?V�=��{0E�\���������X�O#��dE��+Im����y�m����	|�����@��l���8�^� 3i���J�{�ϋCU�" �	'h-FV��o<Ki�ɫE�{���s�<�)5�m���a>��'�.���8ν��s*��Y�� $����om���^���ۨ�?3�_�6�zi�7�����R�Ic���y�.f���eo����f$@�n����3��3qUBË6�_ S{m3?�.�+W�d���g2�#}g�S�G�oD��Y�P��3��ᠷ�q�ǥTa�̘�9�A���a$��zB��|�{��e��z����+	�>6M�t���T;O8������L�*��ɚE��ZX�#�a���1��p��ћ(@��iԇ����	<K#�:Ŀ�+���qZ�E�<�k<l�0^�N�'B̔��	S�r��z?('��ףDR�M�����M�.�xTq .Ǭ��ٮ��G1�Kiw���#P2�.�o%V��!�o0�kŐ���`��b�ca2�oj�PI&�3-9���l�s�ƛb�v�g���UI��� ���'�g@s�f0l�Q���\�3�ni� �G�S�z�|Y�����aO�\�kV��h�ps��mWc����J�v���Z�7��d�*�����E�|:�k�SJ��5����v��R��� ��������X���r�UC��D�0e�ɜ���ӓY��q�%ti��"��`@'��� *�񎺇��y�{-�b����*heIڤ�p�W�G+Z��Ơ�y��_�%�>;��QGi[���}(9a)W
�S$(�+�	=d�O����/"'�c]XZ��T�X F
R�2T�D��:d��W��]f��[�THC�<j��L�~N=b��n��Uh@�\7�*?�H��y�p6ZVm�@d���J�_�r,-bWҝ-����2�"���"����zOK|Y+)��8����iQ�"-u+Qq=�2o�F�(�O��_��P!�o��+7Q�LP��)�H�B��<�Z�C*���I	T�AJ�l��Zo�a7�a@A5���	�zQ��s��IDap�8k0�B�
C�b:��n��:`���t�嬆�Q��[7�}�o(ĩ# ��GK ��5���'�QdH�nO���Dzz#{	l�(�;�(�7�����zu�{�m)&R6C�a��|�{M�Uh�N���^{�	���}F2���%�Gʧ��YШx?Ї��Z,zL����A���KvToKY<Fd�� �:���A�b�}����-/�=~2P�b23�R�R�)�����TV.ƃ0��rZ.�x���q�KGK)���+)��]"��7�������oe�@X4��h<wu�/s�r�Q�t�kV����W,�_,�/Dw�W���G�.ϛR��������K�0�e�QyW*�}KK}�}����T�CH*B0����&6#�^P��30`F4'*�Y�d��G��C	�DMH�]s�Q�a�7@VG��Q�k�>P�5��#�U���4�;��A��N���s7~��A7�y*�Jh�<�t�r�$�+����4>�Ծ�S�Y2_Rse�8���X�@����8{�+�M�_�"K��ehq���x��B���X8Z��~ԅe��O��D>2�w�E�i���ʈ~��ѕ�i���˳��Dj��nF�2��e�P� T-��B� #��T��U枭Š�4]�:$f�T���Ӓ�E��Cf(>�?��Q����'���&~������!?�����r��4���\��jzAD���Z4�%��z5�R���sCnȸ#�ͬ׽& ����k�#��1��g�j�1r�?L�\���q�]�YJz�B��|�3퀜�uW�7'%^���W��pc��"�7̟�t⫛8~?_j�A�K�i�W�s(p߾HD���=M��4��RV1t����<�&�v8jg�q%����t�D`�j&yKw���c�ON%�ŷ�%m�*�-�3<�sPu��2A�p�!�CѴn�kM�x
��*1��\�5��a!W��gR6�p�YF Ŕfne���N���w�p��eb��A�{bZ���!eqz���I0�&�'�f��[3OF�^�(���6��o%��������6����[ۄ�o��d?	��M�'�@p�u9���|5X~*
�UI�v	Q5�x�B��廞����C��uur��(�f�m���E)R��8F��IK�����R�TcQ�3��̐g�S���3%q�ϚC>��#6;1=�O/��.A쉃q�D9��K:&�L��*�q�,J��!]pߑ�ydnQ!	�	��	�ث��h��\�Q|I�p�~Z�9Gb'� s���0�Z*�7�n�Ǽ�/��'�ԣ;����82�颫U�|6���[�� ,[_z`cOFS�)��UjѯU��,�m}�dH�QMC�j�3F��U�RGL���m)y�s�i�i������'�'��=v�7�s�������5H��q�e����0A���x�$�+_�z�c�����̊��r��ֳ���֦i.U�@�����&���l�6a@�y�P�T^(������?�Iw�_#9r -�1�;�!hEI�
��,w�6���=�˿gq@���s�5K5|R9��.GK��`V�`�h���"U|��$�:F{�+/��ڷ5��~%]��1ͽ��w�p8�՞4u<�m9s�=>MnO�	�g��xC�\	B��b�i�[��7�Zz��k�1
�20���-j�\�u8'j6Pӗ���qӣP�����=����~9�>u߽	~��6���Ikz,��ǦVg$d��?��{�Ơ���)I!W�����A�6�X�b&$��<�Ts 9�Ʋ��G��dT&y�'��-� ņÄa+|	"��I�s�����Sڀ@yE�����m��9)��	�'� 燺Ú�o�P�<�t��Z����v@�׈��i�i�w:�s�BJ��9Dv�Y��<m=�a2�f�=��G�k3�4���p9uu�b_�S�?:�j�RƝ�_����s�f��uJtm�Fم���e�