��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �	U>��h@��
}c&���`=����nB�&��=��3�&����C�e�4��U�Q3��\�*|��;y���#�՞@4/�6!��	w�A7�).l֬���32#EPڰ}��oS\� �����l{����l��,3���M*�X>`��z*�j,�z����?,i{�wD�>YawĲ���������9�}R�O��8:��*�l\�w��À��AŘ������S�x\��2(�ځx#;��R5�g�)�F�T��[\0.GzM��9���v@���ƣ�l��]=�ƴ�Q��ѽh�]�|=\R`���M�
K��\8�ӑF�Ӳ�{��Q4� H �����M��z/Y(l�/S��y��V,���]g�h��K+cs�CJ�"�+t{5��|y�.��M���3U�@�������Qj�H?��%&��a���?5�o�k�(Z�2�Bv(�N,.F�J�UƜ�����_��u����	��y-��6о�4b$��o�i���6/2O��$�g���t�CC0���H�Yh�
��'od�Ac�\�Eu+��2��TO������k�(���3�7ˆ��:Gn���$�����k��O�z8)U{L�4F��Bxǝ���:s�
��Vnf�����_�����_�l$�վ�F�Ъ^b�]@��MV3�4k�z y�7	%�ə�iň��a؜|v�dՐ�����B���];��x`Vq��e|X�݈�8ZFd�6��0� �g9ޕp��|tգ�!���5h���z�O�i����*l;�P����mn��͒ߎ�P��}���,��d#��;��5��ͧ��"��f[e�	�+�{��l�+V��U��K���TdFS�0����pC1;Z��s��M�
-[��~0D�];�H� ��;��%C$��'{m'S"5��y��Ě/�����mر��	p��-}��'P�ekTGEQ��t�����"�z��)��,�)oY#�D.�����Uf��!6�D_�39�-�Nn�+�'��N�k�C�鲊���SҨ0*�pU�ظ����Z^ģ��ŭ������M��lD� Fx�����G!'M��,�Z�w���4�9u��v�SD1J�@�F�HE/k���t�'`P����� ���T[���W�{{�5eG���VM�j�j�}�#~�����j�3�H]Տ)����4S���v �J���ކ� ��n�Ec��M���=a�Ѽ�;˾�^���
n^Â�� Cwl�����l�X�����7�IūA9���n	��W��/�;�D����qOd�w�� �{���ʢ��qLY�ឬ'<��l��l��ϖɪe���0��4E=r��/+��\�.Jr�n��`�,��7js�Y8��"yRp�?ܑ��NK��Z��~��Ϫ��6[�ӹPH��5o	;��ʍ��:G��5ƅ|�+��Y}M�jj���u��>�Y�vJ�Ȫ=E���,����O^��#_\"c�:?�bL�Z�WV�-<��]+!��*t區o�������y�C�]�9e/����:/�Ë�V'��p��׎O��#��O���g�R�"SV��H�g;J���	�q޺"����K��W�e9�ܰ��7�Щ�B=�`��~_m5�B �x��J�@�S�(jWˈ�g
��ʙ5�"Z�x��[��A�9T�I�Q��4k����r?���@5a�yk��8V�F��2/z�_�H��V��zu�
ܧ�����N���?[�B�����/֮��#���IC�B�HB�v�3��#�A���9�G5����N3�3��E�*R�h#��9aW���>��4�u�-���;䏡�]�U�z���ɼ�mj�b9�܃okXF����Cp4Z3�P��.�z}*O�/��Wc"�3�Զl?�x9o\��V�q�O��@9�/��PR����&%6�S�,0�zm�t`X'N8xvi
�Q�6+b�]����w��v�7R���<���b2����y�L5�(���\km)���Ҳ:�G����٪��m�X7
]�΅vf��T'���*0m*�R���3V�\�57��rR�ȩh|�oxN\*�����ƴvh|���?��0�{��7ю������>�a��ů�f�XU��t_[����\D��MǺ���t����Yw1����W8�ɉ�4<��H��	Q*_�9�`��x\s�L��%��rb�d��06Aj�}�<����>�;K��s��Wu�Κ��^=X�����
r��0��@�C2=�U@�Gi �q��J%o �*����Yh\G�%��ǎkO5����Mf��@����0#.�' � ��ϲ�*��3Y8��
�&��K�k*�q$eE���vHo\5I�SRɌ4{2���/v�=#ϼ��bO2�&�	��T1��8�x�%GB�5�� ���g�J�)����i���E&��?���˵x=@e�?b*���[����3gO[���V�ʷ�}������r�X�b�
�O�y�e�a��CKζ,6��#2��^�;9i��,�3��љ_�0���ژR�2�E�C#�o�J8u��W�xq
]�PV[�~*�X*G�~͖�j/o-���l+�X��YJ~h��Ֆ?��@�`a�kq��&LVo��������2�G1�&��$??Dl�'~*6�Z�vk�*���~g�(�W<@�oQHu۴8���3�K�[��56Ou_y�s~������<+�j �{�I�yZ�#��f
�A弉:�2�.e�[i���,	��:�ӛ ���\~3m�h!�e}�˗�/�3�����1��qZ��vF���A�P)~�g:��v����Y�(Ax.$J�dT9���f���� lR�2-�˦+�����A8�I�*�kn����ߐ��<�EvW�j!~��Ї��� %B��Bf��8�;!�>��u�e�&��E���+��4�i��������u@b���T���X:�n559��<�s���b��s���@i���U)�ɫ�?��ۢ�56>��F_fm�")����4��w?��ҏ�r(N�oC[�'�d���	X��7��SLئ�Ȑ�+�k߬����n�V[�eq�n�(j�-D##���٬R�Ǔ��3@p���";i�1b�#<�)7z�2r��d����۸	��O��^0/2�h�r�n��q8�y5dI�<�2�z�2���KUX��>�W̡��V҈�.�A�+#[�^�O�,�?_A�}�Qק��w��SCfg""h5���SX�_G���*�ew�菢���PN
�i�$Y[Ȍȧ)�U~h�V�7|�w�%�7�V�"F�=��.}b���Y �P=�4���t����%�Oն�ND,�Y$����v��!�tT�[��^ދP�C�g$)l�Z^/����T�x�.�x�#�����8a\&#*�Xb/���Z�\$�&Cǲ���"�F�Ұ��G���	P��}�8�c��m,�W��U/n����e�z�3���O�~��$S��\ی����� ������!ל8wm�p����;4F�f\�<��T�SB��uYP���G
���&�]s�g~Qg�b��oG�@�*���1D�mP*�	ZN��D߬r��V=W��M����j�d� (<�3JV��v�����ˡ�L�B"W���E��r��A�~"u��Cf,��9e�=�h����4���w����E��H���?��g�t	�W�������0�B�T���-���|���sw47��<�O�Ah��҂z�� ��JL�V5�p�`2��^��6�H¢E��l^��7����ﳞH9�f�²�������wiko�<e�_A#��ۿ۔8���0�MY��삎���H�&���4dܕ�\�Iw�*�)�~d�qoEm��Q�������^?�!��?T�6�q�A��c�A	/^���ˆ�`?>*i5-D��8̞�V��ߜK�����3������r�9��̈�e��L��d���-���2��(�6���>�^�`Հ$&��l*g�R:�[6�xDe|�v�tC!q�����=@�OZ����)� �����tN��|x-����A;��a�	����a5����n2�w�p�e�i�!q,|Ʃ�����3H�}��+���#���������rꅠ���Ի@봈5����0�6MO
�UА�CH�IB�=��� (NϦӭ��)���֫�Vk�O.g��l�}Q���`��Q���4P@pO�����8n6H�Ӿ�E�X�F]Y5�Om�6��
��D>/F�m挡mҒX\7��[3������ՙ0�������j&^�Y��T0�`�/�>�cn>AZG�oD �q��޹�8]���r-5�� <^��@̛2���/_N�6���U�2\��X�vL�C��o�0�d��%˗Z��K�ϯ`&���&H�I�n�0_�_;tpK��P�[ά�Ja ˙	���V�$"tϏ���+�M��`��;�'���D����6z�p�ʙ�8I�o+T�ק�D��L�s��ű4V?��ID�!U��DɌ��Wy�n�A��ʂ���v�hb�L�c���v'."w~�[\K����H�t5 ċ�%��g��3FWD�E��\���ӭԤZ��_|/G����?���3&f�rԩ�sGBJ���!������=����?��o��Q�������]�IW|	�[ I`���ا'!3��"9�)� ͼq��$H�_��?+c7���z|���5�P�{ �8A/U
�X�Ɵl[��s>��a�������	��ܼ�*�THڥ= k�W�2�d���Ä"S��313%x�o٤��N���܏(j��گo˷tL�	c��dH/��椞��ǆ�3�Ci��U ��!��u�Sqas
'�%���p�|/3Lv����R�3l��0'dhz��faB/�9o}�v���FZZ\�֬t��;���Zko��^7��zל�V]�ǌ�g��� ��E3O-�	�E�bJl�&�M>H��^�����l������Р�k� )�or�x �y�N�-�]q ���W�� hL��J��$i�%�����9r�R{��ң��@��`u��3T�X�C<��A]P���t�j��#.���l�W�U&v��J:A�o���A��"����Q�7��c��ԥ.�BӜ��9��a+�u2t��&��a0nW/������y�`,:zqU��q���
��OI�g�/3l�
�6#��xV��H��3��i�"�� ��
8�ؓ�����,�2}��ٙ�Ad�"�``Pآ\b�}(A�/��J���j<����"G�jK��η-�P���5/�E���Q���g�@A1?Ъ�8�� ]*ISp�f�0u��|#��� ]�+o{�X�%P����ܙ8���|���.�X�xvb�g��aF��#O\h�z�Zv.�����?@�R&�Q��~�`Ӛ���@[ǎ��J��@�g.V�Xe���a�"b9�C�����#Jh�w��������F�-�����r����[�	�y�6�W��d^�-+%�0�A���ӡQ��Տ��f���I��,NMY��E���������q+�����W�?�rp \n��zBx��Ũs���<���	5�����'�xz��K����f��6�x���J�pE"�k�_׹�H�8K"�M��O�>#2T.�y$<w��}����H��z�%���+���1/��(��Gn��8�ێ-�Eo~�ޢݵ����8↫�&)��X��m�FGdlW��b<�˶�e�v�SJ��#�oZ������T�iŹ$����g�D ���)�� ���^�W���*L�$Dr�*
�����[ ?:D��m�ͅ���? �o=�:�,�%_�	�F-�R�ٱg��uY4�`��
��,�V�󄆥pI��G$#�:������2�����2��D�)_�B���޲�����e�G��oE�QI-�[r�g����3%Sh��㼬�)T���o�����^����3ÓvU6%1����l:|�<��O�ٛ���^*��Y�#:�PҐ���mu�`��$�eT����-��ሩG�i�
���r[��<R��wARH�T��Ο������@�����R�꿢�e������"�Fx�0˾Z�F��hX^�Pgoh���
��|Ξ�j�]�N��L�*{�gM�\�ڭ��oKyO�4=(�p�qWB1w��/��'aY�T�@Mi�p#J����[�<�yE�l��C�O`^�b�4��<��w�$�Pe�P��A�'U����7?$g�}����a�{b�����<��4�7V��;"Y�ڭ֭.��UbS٭�bO��$��f>����r��W3. uO>��7�bD�����?��៫S�0[������������6�A��A���ω9�O�vx2�����<g`�{1��T��ХNe(&�d���o��ǯ�����)�Mi���)�Z8�����k0�m�l~T!�Y�G�8rhq���x#�*L�3c���q�dݏ��`�!����^:M�wЛj��3 ��r�8�IM'�mT��1�z��{K�x�-�#!I�����r=* z�X{/�ѧ����|��F�"��`�)p���KZK�*�W��W�L��T�(bQg��~4HsY�~h�ި�Ӱ��5vmݖ��|�H�;����U�%c��6���bx�r��$7wㄨU����jE�ݗ�m�Ȟ&:�;���! +�/�u���SbN�Z�֋Џ5�2�9r5�iѫ)��س�lv��IA������^;V5��p�b���:�	]�?�s��R&�)��Z>��O�I����7��Mn3X���f( _�iξ�Y����oR���3�W3	H�/�P���b������U�� ���{�v�u�~�_��}SՊ<Dj�;@L��sJ�F�z��
����bgڮԠ
��t�k�2�8����"hfIƜqE�����WWo>�u|!��Z"X��s���*T\��Z�"]��$�c���~"nғ:'Lm�[~��j{���CU��0��A�_��)��M�$��6IĴr�?9@S��v1�A����q �q?M��9�:!���!}�I�c��l$A #�YC�x^C���f&�K�t�3wj�~p�AA�e�����>u���ϭ��
_�?��Ѯ��^l��T@�
M���!P%�\�N��og;O�V�}��f���.maWp��R�_�QXnI� \տ���=M2�y�
�SF[08P쥢��� �$��ɋ\��7#\����B��E�n�~zl#z��b�V�sm[��utN]�D
fQ��}�c�m�i��?W��S�l�A�r�
�)��_P�Ζ�bOux��Z�<b���\ƾ�A��Nk,.����-o�p^��޴��7=X8�-K��	�s�VV��ӷ�w�8�ֵO>O��e���[�}��4܀��v:o�\+a6!k����^���sS���
�����H��t$P�'���Κs��"U�j����D^_��h�<6G�����Q���$'�i�?���z���E���0K0�n�]}m�KL���^`��F���d�}w2À�Uhw��*(M�u��5����Y'�LȠ,�,�̈��� ��{p�[��,j4P���D��x�!e�\��#��OC��"�<[S��_T���C��[:b�	@i�~��"�LV�d�+v���$D>��I|�'T��w���N򗾏�{GHq�w�;�V�{��!L<���d��u��#.{0�U�'�LC�X3rt���X����wxP��	bl��}���^��9@
�s+�P��=���mE�|��0t�r�&��w���o����n.�%��C�ݚf�	��C��S�ȨIs2��8)P�~��'K�%�2d.�*�b1)o���ʂ��W���ͽN郯�X��<��
ϧ<EҔ�!���f���&zJ�w�!!@��5��L;���RQh}��B'�|d�ޔG�w���ѩ�?JG?e��JS?�+�Ccސ�<P��f]��~ܖ/��l�4�Ѻ���~���!ʿ�?$��Γ�|�g�CZԩ��i8�J�*D_�0�ʃ��*��Ȋ��[����(ch��N�&f��q�!C�=Y~-��-���V�{W��n��Vw�yg�����o�ɏ�����yr"m[��ػ={�`��s�p������B"�ؙ�M��P�N��`�^p�=�E�y��Xa�e�WsAgl�����XT|����{�����4x��IlrJG�3i��,Sv�RZ�!����Tld=8��jҩ8ޥ ¯%�D��xCiYR�w����ūOCR48eN25}5�=%��13�cxn�/�*�󊾽��ɿևT��?�x��S>2hd4i����g��׳�ܵ��Vɳ���z���C����7Z��ч�hx�0%a���(�[��9;X��7A~�����̗8т�9T��-�����1Kb�	ܻ�_���%��m�H�[�?��ZD��dխ&^M�� �[hq5��w(�R��i���m���o��Ş�HssR�׻Fd��S���8	w7)�
s���M`&��ԁ�Ć�!w��6����
-�D���6�p����epT]p�����B���4��}�����V�;�B��d���X�;�2�$�n)g� �0����7�}���bo�O�F��O����mF�8Ҵ�T>ů�[�fK�e�K�i��HT_��4�@���j��V��~����\{ϗц^�+�`q�������'C*0�v	m4�G�Uq.8�.��:�A����шr�W�D}jK��]�h�FJ�ȉ3�M�TK�	���J�OA�ݚ|��SD�� �3�&FN�l�Cqf�U��n.'�� ��'�MVЬڔ�,�9��Z��YfT	�)�.��K�ZZܔ@�m����J�?�B9�sLC"�������^9���TS����1[��6���L���]��0�Ij��b���V}����jc,��Q��B;��o�(g9��\�|�nW�U�,89zRz�|d��&5���v��Åը�.��C�N�9~�+�.Y:!���>��\E����T�"�T�l�
����S��r�3^0ݒ��m&QG�3↠�$A��S�����[��Cz
ݍ~���*:ar��4���z~�:6?-x'��'�*f�Ut-����	�bXr3�]c6��6'�Jw����)�����ߎ�Қ9J �TYMV����)�~O7�d��Y{�A?���L��|�l�um��|���{�
��R�ćo�亊dp�2z��oeί�B-��e���]_�+#z�w��"*B&`;/�`ߛ.��i���v�c�q_����?T�ăC����*sz��2us� _7�ze�kEI���8S	yå��v�q�|�V�WF����)M��Yx�$�4�u�ʣ��}M����ô��Pz���^#����~���`���u=��	oְr�:Y����ᅊɀ@���&<�_x�"ĔI+�vƘ��E��趰�1��ze�Y����a�cQr�Fu�y��4�����
͕~�Bn����r���@��V���T �*P/G\嵽x��{�$iV�-9��9�yEg�;_�����_�FL�l��b��d[�(=�\���eNIGV2�M���H-q�"?�f\vP?�~��CQSu=�$o��*��jX�t�$�}�u�K����=
Wg��=1*+����¢�Z�D}�܂����(���B󌛳��~�}�}��(�ex���BԄӂ��0�a.8_�A�.��ef0�L����?���S0CBm��z����Ɖ�n*������8P�Ȣ߯9h��L6|�x~��t[����/A�>���V��w��sLo�H��#9�����2�.4�E� ���@���0n�S��LB
�h~�y�zq@�T?�ElE����Y���GRm|�*�i�uQk@7Mƻ�IڋN.!�i{��Q� ��M�(̌"���i�*�Ŝ�7�ݵJg	�!�Y[w�I�;KILk.T�F��kR�2�]f���M
�fI��\$J��48i@�|�x�TK�ٹE��F:�xȞе�����}�K3�y��M�2��^�SE���W>��"��"���������PA�%F��Ijf`���,J x#&_a�V_��RK����M9�`W6�` � �At��^:JF�K)ηE��jhW٬�P\��䙀(�;��e�)�ޚK�x�`���u�m�d�u�IO	��[�0=��⺝��j��B O��s6Ql�X�'%�I���V��ED��.��|���?&���f��hlo�� �4�;�w_��������iQ�o��ۍ�|���D���E��Ƴ"�ɛ*�f�SX~$'r�o�x/i��;n�~J��7����Z����+��|Yz�j���]����hH��P��6���wbu��ޓ��m�h!�G�����2 �bF���� O�D�#k�xʘ�`yE��J�im\E��u^�KO8�i�t�&r�����%�ap� l).�5��Ìj)���a3�/�r+^�l��:J��cd�hLa:���z�R������[v�B�u�z"��f��H�I?� 	�mWZ�܏E�
rZ�(�qe
"tcl��J^�i�Β{�"����/0��ؑ�?)�B6����gi��b�,�O2�e_���ȵ�V��S�< 1�����ɚl{W	w�#�&�y�H�2K�h�d:Z)iot�~�w���D-C]�UC�=�'���6�s���@ʷ>b
I��j�~�m�)�����UK~�E냻r��@�%��iK��^5�0�=I�zC/\�e�}T�$�3�t۫{8��n��~�F����?᲎	�ׯ,����3��)�.o��t�L���+wA,Ǫ�\Tcr��#Eׄ�G�
�eMJ�1��&awD��%�"���W6��F������Wk��Xo�=owk�x�@K�@\��GG
�'��j�:�Ň�&����Z*{(@�E�:\���/-"KWjRug\ݰ
�j�l�{��ص�����Th��B��@�BJ0�{~�k��R�i�Vb��*\�"�3f�9n�]�T�;0�7*(b�6�:s�J����`�4"k^�Dgv�1&�����c�C4�v �7A�A��a� �*^P�.Usa{#yl˱9-;��2!�u�,g��zu�Bvw�����&ʠ��v�E9SjB��� S���|�?��:�L�~����QO|��E�";~E@�.U������E 
�����lG9�XpH�ţ�B�h:�d�(���y�h�n�9u��@�I�_~���źa<��8�U¬�I�b�������P��
�3 ��g�hd���L�l�`.TaA� �%��
�"���^,]�+-���f.ּ�����X�Q��&����;.Z�w�VI��æ�[�00�v����PW��եu�#�N��_y��a%��2�l�>���aũ�V6x�����JԞeu���NE�Xs���óT	�J�Eu��lM���e�X_t��*V�q��q�t��u[�&�G0ߢF3�9b�q{1S�"���<��*����ғu7\C�
�7|rC�=�)���?���5�3��N�#���1�����єͽg�U�a����>:!�x�a<��HP�7i��k���v�M��d��c����
X�	��(����7�G�2�d[�qn�2����ʣ�?���Y�����&@�,j�G���<��I�<n�������b�5t�|������aJ�vò��O��W^��\�f]4����:�;Ŷ�\(���Y,RW@l��I���I����������9���
���yYHޠ���8	N�C�{�����C���������w�H��L��^�k�S�M�KoM7�_}W6���HCN��i�͟���u�ގ�ԉ��$76�妤ŋ;L�>��S��e��L]o�q�gi�K*)N/v�ě�P�r�#X|���z��u�C�6�_������Xմ���2-oZ����勾S�����`���T�A�Ϊ'7��amї��꾇L{̘`ο�R9~X����#��/J�Q��Ma�8�-�Ћ w.HC���'��|z����O�h�S�?�T�5���D&g�;�>����׀�1��z�!�m�X�g�@@�wW����O���ʵ���E!n�3pZ!}JL�1&&�PE����+A�:��v�������e�bO>���a� ���������9B�4�9�T�2�p/a(f�m�a�%!ɭ30����s��"j�.a��p�8`��t�/h�qf�?�,��]���m�%gh�^1����~ N�u�$��#���,�#��+ϖ�n���V�Mh������5`�Ii�:��
����<KC���$u���i^�DN�<�g3��;���0kMoF&M75��bz�x�$���6~�;�%,��)ג�SO����Z���/��}���[)4`f�Ѧ��cbl;%��1�����>:�)��T-ܤG�T�G\R��1��剽��(���Gx�G\A��x&A�P��+bv{	Um������?�,��j|>Z���p
�ӵ�F�j��f��ldܗ|8$mׇ=d~b?\T��GԤ��~U��J#���_K�]�\ �G1a�;���%&͙>�&��[6`�6�M��&V��ġ�x�B�KF)�D{c��-i+�!&e�8@L����	2���M�υ>Yù��� ����(�㬮*Y�H�_ EgX�E�س��g��lnmbEZ[mʱN��5��1~�`UO�)#�"�s��|Z�@u7��މ��y�M��7^+�	n/Y��%wj�KlAcC@��0��|����o�d�c���J�_D
�i?&��f5,����{�8�l�(Dk�Ԝ�xg����-�Ne���Ot�͉�c-���
����*j�<����?M��$ߥL$��݌ĩ�Sh� �!�ր��S�x��N7%��Vl�A��j	ח�½����Ǚp�Sv�u��0���<�ʴ�XH"��dm�_��h���^��R�.Ub%�X���:1.u���rA���lS�Ǫ�v͜?�
��+ɱ����<���>�� ��z��S��P�eP��o�F)�4�]}B�Չ������fy�p��3�x]�#�����sb��:MI�FS���1i{���<� ��#F~lK�u粡7�ɮF�z#q�C�j���?�X�0X�vj`�����>�����J,���%��՘<�"(ξ�W�UR�n5�[��Ϥ�5����/s�.�>�	�r����	?~&~�
��D}�^��絿������u�#2��S�v�-A�
�2��n���I��}�:79�o2`̪ˉrn)� �Q*������ڍ��_�*��"��V�&�\L��S���s,	s�2�I�s�q�!˙�{�e-�1]W:5o�D�^m&��>|{��9V>NYvB�㥼��*|`_d�>kZّ���Z;�Vٰ�0mO)}��J{ZUQw��o|��o;�Ί�����A:�,�_k�!��|���]��Խx��X���T5ŷ��� ���:D��
"Vߢ�z ��{Qɛ���o
�3��Ij���@�m��&g7,�Re�i��K�x����.*����f�1���N]� ~8�D�^���.;:X�<��X��2T2��b��0�H�$�>t@y���= ܃�O2S`�������@���ݣ�]>m�k�=����<�+
~���-=kCm�]��v�0�P��C�
tLMԦ���z�2��a9m��l��A����(����"ή*�k/��'
CU`�����m���6��A7�o�5�N�mq?xx�q��I,����� i�-v����1/V�n$2�pbĵ�u��,j���ć�=뻯c���/bgԛ���cn�:��f;֊����d�t�P�f���-%�8���R4�����f7��Z��
��,O�k<������	�1�A��c&D��R�g�����8����N��Y�p���s*(Ta���
�;����	jI�e�i�tT�&A0�l4l�����PV�ۄ{6�T|!d��#]�OTɟ|Ztv�4 �)���ɟ=8���u�oJ=&P���f�Fgl��VZR�d�]bq�5�^�I���-�M��Yf��?̀>xa&�A��%����'�&����K=q#zy�=�C(��ns��nc>�^��{_mv����{KS�Ba�(%��5ź�~�<&l��nho�Ԏ�F�v����~�
�mL+]��+�*����f��H��sqZg(���)v��	�Quێ�����K�`^:�A�U
���ܼA�|�����pv4���̝���d�Y��<t����5OJ�=Ua���!5@4���d	T}�0�L�<a/�B�hP"�u�*��1��5���O��`���$����{��}TĹV��q���wF�`z��I�w!����1I#M���´٦�I#�7�M"lS�H�x�/��#�&+����'p��:���#�f��U��atn�"p��%9�ռT��Zt 
�00w�>��YK�\���HjY���_Q[˽��~�i7#W1���/��/�\�#�&H�q��R�&�}�WO��`�����\L��X��hu�����4dfu���rfԩ�嫦tn? M�ш�1�M���M�S��%,�̨�v��Bt�'0��V�������	�	���)`���*��eA��4���>����4t)���m��o�iP���WU���R�,D�l�q:�uO;
�ʄt�<`yq���}UŦ�N(݁u�31�m�|�v͆s�I]�O*�J�u�b,ْnuT`�7,K�l0$�)�+��
��>>����	'+�T�t�D�&6�������1_�'��|��G��"�Wq`ra%ػ� �����%r��fN�K�F*���H0��W~�2u�8���fE��f�7����e�����O\S��4']�9M�l�7-�5��,��{�ԋ|�ڏ������{��x�֟�
d��1T�����$-&�.K���4�Q,�����~��0��a��\��8�a%⅖/�`��.xU!$�.�$,1::�Od�Y�paK0p&�ɸ������4
W �x; ��qE�[�M��C{.��/m�~�)�Kv��T~���}l��?��:�hL͙�J�	݂�������0��3���e��#����,��i^`����q/|�� ��QP���{N��6G`!���(z�:@���G���e�J}��U�
���\iO�è?�N4��K�N�/mԸ��D��� Ł�`XR�L`,�U~�{��<]��H@�"s�_R��	[�_l��K�ؠT[j����Q8���\�8g��w�j�V�����Ilf"<�kp^��.�g'����ˑ���C���V��$��|0����'u%r�h���,��%
�0�~�y�+��d@���x�Pk�0�/���a!�p(RF�k�M{T$�aP�<�b���@*Џ������&:��8��YICξR��,�TX�����r*-��d_aL8�&
l�x�f'=Gi��Qaך�����	i0�8��Bw(e0`�+lZ�����Rtu����"�W�q(�&XB�hNϏ�֬Z��?��j:���1nҥ7%��8�/��q�� @��,�ФGqx+�;3~O_��dw]X
�^��׌Yt������Fq?�P$?ڛ"���J�[�����������k�n�)���s��[�[N�җy�CφM�q
X��Σ�8��pbGB�4�j޻��! p����hS"��g[7%5�Gw���~͎b��H��xY�������^~�~\!�L�ݞ3������Q����[2�GtZ�|���������CI@���zglOՙ�6��N�o3�)��� cvE�m��ϣ\"��e���F�h�J	y��R��dH.n���"�Ϸ8�˫N@dIy4����XY�L��o���-�%1ɰN��.���)̗�Woc�nkf�e��7�wH�����ԥ��Π:�.���ߴEP�'�0[�d ��:E[���Ę�x��wRM�r���T`��k�~ϪWSH�{{@�NB�X'��M�P�~�a� �H�2�_�>#�Jyxz�W����	�6�#�j6׮�s͕�'rٞ�,!d��'1f��F�D�*~�+S�S��P����-}u)0C�T���FT��/^�!�и��8��<;MB��� 7Rh|��Ȇh@`�2F��Y����e͎�Qњ�"�ʌO\�i��X��uU0|�<DκБ󚿂1��7[o��e��],ŉ��G1.��8�p9�J8�DH��s��f���uwa8����?�Q� @�∺��|�T�8�\	���^![:Qn����Ϯ'P���f�2��A�ߡ�e��j�^ۃ�~��v����-�����x�K_�\�ߌ��d7[�1{�Č��.V���C�L�~������	%wi�D�W�P�I��T�2�ܕ���Ri>���T��=l�,�C�A<�����ҽ�̉�MZ�L�P��YI���`��D���::�/v���j4�����e�.�Q߿h:�Z.�%���Q���������%���ҝ�P�Ǥ�ed�3*��R8d��<��q!�4����:��aFU�gVs��=AE;��&�*�h.@hQ�Y�h�?4�@��x_bv4�p�o���A�Z{�����-�,��N3⻺����84� ��X�� �W�$�$.vBO��=E�׹��oL;�L�}�`E����@|?��C���nY����Ezk~,�"͗��c��߲�#b��<��4����W��QA�v����p�`U�9�w�B�S��I�v�_�-t2��;�[RΨ�p%R��&]��M�y:°���+�n�>��ݖ k�Y�H��T�.gVÕ]�c��1��~y���`�7��]@��}:g:7Ì�u!�\j�q��3�8T"��()��>�T[�bx3D>�'g���iKQ3�ˁ�A��q���;�HB�&�,	�j���Bo��Qu�ORp���Nߣ�X�	�35M�WR�o��?Zߊ�)D�X�fqk���9S����*���`(k���%�|�ioLQRr��$X��|�.��t�*�A"T�@�RBC�ˊ+�bd����I�+�֨�v�v���eF���uz��5�r�����m��3��M����M\�BP�e�`�`�w��9R@�������'��D</�ڇy}����kt4�X��3DV�jߦY�Sg�d?F�X�� Ђ�5���i>ls�����I���q�t9��b�L�wd�4}�	��@\�M%���#O�6ř����Ѳ�z�GS.�i�6�* ����^�hߎ;��N�@n���Z�	�?Z*��N9���-<�6eA­{3X�c��+�r��o��~~�J-$��Q�J�ۂ���?f!"��Ef��j��YS��J�O������~t�9u��d��9�a���m�U`��R�Uo�R����6��V���kɉ�R��Ų�P�#ES�J�����_�K>Ojni����O�����!�Z<N�e�ma[�̩�[�B�M�~6
\`A�<��M�� D_Ek�<B�R��n4������m�����W�~n�-�l&��q��٨Y��/	���0�(R��K��=aݠ}�Q��4�5`:�����dZ$D"�r]�p��H�`<X����iP��Lc���xpՙ^�?k�S #?�#�����(pю�>�S���n�,�?-�F�ϕ;��\��A��P#Ҽ�ܛ�PHi���=k�D�Щ}��`Q�D-	.-�x)���TX
J�uК�_��I�Rj�݃����;�����n��Yg���׼��S���^_�Α���ǆ���8���k9�A��R{�.���g��꟫X��1��Ո�F��(7z!��1��0?��@ޖ�v�qG�n�hS�	@��s�m��>�7oF�]Sn9��Zb��x�x��Y����zo,�=يZ�n	�����v��Њ�2?����Dq鹴��q�!q����[l��\hnLlX��]j}�]a�\�L췇;�aw�k��;������[�n�T���+_d	�'�؟�����(��dG��@�U���X���P�ς�Pl�@��e��aBqHWͷy>Q��Hk~.������i�)�C����>`x���L�
�������\��'�M\��P��"�ŧ��*.N�z�Z9�-/'�[�t_�6�\t��|��m&S���9aX&;(]/��|��9��q�6[�MA.@h�:ft�}8D$��$hT�߿$�U�N�*a1Q��^K�|�w��*��J�1�����)�c�m���-�:AI�1r�Tq[~��g�"/�x�ک��.M��\��zN��������zQ����2�{�_	[ϐ�Wx?��l�҂�!���q;ֻצ��i�7�,O��f�>�An=��q�_��殮����ଭ�Yz�m��//���L)�c��˗Hi��h�u�����և��i�����Q,V���4t�[a
���<�K�]RkF-��݉zF����� ��E;��������8������I�ؙorpF��`�~ii�~�M|HJ���ˠ=d�z�Ѹ�U$2���x�)'Cm����po�OӺ�@}y1J����Ћ�AB��>}Q�����rʆ.�M59�0�Z&pc� �#pbB�|
�0F��f�;��~2U���wmp�R"���{�U�[���k=�=eUI,�7�#��WK� M�ȼ�����9��Q��6N<�����}��u�!��L	XD'X��/���am���#�A`C�z��s
.ۜy������.��~Dk��2��{��:&?˜����>�蘸wz�-���d�L>����c�'f�8ic��:��)x��e2�@-p��:q�v�̴����fA�R�{Ӕ�4w[K�R�~����<!�f�_r��W��i����Pz6[`�be�&���,k��/?g�Μ˂���sx�,��~-ա�r L� t���2���U��?�XNQ�J��sp�R{v݋L�l)�&�xv=�ۥ�V~�YG���(�BB ��`�|������Q����<~v��
D-D b�.���=+t��*DH2�z��1�qP{�I�A�`�������6U²��U�*���}�-�������W�upa� Ь �=��Y��srُ��H����s����j|�����-a�F_7_��9Y�%2�Q*�ׂ�����d��uf�Xh�����4;I�=��S�ǭ�6O���zH=���׈��-<Y����"&���˝�7�m�7,�OIƂ=��2dE��B�|"�H�+�y`;�uox,�f!��u�[ �%��[ v#w0����܃�|�7e7r-<���2_o>7ݾF�	f	;*32M��m���+p��ʼ��]U~�9�u(R�au��� ���FwB���/�͘�=o�;��հ���� �w0/��F�GAL�=O�k
O��[�{ƥ�'�v�����cvu���[e��}M}�u䃥��G��xA���������d"�N��VIuQ������l;ғ��h�/̈��:���zV}�	.V�4��/�	��n�B�-����-�E)"z���V.��pt�,X-��
2z�@����[�c����&)��54��t�C=X�'�`%m"B�n�Tc�F��<fʢi��� G���6~4���1b�/d?F��~R��Գ���v-$�:L����v,�(���~��=��ݛ.Lh(fۥ���R#�c5�v�Mu�Y�a�6�8�Lw+����+�?F����ۿѷL�Œ$L���]�A��"�R� ���}v�*�0#l��7���h����fr��N �\z�G&�dI��i��:���%��JA�`*#�) �yҷ�_�0����c���= 
ǵ^�ՊEc�X�Y}�	Fey`��+�� �7C��5u)2K��ne��}� m(�6���s�ec�Y�E�0RDi�8���_�����ɨw1zI���TO:f���;�d|�
��K� MN�4ZK|����K��K{�L�Btc�a��1�S)M֞�2Eb�:e~� �ݥj)�J��$�i�ϱ�B��q�8�4����u�\N:��u�q3�~�,%�֕~���,�SR�T���2c��s׬�c\oo<Z�y�$��1/&I� ,8�?'�
'���T#��!ٌa�=6ޜ��;Μ����`3�*S1o�3ji��8mT�t6;&�a}ڙ��:��pB�GgWǗ��	�/��Ҥ6�bk�9��؃��<�v��sC�H�_uD������vb��3�h:�X�%I�-����}R�o�F �P�Da2O�CJu��l0DL\�:P�}&Ȕ]��'?�*'�����h�wt�aggq�8��)M�z�f)��?d��}I��JM�剼��07�;P2��U�M���LV�BTz�F�A������Լ�� ��%�Vug>�����}����F�lR�U�BiAM<ī>���j��K'�t���S��I�'C-I[���VΜ�����@&.����r�m��s~�é[�%�ZV���0��`c>z=�����H�����HU+��)�QY�-?�-)z!�LZ��ݩ8V�6�F�g�3�gcm�sm�Q���jj���S��+�4�	��҆^C��"��eQ�R�W4�~�ڂ����!2����"!��?^HDQ���ZQJ�0PbӿUe�� 6o��>(v�?0r����ј@�#�~�M�|1�)����$+?�8:Nt��q ��!�*�#�6'V�_nKޜI�l'x���m�|}�O���͕:~���9M&�A�c�$��n�U�g]�{gWr�a^��q���Bj�Q���ߜHX1Ϊ?�m�yŉ%��@���`�±B����G�R��
ΟV�:���M|��T�i�9���Cɜ�s�I����k�-/��h��� >ԫ!�+9i�E�^������*^u4������J�[TW����ׂ���l����,ck3K�ў�N�h� v۲y�O��Hm��4ܐ�%�D��ٻ�tr��x��{'8����v�9sE�I�@�g�]X~���ר�-vV�
��]����dе��Gp[�0��u�3ɜ�u�9�[2���}���wϩ�_�Ap�H�ӹ�4,���q�O�9J׮��r񽗔¼t���� �	���!I[���]=�*-��N�V
�)�v����F�u�@�b.>�C�KdaF�,�L����\��Zqس|��GU���ƞ/��n��i�>?�����+�5K�CG��i?�4�i��T�XE}L[O1���>��fi��v�쒟pd���^f�w�/�rpUht'�H���r	T^�u9/���: SDǀ����N�$�V%�SX�CA0p���6�c���F�$-`���5�}�@*�vSN#�N��2��B
�ڛecV�r2�=�x��9��bb�$�_��H6�.��R=Y3��j"�ؖ&7W�G��r4J!��bBr �i�펩�7:&�B���[U�$A�b� a���C���r��5��f��G ;�Pubަ�ϊ����Wp0P��~�^��@�z@{�O��[7-`��C$)#!A��|�pM�Ζ#܄>n�^��o��l�BZ ��-�c�T���rԔQ�6З'�#�z$نdh���"X�qw�����P�c$�����<�8@YE��UM:��q �+9��:x��1P��&_�Tq�buިѪqv��\0��_8���+��#���ҫ_���E�Nk�٤�0�i��{�5���\|v�ה<1��.��~�U��t�H���;mi�	����ɴ��oo�W���/L�J�Q��'�F�YѮ��A�"N�\�'��}#�;���嚮� �jlzt��>�U�^����5�����پ.�zo&�[����'}N�Y���Q_�o���@�NAoq9�Ne�����_�`��Vf��Z�b[��t�) � 6�P `���i�E�i��/���Rgx�:1N"R�����MI��ϟ1�8�����ZU#�Շ�V��x�����q���ں����0?/Bx�H� �`3�sn�{q���ٯtSŏ$� �@.<�R_ң)kT�?��	�p���l�պ�����S��}狪ᵉ��>�S^�':��D42-��4l=q]���9�נ��|�#�9d�/}3���k�b )H��g�$c)L��[֞�1�Ѵ�m*ZJm**^��V�d���W�� �)������[?�x��Ka/m��AtD�����P'A�v�|q�(��k!=�����3=9MJB��bb�;���<���c���V����?