��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�g�����B9>z���SEޱ\��c�)�P٨V�LB^���l �g��V�P�U���,Dc�ך�9���}8$/��w'ڵ�=e}�h)��8�E�j����h��B�&P&rV�� ꊔ�3�4���Jb���at�$�Vk�tt�r��j���'�4	<_���s�I�H���E��A3���^�.�1h;�TmYS�������@��_=���y�@IA��嗱O��v8@�d��l�.	Xe�*���p���/�z�e��bs���A��{�Qމ&)l�8Q<�%V�����4/f�Xow0X�����*�d� ���o�l7�}/���n`+v�ή��}�*� �Aw
cW��w������婢L �\
ң��0a|:>��6�ۿO�4p�7*�#	ʪ`���̢��-�<�L/pl_�(�Ꙙ�_!)�V�e �����<
�#�A���.���|V���]�B*ִ���E�ǘ��%5��-�d� ��9�9���9��E<���wƄ��Vc��Ԏ�#�z�
P�1k�C�0L��E�S��˜�����F�O��&�$�SJ��w�.H�*m��t��D�,^��m�[e�<k��Y�LZH%\����)��o�,��<��z1��IN#�k�q�-
�5��=�b"pK�����>GV��&�F�t	��C'V����ؓxYBu0��|4�fV����c�^ಷN'���5�}ƃ'_)k��������7,	�k�ՠI��?�:E,y���h����2�~
J7�8\���2�~R�J��`��Gnl�n5`�s����1�o`M�%��y�#ZN�)iV�i���f1��!tv���U�I�|6��_5C6��")!1^���qĲ����m�f�r�@f���!;��~����ս�~@����#]�����U�k9M�(�r�y���Qa�����Q��е�b��X+(�$�ebm�"�5P���+��|�ū{�(�;/\%��s�&�f#V@K�#9ZX�C��>���X��-�=Rk[2q��k�V�Os&���Є���t�� ���w`\Pa<ኪ�������|�myT���׶C�}Ŧ�*�4��L>�����B	=pO<���$"}$}�Jf�fL��<��m��-oNkA�0���j�}d���W���r;C�+M�����2���֨�!Up �0j�b��J}�84(�/����k!^ڻ؃�F���{>x�*nJX/�*֣�D��̀-i���D�q���st�´�{�Ѓz�(S̇E[��P;�߮�h�a-�o˝��6W>Ü�/�[����)�����
�U%��/��U�22�P=ky2�:i�ջ1w.ne�V�F&m���Ɣ���3}�ڃ�y�J��� �R���&m��<oSiQ�h
�D�:0��ٰ��	�X~ ������%��'��6����7�ł�����V��70��9�����K��C����_l�{�;���[\����ܼj�EC<�� �q�-��E��@�����]e��E��n����%J��~�W��\�jV"����q�O1B/ƻ�0K{���K�ޜK�8�ZX�4���=�E
�z��P���lC��E�RoC�7N�[�h4�f�Q]�W�A<��ƗsK���6\��F��)�ԁ���M�M���v��Ar�F�b�&��ڔ>�T�z�_#�gL0�1!:��6(G7����w�$�V"t������.kv+�6I���?���[��U)�V�Ī�J�U�@�0Z$גT��lEј^��TO5������_~tX�1?�{6Z�KL}ig����WK�w�8ouY�^+�� �?Z9���m�o���������7�Ϥ�U�O&��rW��9e�f�k����Uw�#P���N��:o7��M�z%�����W+��NB]k�C��7﯉�ݲ`
���y�y��[��X%�-9������	h�g���N�6������UW\E�N����o&d�Kdʥ�M�P�v:��v�����^�6Z��,�ԡ�eLL#�Ş�4(�q�
�@�q<��P�h�	eA�8sȔ^�v޼�MU��
��l-����ӵ��� P��dј��y�E�p�4_XO.�C�Tm�?Sؑ����%�ȫ��?b��Tt%��7�2�}o]���s�i+���ŏc�#Ɇ�=dٵFiW
}$��p�����i4a�\���2�ûŉ�X/�1 �I��?V5�"�)o���Jy�V'���$�����&p����	+�uj��F��F6�p�p(��:4r�C�0�Ek�\�L@�������=PV���b�o@�C�*ir�S�0���	�1���e�b8�nQ�-�b�%Ѡ�L���U͋�����5���Q�.������L�X>�Zc,�b+��#�����q������Ú.��α��-����$2���=��)73+&!�(��el�a�.C�P�czó�"��<-�,��3���7:W�����.�2y���:���w�)�m�%��0:;��[�S���T�%��6��/�a�B$$�6qDj��(��X�j�_[��`%^���9Le��	��79t��W�
_��l��c�(E��]���]�r���~�E��!�K�����|f�5mD��ȁ	_�ĭ>�W ����p��]���o8X?<̝��p%��B\�c��N_��
_��� �'��ン׻����9�^"~n�mY��d��*v#�Ŋ0<�7a\���-}p��t�^g�� ӟAbٽ�7�� ��љ�O�)�m[���<W~���p�1�l.�>b��	�	�ʱ�
#F��h�q2�������YpkZ�+�_��58��?C�)��8�)�5�9��� ��fѲ?�+K5H�`{if
����@��(�[-:9J5��^p)y�vf���s���l�(+��y��r*��1�((�۱�ΕT����x@l>���?(O��Q���Ue�W�=)�.xTq���ƫTk;��-σt����{d��y��f8~���ɏl�".����U�G����<���0+�Z�}
�!}��T�q��V���s��N�ր� |6i������b��c��6[ʹ���:��aԶ�͟��U�>��hP�q}�1��� `w�RF��q����sK��\g~�˿�/��EMű����;�%HEd6�����6j+$m�q�2��n��[%CFv��ޘ/��L2nF���{���Yg���i_��4�ԛ%�5K�S�v��5m�8����s�'0&:-:�z!8��"q/z��Ӝ*�Ѣ��v���#�r�*��0�W��Q��k{V�p�8�h��F�C}씔ϖ�E-gy �l|[��