library verilog;
use verilog.vl_types.all;
entity flog_altfp_log_csa_0nc is
    port(
        dataa           : in     vl_logic_vector(7 downto 0);
        datab           : in     vl_logic_vector(7 downto 0);
        result          : out    vl_logic_vector(7 downto 0)
    );
end flog_altfp_log_csa_0nc;
