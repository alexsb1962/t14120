��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�������+C��̐����ѹ�b|���o�ud�&I�z �]�LE�wgn�8�F�(�˕f6�O�� v��"la������#8��Y5�O�a�����������$R�	#��p��MB��
]����|�" �n��:���}����ڤ�����*���g�{d�d����"?�pɷ�YTE���F���K~ػ$К�������Yډ�l��=Vn��dh��A�J��T}�<O��ll�.)�]��߫�+ڢ�[���]g��e&	����h�5ȸ�:4b
v(���D���>�=�0%�:>��2&T����Jq*�!����#������0dS\��ςT8�i�[��w
�R�l��!ă���I���^p����< ��~q>���0�6V_`"?����yV�)�a�H��k�F��I����d;�G�����q]���PE,B��r�I�/�{yD�=1�î�y��]�ZrL�<vR�4�������ϲl�0�5�fQ�Т��e�W����/x5�hu1Vl��ɖT/����XL�s��!��ct��x5���@�U�:!YJ��ę�j~��).�z��6ѧ�w8���!�j}0op	A��/�kfD���F�l^�𧅤M��q2��n��w�W:k��R>O�b��J��6�F���u����s�S�Dsm�P*GOp_W6=	P��r����*�||T�r���ށ�%�j֩���F�R��	���e��3t��!�"}��hN�<��Q��0�9��y��/:��1kn�!���zD�wp;�����`����6V�k��� �fŌ��jß��	����jL\\��76wf�:��L�d'�x[�x����W�Fb�w��Sȯ������Jѭ��(�����^L�j��)'��e�N�Mќ�7��f��/�r��RӐzP�E����|��Aq���uX,�T���1`��A"�@�����9�kh�3+=2�<aC�Pe�=f�jpQ�pk�C��e���H���|f~�ٰ�x5V��g-�k�\��8N�e%����#�Vq4��)� �yiF�ܕ9��L�e
��T���n����� ���6g�C �i�����$� %��~��u���d����*ҿ ܍�|��� {�R�����'�����S�P�dy!�w������Li�^޼&�E&���5��ι�|O}�J�c<nrA�D�ϰo1����DA��gRِ/�yi�N�~��H�	됥+z!�{�E!+g؆�d���C����ß$�	>ŭ(�w��Q��������g��A����B�!�O����6��9��h���2j9�\A�(����=���W$]��]|=Ù~�!l���)��N��1)����>�g��Kr��%���'/i�׷�~�alz�@��=��V �^!JffG��IM	N>:9�F�#�oY8y�pY��\S��_�Y^{\yl�P��As�T-��3�JN��?k[y#�3�=D��%����tt����p<�E�����m��;l�VM��4��;wb���*����/)ݰ���/?!k�1��e�-�j��ԣ��D[;"S$k�>��aV���젆& F_pA�Qk2);�O]f�V.�%��d*4�, ��]_X�[�4��u�\�ʥ����aN�`^iߗ )DdF�qO����p獞���=�	5j{8�f�ߔ�Mҗszw�#yq<�M�ܐ�A�P�1W�afmc�x��Ø��4,INAB8�=Rg���g-������ZS˖��^��By-��RjڐsApQ�X��!�G�A;Ý�T��e�*�V����ȁ���b�-�}>� 8�kx(I��?��������

�3�K��v5O���������M-��KO��;�Ga�ft0C�
��U�@�}%~�7��J�J��e��C���G#wA�^�tF�X��\��M��]�G�SE҄f�o?���~qI�`����SY�b�~;S:8 �XCu�9�5��8~�6�W����Q��Nbm�j�Ia�"sW,�	ƞ�CR�Y=o��%���&}�ݧ�i����LGPV�j��A��Nϻ1K7bmLw[�r��6R���UI�m�4��L-�Q�'�~JBο��j�`���0��AR��x��i�Px4�͐x��2J1�h��[A��$�l����W��9E��o������e"x\��B
:%0 �C5fD�=G�.�eq�w�]ל�ac8�7�
|�!�=+� `kkt�Z�����
�Ve�S�
���0�d��͚R�f���j@7�_;�4�����YN~mt3Ȣ؞\�^�b�s>��Rs0�@Oq�A��D �gQW�^�n�B��>I��)sg�9�xiMP4�=�6��3,�O�yeP�Z�&����{�_NJVX��j[�[GvbF��YD�?Ò���7`w/A������`���JyK`  J��[���6w$(Ih"�{��2q��lwܪJ�G���ף�+�+!���5ehuw:J��s�F�+bV��t�UW�PA���d_W���fC[�끝r���T�k���H���Ha]�^Y�Ń�5�Ҽ�r�3������>sp��>�~���%�Xo���-/��KBI�5��	)ˋa ��}Ǯ0Q���!�KwB��V�j^�t�WJP�A�����S��Q6���=�	�^���C2>�px�Ot���C8�����O���K����]-�ƅ����2��IH.WD���]`�ݓ��VM ���@��Qb�;�f�Q%�ח,���3��a�;:M��"���<MQ�=��'�װߣ�LY��7���Ю������q菴d��$.̐(�1��#rn����9��wP#�>�:�w�~�'�(�&p��Yp}��u�� �����MUx:�_������)Lm�T�%����\�A/�y�O6���&hjV틜g�Aŧs��3��NP�%�PcvwT��q�L��#���d�5aF��+�#�H�Q�5jG�e;��H#�+k)���ai���U�eb�Aʟ*Z�~3p"�TUo~m�G;���B�˞�9>��P�a��b�#7�+�ٳ�uP�%d�#W=�(&UW����}�����?