��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h���]��ZBq'aN#y�L��,�&8RG/���.Rh-��/� "	m)p��N��ï�li�δZ��U$�/���зk�BR�:���M��BCz��I���>D��ߍ6d�m���:�!���s���{}��ca`�f!L� =q�^�� �fggK�4��[�$��1�)�f�p���لt���&r��<p���Q�H���H�����%-Z[����*��]�Y ����I��F��4�[3�t�#U>�̫�����"a�9�Ls�k�C�Y�l��`N6m�$-�b��,�&�
����@b�u?Q&�ߜ��0��%���|\�T7�ۺp vJZT��&�#ܬ��������]��O����Jg�
d�8��5k;�������f�[Ac�pq;��S�)��>պ��,�:;�r���з���կ�B�����h��kcT��������/l��vb��-�^�9M|E��.�y?�(���vI�w�d]r)~�v��R�F����M#~v��K�.F��Ҟx���k|*���M���g�9 �w	���֓�lY*���Eϑ]��dx㒁���E݃��M��7O�����;nb����A��������\m�E�<xZ��Ns�-I[����Z��5�[F��B|G�y��o8��<eAZzw�m�\m\8M'�DX�4���k�B�5pH��u���nX:�;ǌ@�P��x�����\D�(�_m���Sp�*��ʑC8��iy"������L���e���p� ��.�LP՗0E�4G�����FND�C �XjN��������犀P�ۃ��o���(��m�۝j��4���̖��¾���İH��\���p�B�;j�{���Q0�Jp�3Y�׊C�"	]m�"�萙f���b?�y��T��/N�$�=���-f�.R��Ο�I{Q"y�Aу'_x1�;35Sa'74��
#F�-�� ���l�Yݿt3�K��E#+�qE�V�����)(����������K��qd��(9[�9)'��~�$��9�������77�fO#�su]���`��@z�!%u���1jT�ii
čv��`}WM�b��Q�������G�4"�vm{s$�����{�L�^�zw�N��@
r�T��X�[�QnT����̝DL�@Zv�`�
�d�b^�A�kLx�͕�nvt-:�P�N�.��K=O��'�y�v�����X���6(���0�hZ'2q��g��^��ۭ�V�W�BD�EWx�����,�FI��^w�;8a�H$�+}�b�2o�;��N��"6k����s0�a����)yD��c�ٱ�Ŋ|,��%������1�FS{��d!n�X��[d�В:�m۲p���ƅf�L��M�����w�Y�/���ˑ�p%��[�)��'�9���آQA4/�߉�r���'z�2�Oc�.�&�Rlqg��Eњ���&�aʄi~9��A�Ob���
R���
��/R#)�O�RB�^|~�=w�)6���헐��M��˶*�@��	޷z��)y.ی�R���!/ye"���Y�0���ou��7�/u}�.�_X���V����+f�Pl�\V��O,ADBFR;������aY�N�U�S�����T����ʍ�pQ*�hk���$+[��@+Q:�"�i�h���]�+�㞼���;y7a� �ֻ@f"�i&�__��cI��P}��	s���v��~�-�2d��gH	��I�7�/���H��ط���~�UݘD��O �ǈ^Z5�Y�&�%�KW�r��~]��Z�XY@�!���/#`��{�7?�'�4��iz9W�+�ζ�U
'��2�N��g+��,n)+=��z,C=����y����ڞ�dm�~eKL���}��ts6W��6+m��R��]����z�=X��B:C(�7���Niw�����
�����}�23pg�=C-DdYh���q��4�&�����ޝ�zYk~�M������t;�����5�k+C���Ո�9��(�?1���K;�AO��J�}�윢*l�j���Ҟ�*����/��a�%�n>���ѵ�GP�"l:��w�ǿ'����9i�&��aG�C>XJ����U5{��*H��7�z�'w aW^��L�K�s(�*�<� ,!�=�K�&��7�#Rq�f�\-ò��&�|1�K�������"}����*��ͻ��+����S
T^D��_�7�@u���Pա�$�z���˂%˙I!d��mN����#KD.r����n&� 7ښc;��K0t����&��g����ޱ�H��\n��G�9KAF�8�2�-�2©3��Rψ�D�N��>1i�a���L�L�6S`�]d�,�6Z�]폯I�D,�m?8�@2��f��߿���&�%� �Z`u��"�0R.�F��Q9�"�}i)v��@%�_��[�-83t �j��U�ێx��t���e��n�I�Ό��/z�-R�������D��ذa,|���ߍ<e���$_��~O���]RI����w�C�/�b���ob/�y���oM������ߝ1&m7/�,o����L��_H�ǫ��&����L�k�5���W�Q��C�ǣ��	'+�F���$��g�pQ�Ϭ��.�Wq?�~���a$�S:�|g�Y�t�n���n'n�l�RF���.���q���0!��2KH���Ui���^O����p��5�I��+�K'��ǔg�V�6pB����ұxy��Fj����W�1�52K0��Vp��e�wH=���ɧ��D������	�er�/:�4�;R&��qNJ��=�,��@�lɡ`��e�`eM���76�h-�����B_�U�yv�\�Z�2�M��������n#��'������x�>T�)�a��F�,
�T9�q�����&�ԕ?ῃ�|�$;g-ӣ5��x����X!���{_�	��?��9���H<�<6|����$U��W��>�y5���=�<G7��S��o��~Qc;�R�nD�5��F5��ֲ�
�c0T�4���iZ����ꠉ~H�2ǟ)]R.����c¼��M?�D~�y-��}��J�{��eܦ	ԚQ�ۻ.�@PP&F�B�P~ ���"�PE��:ۣ��������-u�C)ߨM�/�λ�������!�^%?\�ۧ�C�DgB1��V�x�%q� ���rw�Z��!sN؏�p�����`��+'M��/v%x����xg�а��`�ח@��)[�B�1��#������Ը[ {Z0�B���)��G`�2
�����)�QX��
�1���fP]9Ytb��2\Q�}���V��.��j�D ����䶆e��I��P�>{����U��B��Ў�}�����1\H��0�s2��.�2$9	+A@ŉ)�K�}�mK��0q�?�Fx�ic<%���:�u�k�h�r���X���C~T���Bx���7�=
KB�4�=ꙮ�L�v�u�ژ멗M�S(%Ȃ�䳱�%Z�-���%D��2�f�H�勪�f�qβ�D/ū2��f�O�r���w�5��`0�볩��s9�l��3'������>�cx��4�U�����|���>��g�.7f� z_����I]vlݪu��(��W2}���P��Ml8�Ұ{������q�f�u��g��m��(Y�J0�����z����`x�+�J����S�j��+3�$�	D>/�L��hY�.$@.@�hVg?��#E��Mj�H[=��ܳ� �Wd�#/ct6�b�L�?�ԴC&�p��F@/ �W��7��luՋ��??�,#��"�yn(� �� ����1rf>Ϝ�Ġ�Y?ݾ�PFO�ܝ3��(%s�����j)��`���Y3�F�K��B�D���_��E��S>�y��k�6 �Ln��'G� %%ǌ�rE"]Mi\��/Ʊ�@~W�ڎ$�p������{��f�}޺�9�Ï��=��_w�,���<�q�?�d�S�҇e�K�e�1곮KT�T���7�/�7�K��E�V+�𡙑 E���7��L�ę��g��������P���*���t���f�®��=!�q*�
�N�`kK\4�Vm�]S�0R�+��el���\�h����gZ�����WM��K�B�8M
q����D����r�ڜZ�~��e�4�i ����Y!��p��qmE8)����˜�����B]#��o���$)M�͂�	O����V(@��ү��z�00��v9e|�c
�By�]�5�'�1���`��ާ�ǰ��K�G:OjSs��^���4&b��� a�O.(�t�wp���8�p���_�L��3�G�����s%��g��[���xU��v���ԷJs,�a�]��ݘ��|�d=D��C%r�h��ǖD!'š��8h�ᩦ�8�;���n����ub�y��� �`�������J�<�����p)�.8�:}d7�JP2�X2�F>6�{ǿ4��w���̄�x��_*a�p����>���p�p�n���&�0�y��֝�O��Fp���ءb^��V��/K�)X�7Џ�ѕ�ؾ�u�Nd�����
�{�k�f��	G6�	Y��W���5�� �$�EG�<d��Wá��:\qd�1��oॴ�u��]7^��r6#��@� ��O�_���Է,9��X��:l%��}���F�<"��,��O�.�/:�xcZ:��'��w�Ģ�I���K�#�e��:8>�+��gJ`�dFL9Y�+Ӓ��W�R��x2i��ŊV�\����'��x/)RJ���EO~))�P~�(�I�߆'�,�+{�v�D�\tV�����;�mWA2�YX&���ћ�?�@C$$���\=c.k�.�2ȁj�k�h�y� ���A_5)P�;�_F�K��x^.;�8�\��W��m��&��Z0�����g�s�7� 3�qh�h�G�X"�$Wծ :ĕU�X�&�S�����6�ޚ��V~��+^:�	%��(�'"1MnP��P��`�4)����O
�$@�W<^B_���Ψm�aX}<�8@��Pc�w�G2-%�!�?�[!� ,����,��_(x�.�^��ػ�<���*.0���}�����\{ �\#�-��G�C�FB?���}2|���"��.��ą��zRʑ&�Qy�v�?6N����_���s��A�^ߓ�"e��W�2���@H����~�o�F��g�n�z}�u�X+��������n�e�u��Wlu�'s(�٬ާ۫�rp[��][��Fu$}�~ߩڬQ.�c��f2v��#�KD�'r$k��l�\g���V����Lb@v=�yS�F���9�C�L-����)q�ٗ�R��93�ra ,�$�n��0������A��}T�0Q��W��@�+b�?�,�$��H	���p/dJ�8�� �.���VT�z���W}�gm���܎�v8�W��J�7�by�>�C{�S��
�yޤ4�s�Z;Np��kGq?܀|VʐH�m������
�����(��]��X1dl�<�yG�zJY}�0!�q��2��L��~�R��5�6�4�x��A�Vi��u_,���ڤ]c̈́6d��͵��i����W�򿂋s��L7�n��V&������L��V^3���tO���
{��C#F�s7�7ɜrE��y��A1,ªS�����*�?��kCΏ 5������Q�7�Z���6��l�g~m�ϫ�\Q��>9�Cm�Yу��U���y���|z~�7V$�p�*ȶ��t%�G��R��*p�o�L�;�� ����Uvxwr�EHE�l$Ly���C��g������Z����\D$��ֆ/�Q��qs5؇{�T[��<�V;�e�@f�Ue5���Y�,�I�����*��h:�p����>�� 	v�C��*����C��sWv�w�f7�#m����F�l��-�+p������~��	�S���p�l�t�	��?��	�X�(#��S�a 4��VZ�8d���������tDEjT|m~9�l����QE^2]yѧf���<�{ڰ#ɽ%���[X��ܨ��/��x$����X�:,{%�\|�!�F,�ҋ��*�{��ZZ���]-�W.�j�i'�_UR� -�\��J኎��<����v*�cV���a�����"b��@�Z��G�6�q��g6�w�OV����܀,b_�^��  ͟ �u+�%uz/�*�GV9\��F��	��Ma��^�٣>oj�"`���`
�H����X�&�z�깈�Y衔�Ӗn��z̳!�rn�p��f��yC�^�Ǿ��y�?+�s��מ��3$���z��B�?i�<B��8C �݋J@�(%g ��I���>g�d�zA@D�oP��:�\��R���r�,W����][��ۍ�\#Z�Ց�����ҳ��e"����K)U����|�wD���Wǻw�&7i����;�2�sdl
��v26E�/��h��F��,�g�=k�U>����!�Š(Z�
M�o���"�^BhS��,r��˼�=�M���f��?�{�ju��+8UF�M~K�F���T�dW�����+�ᩲ:��w�g:�Z'dG��%�/m|Y�o����"ܫ�����|���y+��ZP6hUT=v�ď�  �ٿ�0O\p��%W4�'��\��Q�eZa� ����[ޓ���5�)�Ċ�K���a#�6�|�|Z�kJ� V܁��c��]�k�PǮ3Y���i�~:`!u\c���
�9���hk��u��i˘��$��l9�`��%�6�2��Ʊ6��ԩ/�R���L'd�@��B>�r:�>�K�����/����������^g���<�����z�>�@̡��u{%����wF�-&�m^��w.X��E��OMDv��ϩ�3ҵ��3�������2��J���:�m��Y�W�<.���������j����(BL����˓[�uN�,�x跖�]mOu����q�$��ο;Ŧ��^�"�x�Fc曶�\R���%�D�����J����U�����Q�Ŷ{����m�E���h;f����эC�Q�D�]�¶�8��3/d�g�n�1XoZ`b���Nb��Ɋ��
�?H��o`����D�	f!�M��b\ 	�u�{�w[�s�������ޱ����
	�pv(��	����,��U&�[�x�7�������M},k��'�~�0����?��h$�۵��<|�jUT!��pn\���@C��m-y�\���ᷝ�(��odA���D�LN	#��;��W4����Ј'�\QSx��d~��a������Hn�D���`�*���VOJe@?�*�(pM�)���uC���=��U&Tj��e�(��l����p����Yq�H| ́����9�mM�y��
�˹u�X�SLg�O���@�����C�,F�
,�/��?1OU�Kx����'5�Ok%-���6Zhp�$Kz�짩�Z*���w��_�oG��s��``�x}�ߧ�#���Ͽ�ڹ5��)��M�O�-�C%�V�n�Ɵ��b�Q�����5L}`4ȥ�C��aw�h6~z�썍uH����ƭ:�6bͮB�B��W�4_&nG�d&Q:܇� ��%�S�� ������H�ZVwA�=km�hn����[��_0���w��z�Ӟ�ԕ�5}&C�>8\�O�?�X0U5�bZ��Sǲ�1/l���0��/�T�:�z��O�s|�5�Kn��1���Hͅ�u�&��Z����?�K����H%��cR�}	1�?ꧪ���\Q1���N�����g��O�����5����c�����C��Yq�+�tƍ,�,.�S�J��L8������8ϊM�'x����Q��'�0S)�|�r����?�b+�D�]3�fr����`���x��&=���9�S'��s't$�m>��@��\<��0(������9����Z�]�eY�DU�K��w�qUطL>�K�P+�7���w��hR!�H 4��K�J�u�"��c��Ȑ� �iL �P�t��<�gs�����,�I�S�fx�(@K�nx@��PK��(��~-�X_%K�nU�X�r���%%\"(����W%+ �h�p�-�c�)a�sS8鋊	���@�����R<Ҳ*� ��zY��)�XN`�Q3<.�����vp���"%�ӎr?�߯RyOw�t��������ajptNp �ÿ���t�ì'�0�>/Eϡq���zUv�����#`f�ɾ���Kp�j�0�ѯ��c���*T���SO���|nQ�b*g�����?�ս��e1���l��Q����G�����;"ۢв�l�;^�2���?L��(���i�G���Q1⌔a�
���2<Y�� .��gP/��q��V��-�/*y��ɝ�n�I�E@Kd�M����b
�ç��┒D}WS'6�1��qY�D�F^r���Q���T�7�eP8B��!2�f��c��қ���-���[�C�c_��n?�c�7QԲ@�����#���N��>C���8�8h��`3.N�W�e�N�[=(� a=]{���-~��pD;�^L���?��l��@_�k�d9�����OQ1��c���g!X(�F��G	I�&ZE*z�S/$��+�!����fX4�l���/Ew��`3zu���'t-z����#���p�e¶�đ�{(��'}�����xM�m��2r�I�f�<�LV�qW��⃚��ܿ�㍤p�d*�>s���'#�d��,�\�!�m��6�a�p��b�� a�
��� ƒ԰H�I�r�ӕ,��f#Eq�$n��͡DU���;C�yg%�1����U�DjP���ǡYE%���l+!ߌ�w��<�_x5eO8f��}�KثzT6�[;�L�Zy�1�"�ۉ�]��,(�癸��T�PHw��mh�� ЗM|TC]U��h�$�0����� 	�U,��H���>T��Ȇ�ҫ������M�x��h?�0�=s�bpL�S�t_��S�:������'�f�օ��t4��0�v��,?�-f�P�?�1���d��lB"�x�f9�3%�H�`J��^V$#�R���&�3����������$�$���B\d���KR��6�W��}��rY=P���d΀�B��l���{Iq�X�Pl\�Cq�2�Ha�Q��ڷ�o:k[�E���nlb��hjZ�2�LN�S�ŏ����0���CƄ�l��,#�aP}^(�ǜ�[�B�r7��z�������w$��!3�EnlcM��B�ӗ(#�s�j"	�.���\8�a�����}���Ԑ\B|}�]�mHtM��[���%1%�!�K��ޜ+�S�D@0�w�l�V�e�&�(��>4!Q9Y!:�(�ײ��ʷ �V��i�2[L��ǟ��g'g~��#�����['�z�[絊-���~ �~Mvq�j	�� C�|��OV���H�5r�9T��:�D@� �O5�Q�c�@3�3+��1�jWy.�}
��?h^�7B�%�Q�7D������O�j6\ڑ�N����
/�(��(Ll�\��
����Ny�Pr~fU�5Q�☤lhZ�gOv�{|��ݷ�Jf��-��f9q0�xBE�2�KG"cqn0Q�D)9�*�ws�t�g�QX���.�������K��/�Y�MG(S?�(SD��y���F5��c�y�ǹ_l�'*�o�
����B��
M"cK=v5E�[#����c'�>�-7���w=�7J?+rN4����m�qͩ�QJ"R:�y�H�����Rz]F�Zj�_�����Au��79��j���;��
2�E01��O�4(�����3p�% ��8Ko�5ey�$�N��B^
`��^_㓐 \�}�~#��y�=��p]�����6�C������f��S���ףoV�>@���s����4|��MDoo�-(�=*���9�w*�Ԡ'0-x.@�����F������P2���/􊑅��K�z�֧�ޯ�=	��5�g��Hm����� Nm{-͔����������Ӌ��P3�1��J*�ݕ�df�$[z�Z!�T���u�4�EyI�!�(�딡�k�w�;�S�0�Q�T #���A��þ��$��$��|��ʘ� ؼ�=�ñ��MU��ƕ�����m�pɝP�^���A"���?��"��co����T3�_O7�[��K@{{�����a:T���l�ý�|?�a>��(ȯ!��뺛��g��sl��� �d��0n�'}�[��^מ�(��ՇWDU�ݍ
���DĤ'��*�d=���%7���oH*��s��_�]�$���f��>�7s*(��1	W)AhFx�9�Gů��Ӝ��d���:��ю�j�yB��M1w��[!g�ez�����jo!�O��2Z�1˅Ӻ��ba���%� � �-a^B�b{��SFF�ͽ+��\���#W-g��~	{?�fb��4=Ό��Y�7i@r�����-N:VD�n�uW_?�{�B��r��׀D��{���.Ĩ�������͙�A�@@�'�[�'�8��B�6ֵ�-p.�`3�4�Z��Dn,��ʑ�-@'�O����)z��� @n_��
�g�l�*JO����&a��bgN���Z�K>���
@xҍ��#:D@ְ�y)S7T���w���0ϯ�<
+a]U�,���ck�l���Y�}�TɂjGNVpT�c'���3�
��q��D0��B�!D�.�����#ԋR�E�������5l��s�����{?���KƢ2�s��l�ס�L�����	�W:���	7��_�6��ق	Ƽu�y�xkʝ9	�aU���������Oox�0�u�\=[x��a�m��r�������@�nv�;��)�Ӊ ��(^�B4c�U�?w��uI{'�do�g%o{(��w@�A��Ea�1������4t���@ĝ,��~�6V���#^�҆��V}��j�+�f��!e�����O*9�~�fo�����v�[:�D��F�Y��E�G�9�"%Aǅ,5�_��B��0�n?���94���D�l���rNqSF�,�V�T�B���;��;�g֥�d�� ��ĵR�"��D� M�;/�ll���;Þ�z�`k;?� ����_ˢ�X�;r��@�Ǳѽkߒd��-l[���P�ء�U�mg�P9
���,>l?�Yzt�O׏4�Q�o� ���z0M�ұ����7_č�^��<���z�0���� �?%��Va�Q(8�.s�w���|_�$�5�G�����%�
��`j�t�!��<zl����6�0�Y^mJ����� 5�A)P��>������9�4)��o[��-G(iۢ
'$����4�������t{����2�G�Q�
T1j�}�E��4�X����=aVV�w�to�A��4�E����P��uy �����g� ���g�u�J��}��M!	�c��J��QW�_�r�<���m<�Ղ�H/K�`lA��u��9����%=�KV�@����I<�9k%�I��_B�Cp�BbJ<S�0�(d��"�����o�z�Y��HX(��~	\�:�C�n��ic\�*a5ZoN���������^�\�Z!	��\-�B]S�~WY��_���GG�������Ay�v�-��4M+�yoߖO�`a���C>K!��Q��[�������G`�OD��b�������l'���r�!qR�g'�gt�&��~�
�?��]��!�]$J�^o$��.�d6
���<Ҹ�]^L+�*�@GlgМuA_�?b8$i?f��Ny=�ߵ;e�&eM��z1�<a��z5�&�.���Ŭ�O�-R��X��z)z&1,�o�չ��E�f��� <g�_*��^̃*Z[;������I�R&#��EA2�w���F�;�~,��/��1gtҰ&���z�{OY�ڏ2�(���Ы�����I�ݳ�L	�u�����k�� �K�'	@^���86>N��<�K� Ǐ��M����=�R�T0�fߖGb�7R��$~�����ֶ�T= P��qJ<��"zSxH	��tl�,|�괢Š]GW�7N��A�a��������O7W8��dD��,Ǵ�.������������ě9v�֍�?�dh])��z��N�Q8#�~��|����8�����PHa�	�^'zL�
�C�8��қw��=O�]85r�~�)N"kc�{{��V��:�=����b�MbI�oז_��?����[�&��S��������2͋M��N�	e�S����ˡ��{:����ޘicjMOA�^K ��m��Ȩ	��JƏE���+��xkO�#LC�b	����Tw��8���27}���Ә~�py{�w+ӆ��x�����%Գ` �l!1M�])���6����r6M�$úA'��g`�<]���f���a�	�����ƿ��Q��X�{��6�����Yd�!�l=N8_�0����D�w�O_e�&�����2�ʙ���=����7���x�,fs��Ϧ(<�Q� �ɾ�EᲤY$��?��T��i���>:G7W��7��rI��2��|_��4ǷӨ�#�����+jC���K �"o[2����Ԅ�;* C����6JIO��o,�P��PNwZ�_d���KsNA�^�	8K㥑V����9\�.c��wR˝�qq�I�[ˁh��_/�{b��,+���Ԫ�2��i	�i_$��l���!�E�#�$�鿼�p�N<Y�Tx�̨�����s�_�����r)R�` �G��0����uj��C*�xqs�Ve=����4;{����'��H����o�8���dw���i.�>�	S�5�Mv:������W�G~8�6�a;�07��j �&x���z�=�f�2$(�`n����og(u�Q��KFi��� �CP�\	s���0g���(:U�;�H�Ҍ���,�&��Ib<.!:�[�qd��'o��i���Fg��^���� .Q������
�8�u/�M-�Ù�%��n4*�_���(�	�#9�׊�k	ٯX���N}����_kk14�dA�?;���&�=��2���X��f^�Z�Bn���Aȟ�V9��u?��|uS����4�1L�<�6�5E�s��B�������1D�N��y:�DEq�7�>�X`*rPh�}r����Х��.�k'|���17Ļ���{9h���M��L�;�����ڥ\���xNa�q�a	�pp�v]Ɋ��'	�F$���	�eh��qi������ձU_���L���W�^���/X���0����W�1�R.%9o .D<^�Q��1�;�NmJ�Y��+r��+'�RD)�}�ٿ��j����M�4������n������R�`d@Z�]�9�+�� ?�xg����2/9��,��l�rw����L����7)��}X�bBv�vzbe�@/ _��"�����rGUg;�~�C���q0�a�$�"��z�n ��&o����u���B��ׄ����i.w![ٸL�s�z��iK�bR�O������b���vn�����d3� [0����8R51Ya �-���>��) %ι��>��p�D1����{�:o���9d,�AM1�c؇J\<�^ �Q2xy[_�J0�"��1�qyt���J}���gv��L�V�e�&mk\�_y�T*�E{�.�/D��<���44J�̉���]<�.�u�����9V�*`8��E����Z�=��G*}J����N�&HJ���L��_�]:|��R�H����v��O�t�:w�� �nà9���kج(fLr}�>.D�v�GB�p�w��e0��r��ާ��������#�%�3J�OA<'�`���*���?,9*u8&r �8s���J,]H�/",L���"����*�۵����D��S}:�cөh���� �A��q����z�&�d$t^�5��HD	�9����"b��5+�-e
�i���-��L;b=�]vgh�ſAX}�3?TG{����RF^�euj��]��+���'s.^����Ō#��Z<��,7�"�����J8ZK�:-��@�e��6!j��[T�4j8�]��z8�!��_ ��¹�������g���zw�L&�9I��{�Ԋ�j�+3�	 [�\&׋c�{B�����-֌���N�|���8P0����*0�gt�y�c�FKjq��(��n���I��<��59���W
�I���d�B�o�ݨ����y��%�R`�G7���յ]+8e��۔ϦP~���zR=R�Q}]�������~��`m�3lΒ��h=I8w�#����&R=}픣(��B*�y��OEH�b.%:y�����I�Lb��4-xr�D�
㝙�+�ᴘ�)�&�oP0�(W����ǲ��Ԯ�r�z�c�`���j;���r�~�lq,��C]�̀���s�9
����<�
N�1}��b���  ��ݰ���K�.%ݝM9��W���bߎ������ϯ�_����ʭ�����Rr��Kh�3{�5�%u7��l��|Ke�8"vJMvIɘ��	K�4Y�k����R�u]��)�]��I������(�.�m���u�i�P���|,=�M�V0�#C ������'���g�B��M�s�(��"�fPn�`�B�J��knB��~���Ƃ	��s"���QoC���`��eo��S�Ra��/8-�9���uFp0q�}3���yLp*�E��<�D>�P�M�[}�����o4:5,�:,@M���$7L?A�8g[Q��%���>��`�y�S�{��jJ7��0R� �"���܈�v�Q����JB�ӫ𶌁E���9q�ep=��dy������^vPe~k���Q�>�@>��0��"��Y���i��Φ�*������vJ��꽗N�6��j��?F�tq�ST��z���p�w:	ܔc�;���Z,]j@3�[�E�/�� >EhD��y)�(3����x���i����z���3c��oű�_2Ʀc,c�|�����ZU��0��6���T�9h�g���ͻ�a��|ˋwǟYO�fF�2�ȔY�
�K̜�һ���u,�Z'S�7r�����SL����'��� N��[[-�rn��L�*��5���mM)�s�����LZ:��J���w�)�s٭����噊Р�j�����V�36����k��
V0Ct�5ޮ���b�8����<�QP8B�`�q�93�6��~�[�6��~2o3��w �>�-�Ś�^t	-�f����[�׬<��H�6�{b�/$A'�+��Q���+�����輰SgI�M�({'c���;1\�H(�m=%E�y�o e?1R�D��^2e)��ъ+L�_�s��K����\�x���o;�X�����1~{�>XOI�޿m"d�k�j�x�����_QXZ��z�2b*O��C�/�4�][��:���tZ�C4��D̪�z�����
8C8����Z�Z�^[��H��S��q�U��Ƥ:}�艱%}�����{����E�u_�� ��/�����<�VିP��7�iAi��RF��z�r�����	��$�O[*(4а7Qh9 ʗ��H<1��woQ	4�%�f��1�}H
V�ه_G�9<h�:�TK^�hOQ�-4���7��dF���}ȳjn��gz􃁎i���^m��
���Z8j����d��Ur��Q�/�Q;�ad]�ě
k8����F���Z9���s7��Y�\�b���W�EٍW�d��Qv�	e�B�a�}lu�U~.�6�/%<C�������o:핢�%�p�l�]^/3JO�/��$� gD��T��4xr�U�&jù���S9��;��Ě.����u\��L�-p��!�v�;fj����}k�{,%�^b17���q2g�E�&<SYD�7�L��7նI^����������+1�X���!�Y5$E�2�g���� -�z�6�r�gH�9�����E�!�vM��;cϒ��ϟ?�$-��l�r���H���ʷ �ݑ��'�	��N/b>��X�H��|	j���W!��:��kskC�\)y�TJ���a@���ݘ.�����.Ց�	�bZ��f����m�2YA<p$��qP���GN/���ri�>��\�1��������WSb��tL���bE�?��O����ld��7\�����v�G�i�y�������7X/��K�fK��V�ESʌ�!v��z�`X˪�@��k��E�7_��(j
h�V/(�X�����.� 3#�N���<�᳞MK̊,Pq�����,K'>�uT�q@�Db�t~�=$R��5C[� {F�k��/��:!1{X�����g�F!؛�`���/X��/3�S�.�Dk�(�� ���4�5|�� wA6�E�tSC���x�q���'���'FH���*z|͌w%��,�d5|B�)����f��3w���	��	=^/ffv!�w:�}�ǂp��(!^G�f�Q��x��,uO27l|��K�;rT�/�d?���JgU,OPK[_f9@�f������2��*��e6]�5�ƉS/>"*QS���
�:��Gq�gU�}?_,����X�E,�[z�3��+O��'gM�O8y�����!t!f�鉹7����vj�a]WUJxrȀ��>�T�cK}}���R�%,Uه=zj_����Z`�m)I>6��*Od�=�_�zA-��Uw�:�_?Z3�<B�,���#��&ް� ��v�MO�w��RPnH� ��4��y�*M�T�1b�Ӗ��3�F��9��(V�U)I��m��F�]��@�ˀ�Z3m�9��ն��:���16ϱ���N��{��^��������8����ÑK	�0l�2k�5S.t��"��];����]�/N�&�AA�r-��Q�2�e*��{��j����ݝ�M2���8*�eb�6�lK�pg����1��T����j4tZB��O�>�<�ե}�xQRӬ�`",ެ��ZglJ��7��C�e۝,�m�y_��Y=l����C�ǸÇHsI+��=�sq���#����ER�ʱ3�z@MH����J)�70���.٤R�F��A�␀�P��mF���:� !p(	2JM5�;8W��9�x�lV/P$n�/��/��H�-�
"�^
�^����531x{6�rx�!�fQ����M����*?�t�SsQ�ÛF$!���̚\'����/�t�¶J��Bm������YBZ��lB�a�4��,�ܫ�FT8�%��WT��eVF7���M�(����B���v�e����V�+�^W��� ���<7rG�r�56���9��I��Vn����@F!�2��7�3�zR?���)u�Ep���q�3�1�_��+r��b�k�4�y�,���TP�퀑��EiZ��:�.��eݹcoƻe+ѭBDMaշ�n�=�ݰ��Z�\ ���2� ��7���$���	�ٓp�M�~���H��n]FJ��S���Cvf�\�i}��W��:X�E�Ư����E�l}��C:����(���/)܈}`�P��2���h{4�oN�wkkc�k| �j��~��L�����ߪ�����E�_-j�~�,>Ř��<����6r���H�$�<?���v�/�
�;5��<O��&#�]�g��)3����E�.^\3�|n�-���ug�.V45���P��u���<��Q��?��2�$�0Z���oʩz͊塵&w� -	�.I
E-�:�h�v��rx�z�S�3�/NtBO˴9��$Ճc^Bɯ�}t0�+�<�����p��%Rj�8��
�;FW�z �כE�{���u��V�Qnɰ��ॄ��CPފ]f�p4`���'v@�����k�"�ŷ��(AK�v��7Y�Ka33X����3���kic��Z�N8',��k��,>��ta�w�����~�H^�|z޹G��J/��X'GN�O<C�b��LUX,f�cs~đ�vB6�[��_~��E�o�����YŢ��n{<B�6���kՐ���U��A.�[�i�0wE���mq����V�;��ݴ�vHˍ�f�K,_������EG��+���$*�,��3�)=Ƿ�)�90\M'����?&��.?Ŵj=�����Bx�m&Sg�<LJT�	��[!�1�`�
p6m�����Y���Qvs��P��70�f&�f������B�x@�����#�=n�QTpHx/�(U�6Y��3;�6>�d����͟�~?����a:|�������Y�	v�亜&��V0�DYT�0t;a
a»�^ܑ��<!1�F�M4���)��Ks3��Y=q�缝6$��j��f$ZV�ؑ"��	9Xa@k���+�B��"}�����ةMo�v�詙I��4��`��:��Q���\D���9�W���,,{��I�Y�TI���� NU-���yL�M�_=��T�KF���*R�]�ө#⧄�p�� N�%`n9uRX��1�����5�J�؆���z�@�n�Co����]29:3;�f��FD6!��\<���1X-�?��㖼S���zx��f��ơB��K!y������셡�ƬA�Dp��ha�D�9d��lĒ�G )zM�k#�`$��5��Yڡk��%�>�3��ݯcyUXC�o����>1�%�cIK�+��Ӧ��e��������S�ʻ�Ƌ2��.�{&�}+����C�zn�H0|��5*�� �x�"��,�(v��d�4� /І)��/D3�e)��f|���T�,SNc�"�;R=Z��"��&�q�5l�%ǻp�>]���i��ɗeR�t�O�c��A��WJ-R��>i-��f�m<x�S����Q��wn�Q��W&���M"�#���]����wNR���K��g�⻦�µ�YA�m��	�
��ɛ^��:�	��S�>�r��%>L�Lyp���԰^�y'���|ۢDPn!K��k�x$��sJF\��YS�%)]hK{���8�f�q��H��;��;�:��05w�8�!=Q����ǆ��TD�'��h�'.R�L�����z�KM���}��V�n,�\�s�"�t���3�z}�����`<��p�K2�z䅿�}>���Bk,)�U����$���jI�J�X=;M���������2lE��V�Mޖ�Ə�9ȧ--�ͭy��noZ�5�b��i,��h�qC�eC�����C_W�U@��d�L��l��-6���X�$u��Zwc˽	�����=Ȼ���d��(�UI�0t&��s�9�'���}�h��X#����=�ǭ��lm��\��Ηq}��
9@po�4K�n4P��W)VNERU`xƦ1ne*,�X!(��̜TG�W�^�@k� )�g�9���䯵�Y�k����$M4�[����D:�9r篕~.m�x�mj*d�l���h���F�Q�BU'Y�-���U3F�s����l��Ƣ�����0-�����=�5��B��|"���_���M�#���6vp[h>G��+��j}D�>1�qr���d��d�#�#� �������\�{��T��`�t�(|��V�=
[_ղ�DXQ�6�f}$rG?�������6�d�w�G���f6��r��tu�avo	�A�[蘬~z왅F�1���I��#�GϼW�W���an��uJS���������ǡ�m���S:4����O��D���c��F G� ���?C����m����rH����Y�5������L�{rm˾]9�*���i�agG����@睴&�Y�w/�ʼ2�7t����4�]���H�1{T�����������)�!d����P|'˖k�8N�9��w��˶)!���� �Ln��HV�uh}<��#�<�˅S��:�N�Dg}�W�₤'�%�c�Rvl����H�gNW��%��I���~I���*+�����hb,˅x�g����yu��'��JԚ!�%NK<�~N��c[�b���q�)+���}��!&���5��8RI��a���|��l���B���kB��Ȫ��[��q�_������XH�܈I+�9n�vD��cM�ּ�<�LZ?hR_W�G�s��8eú�`ܸv�~�Jgq��ُ�s�Æ����}f������?$�Oj5Gf?z�I,��O��|�A�.c��O�]	՜����1O2G�l����2 D�O*AU������]ܝ��D��+v+;슸��jX���N0ĬV�2̕�+�i��jf-#�N�7��l���O��S"h' L ��F���n�d���YC<��m�b��74�t�|I�o��[�k��o^���������.t��1���dc*���C���Q���&�3� ��pE�ޭC��1��8~F��P��>*-ߎ+-X��Bef+�����n�*��[E�4}6\��	���mm
鶌75�$Nq	W|����O�H�0���_/ �xi��2�Y8M��>�x�d��]����WX��:S+n�[��ˋ�����QD�Z����#�߇��|����TZ��@~�gYI�>U����x��߭n9HRP��Vq������
��kB��<FK���m�_W$�h��o>�g�Z,�b8J�!��O��k��Mu"N?2�v��b$	F\.U1�;�0�i?�)�7�2���nyޱ�*J�[j�v>�<�����_���LcNұ��ƕڄ�$�4�L�~ {�t���	�-B�ν�H��V��.��؛�x���ƚb!�@V;���P���m,�K��A�?[��M�.��l|Q�0��������o�J׊��Ы�T���ٺSt; 	廈o��~6���<��ɶ�}��@�Il,w�Ǘ		\|�!9b����?�h��j�{sd�"�%�2�����mnIy�cq����M����Y�t;R�Nг$Y
 ��4�,|�7�n�PL��9�_�a���>��a^�(���$	���º��i
�Q�[D��3��"!\t5�y�K]�5{-@TF��H�k��k��]�=ڮ��k5�5�-@�Z��$������y���$:��4D��s��hC���8���[ ���8w�<�c$E��W���o�ί���l��1���a@|�M�2fqveR�5P���s�W���
,k0�ǀ���M���L*�}g�R�J�#q�w?�~z|�����Fb�a��=�"��ؚ��ce�!����� J�b�1<j�ϞT�5��H�в.�Q3�gsqVo?�C�X���t�d}��*�$~�S@��hA�H��}�6���Ezs�Yg]�϶[�G#5�4Ɔ7����`�P�u�e
����_@:3��<|��އ�n�x�'3�?O�g������IO"���o�&%��`[�R����}A/��z"��M8�yU�t��C�+jc���AtI
bZ<V�ΕyHq�1��W.�+�(<4��Ξ56 w�"�pX{�H50�1--t���@C�O���G�Z/��7��ĀC.B	�^����q+f1�/��B��"n����WM��Z2��y@���v�8�e���3c�dM���]���wU�h��/R��R�f��Ȧ�7{�$5Tc!���ݴ�lO�*�j��Y���!�ܩ����e�8��$d��FN�V��~Mi�l���K�Z�{]{K���`�Y1�c9N���7��e}@�p�K�$��۸0X��7� �(�=_�I�UX�"ᕔ^7L�L�^��w{p�oBMug*N��ޜ����ZRMaڴ�@\�ԃ��	�"O��8LG�&4}<O��4���\��
�\@��am�S��g`�x%U�r���+��|#v�;��w�m~V���E��G�L�����6Zɮ��#��u�3`�]EO��#E�)� �%�xf�n9�P��
ꉶ��cpǶ}��B+ˀ��'�P����4J�U�c��NO��,���_s1���'J���3s�]�F�`zW� 6%����pk��Y�sx���L�Զ��K�ewV��ǟ�C��2;�z;�r�dӉ�a]��u�� ��
>p��6�/��4�S��H�{����U|,r9�q��J��  �(ڧ��v�ɻX���i��^ a�Y�\�2��Qa��{�ʬ�W�j�1�E�-4�st>&E*�^ ���A�����ҸT��~-�UNd0qH%ZDI�����:>̚�����?Q$�mc��[q��ǫ/!6��㥗��3��A��Y�VX!��4���}��d�ܠ��рuZ;ɒ�R<�=�4x��1���2R���H��;F��N�r� !Ы����Z��y��y��:Ar�Adf�X��e�F���Ӡ��'������}�����3d����;��इ$�Eg�����eD���4�H7rUG��Pg��8}�l��ԍP���(28a����#B~*��ԦO˅ݮ㦉wD�x�K��Ҫ{�qPIB�~������q��U������1$�J�*�dQ�S`�FFk7D��� \	�d�0�(�77x�����|Gh�:#�A�h1/\o;�j�3G���<c�sPo����3羉)ڼ��φi��0��yz6�3/�����w�C�TH�7��#¼��)QT�Q����&<$��[�j?�n<z�3�G���CS���I�k��B?�^���4)���J��_B6�i=�蔯=qY簗�0>
&ݸ8>�<��\'qK�&f�L�筭���M��8�|Do$<a
U� 8\��W{��x1�r���J��wG
�����]�J^��ɪU3"�w�U.���;[�]X#ܛ�ش�|���~��7