��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����۳�w>��Q*+��D����?��Df���{{J�����o��'�_Ybq�}��>q3H�3(��=��3KKY&&Y�4��rw�>!1�5]�>�1���Wm �	CDg���VZo��s0�y��P�����Y-�4�,~p��4:��n���4Fͥ�1Z�tQs��Y6��	��s�����h�/��M_���}��O�UR�'$j��B+�,��fi;��y��z�P���2Cq���k���D�8�`��ʐr!T)΂��HH#��_G��[NK=�a����ic���4�NP��熈n��,&�6Ip�_���@�v�Qz~g�$�����)��^��V9{W�9��9E�>8���&������,_}��j(U"n)��8�e���m�V�>�O���Y,�r���vW��u��xڛ.G��k�˾�oY�IG�u�q��j��}�+E^wc�6^��e��������X���_'?��GB<��W4(����#Dp@M���U(�j�ꩥ����痫w�X!&,\[�w�ɓ�߁�[	s�!�(�����aQG~99�'������#	���&e�n}��i�B���jf�T�6?#=�fWT~�!l'C1�|c�ồ��!|�x�����q��?c���FiP-/o�n+L;�xdQ5O�t�%K����z�aޢ��T&0-噖�1`���o��$a�K�#J�g���X��Z[Py�D���-�^�^���Z�S��A���u���y��i�"���r3:��O���N�(��j������0$�l(��m�C��Oa��������?e���k��q���3j�,B$���J�76P�=��A�\Z齿�k9�~��k�9X����Z|�b�Sa�>'��d׮�͜4l�镧HN�D�|�o����	��l��O�h+���6�����]خZ�Ӯۜ��k��z����+�y?�Z��?6�{.�2 ��G.���C{�F�Z;[򼂋�Z�5/�<�M�.��du^z_D7D��~�*�_:��a�G~�G��}آ"�z��L�s62`��RT�d�O���XSP1�-EZ�\T�Q��?<:�����|�n��5G;��?ʭ�%�֑+U�7�����SFd����[_�^��Ɓ�'&s����{��i� rυ��P��ˑ�s���J:e弹O�X�!�Hap�p������ׅ�����&���a��u.�Ѹ�6Y�8(��V5�xǵ�� ���/�M�S�搎̦�RQ�� �۹hb�F_�5C^�g\�$�n�0����Yu�g�Š��7>lI�	������F�h8��WkF,7�|V��%�I��[�_L�뫇S`l�5zx`s��p�g@B\ˑ%/Χ���ȀS�/ox�,G���oQ��!�����8+˔���\Ga�����,��"��ޙ�MjF�8���@�Xh�e�&bUI��q��jN���;�n���St����^��6�F�R��Ƚ�tݣ�򏪮Y�Nȭ��o;�/�I�v�k=�<?��N�?���R��Y#�%�.`��?��]��'����2qid��q�ȠR��Kub\c���s¯	j�<`S�a��,:Z!�v�:A���L�������l�����,}ھ�楡�	��gxdn=�@>���68�l�`0�FC�1��X��%7����'��4�׶���Q#��'�S":��edQ�����
�C\���ٯo�U��i�h'�ũ�c@z�<�=.S��惪Lwr�>�~"iB9$ђb�b�Iaς}�J�����س��Y�(�im����˨�5�&�(��yY��7wU-e���8�����6.��ʆ�gp�o�nH����I�7h�9�&�дX�@�~��D/�;fZU�	-��e>����y������W