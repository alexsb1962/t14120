��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^��������0�G���XYs�s�.;C���m��JW���mx*	UR8�R@0�v`SN/_k���J�/zza���w�T2홈9^�2�̆�ah,�!��]�曰�83l��tt�]��;�T�k�m�{.���S)?a)xf�h�:��C����2	1}�1M�84���cѐ�c��ܱ�T6��LF ]f�@�p��טB����)0��l8<΅Sf?V�Z:U�e���l���g|��W"/:Wΰ֎���c#�Dl5t55���'����6�LG�t��aì�\�-���6KF=�{��B��&^����ˌ��dq��8=�?���ƪ�0�n �t�2������{�x��閷�r�p%d�d�O�UXy�s,��Q�~�܁�va��ǸW��|a!�b��F�OHo�E'����5m� q�4�˵0����������E [�z|�P�&o�9����܎�}�#:�B����J��N���/��������O�c�av�p6�?�,NBνcH}p
[9��;
ab=��xvmca<ψ��C��:���7OA�V!o��]r$��3��:h�j�$������r�6F�9�"+)��2;zd�<�0y���3��!�A�bS���H�l�M�x�%�Oɯ0��H�:��0��i�aL��#e�1���M��6ttLcE	�Ik�~W�����@���m�I�E�ͧ{�
����PP(Ё����e�M��SC�g���$@Ą���og\�����I-V�<���z��V�������P�3���l�A�<��w\�����hA�c����0׺�E�.���{�vzJ����6��*8�#�S�ۍv�N���]��Bp�g
;�FC+O���Ѹ���$C�p)�y�Q#d�^Q ����7<�,�O��O�d^�7��'j��ć_7K H��s�^��q*���`E2Y^M���H�+���^U��O�G�ͧ}Yu�jܯ;uxq+���H"�%�#��4@AhI�t�(��㒻m<Rۼ]!����/6�tiĶ���8�^5ķy����$с;↎/b�K���M�^�hA!�Nf*<	a��B ��p���/�Q�p�ƨs#�:�3p|���sʮź���c��wJo�/��vzB�5���.nI����3A�b!;> ׋?���9.܂��%��`��S��"b�Xn���� O(���Ր�vH{�͠	�R���:����vKr��JC���z�'.�pV?І��a�Q��+��wd�9W��u�Ҷ� `�,֞�L�ѣ+�O��>Ұ'�c$
�	�r�&U|F.��z����9v`J�{��,�bVݷ�*�;E�ε@	���e�k=72'K���D��s #$\�Ӥ6�x�R��+��;�\����"�H��p�b�d]͐/�p_Uw.E�%�w27��r����Pj��$sr��f�������\�<)g���
q�c�SM�о��˂)�R)Q`���Y�T�ټ-kc��I�கWk��ȝ����N�^oy3ܷ�^�|��N$�g��A3�p���"q�W78��z���J� ��p2*~3W��k���0�JP�G?��P��shta�g�fٴ��:��*�f�+\_F�G,�A��B������s�?�ϳWx�G��K)30&�mjY_�6y����@Q+'��C�	ϫ�[�����C~[���,x�mU0\lm ��I<|p6ahu�/�.]��&'�ֳ�! ���yR��������Y�Vr��s}�#|c����}�riڟ4���1�u�g����K�gBvy~**$��`�35e�\�6��Q��f��ľ%�q&���!T,�W�R��We9�0E��Yg�6���3��o�r.�­Q��������Ä���7�
�͹H� �x&J�#�B+��@`»�
2_�%�n�X��5��=x�=�Ɇ���XH�~��d������~
��U>@�DG� �K�<�'��0_��iMb����o�^� ,)�� ��0���{�~��j��m�!M4�?:镾Ȱe�ci2K��E��UU�]����,�������~]|�`�U'vi�3��ρ�=6���	-&-�
��Z?:�	ߩ�h�w��J�ƈX �Q��"�,��ι��^E�H��Z��\L���4_J�c���Ė�b>�J�33Ց���� ��p��c1OI����(��rG�x����w���?N�u���2[�3�a'ۻ�^��bz-�p���1f�� �k�#��&���3���!47E�9�ʁ�5"��7������S�Y�cv�Z���W�Q.����p1��aqq�Ղ��� w�)�&=T2�U�� Lܞ<(�=���XS9t��;�s���4bU�;l�) �m�����`\���7 ��Z�_*��K����p�	���k��)��1Qp��'��y�&g���)��&D����~C�KT��8Q�p����|�FkC\c�gb)�DRǊ�_�����.�f�J�p�����T{�����i�1q:o=�
�q�n���<��eJ�w׳�����'���1�3� �y�4/?�8�ñfU]D[B� ���r�f�)�u��+�ۈp��ϱ��Lam�,�߄�ٙg�g��~���t���-ܿ���gF�g�r��]9Ks��g"���j��b���Y���y���=ޭ.��밈9+�r����6L���c���s7�b���l��<|L>�=���Dɡ��̠Ĝ������I<����q���}��A��vV�����Wh�˳GS�XF3#��2�B[����p|b�@�iE�����#���p���	Ź�/�q��N��b�h�	���`�k�B�@�GN�Y������9��գ��=	��x�/[���Cޛo啍qc`�i5id��Jpo07ZR�!��|��S�!Ӣn���S!T����g���.	�a�`�U��R��&p �{�o��"sq<\��l�m]ɟBz5��ʜ/�F�[n2/A�TL�f|�+���h��N�X�3�%bk*<�r&�+gK�^M�;�T,��lz�?��3S��hM��Ln�r��f3��I�eȦ𖸗W�ǎc�3���1�!�88	R4_@l����p�(`~�5�P�=�������8��p��Κ�6�l">/`ے����ߒ�����E��.�CQ�z��99}7�AP�F�W�3���?�)�!4��F�`O�׍��69���)�B�QĒ��snYcH�|Ú""J#=�|�2=��7����/��s�"�K��M�ZΒg��Lc�l��λ�כPğV�dk՛gJe��M�=�]2n9��N�]`ci5�� ��T	G�>�E��L�H�c���&��"�\0􏵻��d}�}��u��PZbg?%sR%��.�������W>[J���Mb���`�]! j��������>�a?�����ƒ�ޜ�1l���OL&�� O8�-�Y�6(���4�H9�^�7�_�x�N��M
���Aܻ�7��Q��B☝��X�N������x-�[�ʋ���n}��.������ � ;�X�F�q�~u�8��ӷU���u�д�D���:H�ëX��X����8��M�: ӹ�^�&�Cv|
��O�*����]��t�	��U��(u�z�;�(�:�'�F�T��@o�+=v�Cb�?:]�(��,�H��D%���x�e�����"s���9
N��|n�N���.0��;&���*e�qϓ�y�����@Q�~�mD�=y<'��݉G�'Y�YYw��(k�6�~1$�j��.b���K�����=��U��/t�f;��˒I�D���%G����ϐ�?���0M��ݞ><�7�G5^�#v�%�Lj�/���?%,UZ�NL���f�����*>�r���.���n�kcĺ�V�����M�(2����U�J��mh���j��*v�B�%����~���0RL��1�-?M��\���!��m�GdR?��J��o�U���oJ$���,�B�@)`������#�{��R��$8�ʴH���_�"���E�g S�|!M�_(��273���˙3����UV����	���'��ٍ���;�)y�Օ�ց?e:[V���`x �vd�.o��[��3Ʋ�]��9�����L�0�N�I��n->z�+K��+v��a ����]�KI;�%�Ya�	d��/�ZTi|��8��W"eUx�A�?^�z=�Yi�I��� A'`��,`#���_L������g`�#��H���<�vA�i0
��8���2��v�Ea�o��ϩ���V��eϫ���x� �S�9W�g+������wD%�~__[�>�oMvo��(�?��t��j)��)L�f\���X8����z�Hҝ �Q�����6�IM�X1�5�Y�����c+�%bCgX�D*-����~�)&���㹒�ؘ�Y֍�ձ��	��Kk|&���v+0N����E�"&��K%h�V�f��@#x��o��P%�$U�9�Tz�t��΢�Y��gZ�q�I�����s;��j̡)⦞���`���y�ow���2�8�	k���&�RYLB�Id{]
yoQ�(E���t��䟦@�@�i0M���.�i�.�].��g��\i^�;k�h���;��
/+�X��>�xf�g��ev`�cz]����[�w�BUP煕ę�ïeD���&K��t��VE]�j�R�@K�������=�J�F�'^��E@C�!o���������>���� �IuW����U�Wjw�Pq�{����Ϫ_�|��x|��\5ƥRGѬWةj&��](8f̪(�ra��������{Ot�bY˞yj����n�Ք����&�1�
e��l�B��1Q��u�{�os��š�9���`s*K���G�e�m�
���|�u� łҿG��t�u��}8<p�*��
�J�}t�p4F� ��!'w7?<zF�O!���M͐��M�p`2p����%���n����?���B�B���
K��X�N8.3~���4I�Q�ۍ��eT�pn�j#.v��+u�kI�?��%��̦4R��#f@DC�B��A�m��K���խ�����#���^��_
���C\WXyJ�`)�=�y�~���Bh�y�|�[������k�}\mo~_׮=Ob�¹��`Q��)48
�`�.�m�dO�⯢���C0B�a�}�Q�'	�|��W���:���Lbb����������땊�M�k��^�u�V�<�s�����lk�j���g�=�x�D��g��,�Ȼ�cʹ��w<��*�2;�:�A~�&��9{Q!|d���
럑9PIZ��v4>g�/��x�AP��S�W�prK��Mo:\`�}6x�%�(���&��^��gR�[�Ⱥ�9����uFp64Y����oQsGz�Fo��ض��^���V	vzq�Ys�L4H�s�	ۚ��7�D��y�T��j�q�Î�\m�)FH��1V��uEh�x��I�5f��N4@h���_�L3�%-OQ����6�A͍6��ד\��J/ꍅr>�ד���	��=䨶rH�{����I���{-��.O��W�`�O*]�@�����C� \E�Q��s�+�n(��/r(�8v�"NZ>D������}�^E�����s��P�hbB�=:�e��h�����;�詹n��'�|��|M��&Ն���lX2v�*²]H3�ߒC �o�������5�>*ո�t�������>N�sZ�� ��J�]F�`��)]� 9ͮ��}�|�����D�b� �;� Fr�N��x>��-!�����`$&P4k]�>I<��GW`�c��m^�[:<<Aj��^9o���ս�Z�$�ڞZkҲ�3�<m���c�
J/�C�G��Q�۬%�w�
�W|&7�+��'HpI!]��_�Ӟ �pn�9�窤Mi����t�!)�����ZX�P3ά�w�H-8p�A�N<����r�;fnh�\, f}_l����u�'�Xz���!�f)�G�.�T�^�,Y��_a��ZV\Ih>��W:U���ls9�Bf� �|5KB\�J�������V���b<��}��Z]��j�z�
ӵ1�X�*gl�<�l��l �J�w��+�Pj��@*�qө4T��$ɛ����=��kHv�SB�����!J���̎��M��;�u�*E�T�e+�P�����x��!�V=bfacA�Ao����f�\���3j�<�A99:A��%ܬ~٣�����Ï-�wt�#-:!՛�����gi�)�ҏ[�r}
�����ܣ�ǐ�(#��`�%-PuM�>H\@�r
.�g��''��Ң��o�˸l9����:Mo���
��ZK%�b���V6����&�̬�ɞ����۳��׍��Y9\���gx��ar�����d�|��M�~ɑ*fV�f����S�kR��}�e/�ܝ�z��P�f~�X�3֒O*)D�7�GBql"��͔� i.��c�Y�U��`ڞ�$�p��3/�Su{�AwM(�CS�v�=S}���mt`�􉳢�o��1R�M��z������%�C<=^�o� ��l���'/첫ϳ�e�����k�BS�3��xnE��A����R�᝻W}�K��W�C�4L:�Dܚ���YQm.�s�؍�c O��7fW�v&gp-��	�� yiі��O���8�
3� u�`=,c:�^�%�&S�o�
	5������;�C	���n�6�L>����X"��ڗ���{�g�i���2:�)"�fxf����PQá��?_�2�CS�m9�c�.	U����V��@F[l���`�0SP��<���cs/ d��'!;��~A��B�3�|��C<�]Qn���CO+3oW˞�F�.�x��;G��ח"�͍ X,t�ƤΤ��0��h�����Ae4q�`X��}���t*����6V�|�YC?��+�+o�n!�9w�Pp�M\̹_�J\��AdM	�G1��S�1�b2A �K�tt��C�,�" �(&��ɨ�}��D���oK1�sR�hMA�m[��t1@�А����a�R���~� '�e"�UO+��Z{���a��'g{v�(AV<O��	:0g?uR���FB0�3����X�d8�0�##�S��M8�aPn�h ��Z�����
���s����eibA�끄�)�}c�����.�'s�"��_B|<�(2������J;����N�y>u�LEWNi"�s]ݗ�!�}b�-[�TC���@��]vX�rM���R�q$
��.��_����׶6��^� �Y��4K�d��š�6e��6>(��Bij9;�ؑD�;T������Q��h�i�=�?ajD{��x���ڤ��dac<i��!��)�cVQ��X�|�����������~7�<~ڇ�_"*��eS�b*��Ð���&�	�����/oS�4.h
��,Q��)��P�h����.�w5�U�󓣜�nv�T��u/c�mx�YVDי*������p5����u����Ma�rO�S�'��5Q�R є�/T���Iw�晜	 "�\�&�&_M�ķ�ȁ6RZ��ʬ+��<X�j���t帢��Ƚ�aw�G�l.�,~���A��SB ���d����k��#M��1�B�����z~����B�Ø�	��%�Cή~e� (%	��L�UI,���=l�	�["s����E�D]�9��y4����{��Zٲ�|�Y����q�9ǚA�]�ؑ���κ��i��2���W�h�`z]r�������gٹI�V���L�������
���W���NK���]��u���b��F�t��r���]\j��{�X�
��n�e�#�(�梄%����S	z�-P_�PG�N����܅7Ӿ�1؀/L��m Xȣ.�uŎ�&��|V�:����$!����u-�3����yCe�J��0��qY�����՟���J�r�ƅ.l�f�#pJ,)K��{I5Q�	jC�<H�ϛlJ�G�����nb�3�y�w$ŋ��:����u�'+6,������ ���-�J�9n
+����GU��;����u��G>K�;[�����֠x���`4�=���T��*h�1NA��y�_u@a�]��Z����FiU����=jjC��2�J=����=�*y���_��:�>g��vW.Ǯ�esIrE��G_���ݴ�������w�����f�k^��Td���GZ�
ĝ�sɽCݒt�b��D�:�C> fh�猖���D�ͪ�=z��;R�!�t��Pe��%�#��v��ʎ�
���M�![�	9M��)���Đ']��,!2��
_&'��u �1���4>"�}��
���7g���Y\�U0i�I��IU�b��-�'J��@QŴ���Wzgj4ȘG�;��)	��ְ��u�C��Tuq���9N�7u����D�Mz���S�}FaLv*����)��r����2�P�}�r�KQ=eo�u!Y�w�ߚ����Vn��^�|����B4�x(��7޼����C�D����
�q���]|�;Iؐ�H�N��Κ#��O�0��/ξu�@9o���v)��>$��~��@���?Ԅ-�٨��L���1/���㜧�\6��kl�up2�������'���t�"F��"FV�oR�i��B���WaB3@d�՚�5����ϙ�٢8���hN����nWH|�^�����%�b[�2Q�\�;p(æ��|-��D�\�^� R��|��`+CWק�GK5}M������|�L.b�lYps(��]+����r�E�ۛ_Œݲ�71	���Q�jy�J��n�1+�Ϧ~J|�ur�{d�^�{6ŧ}*����X9�|���]l����3�K�>>g���|kG�ӏ�x�990�-��q^��[a��	]ȯ)�%?��b��!ܤA�oP%K�ݘ�A� ���M�?�PK����z�s�|4�x�L��Ud�]�h� 8��R�����k.b������6N"@?�PX��T����lC	�4�?�)#H� r'���q�cג0)M��r��X��s�\R@k�4Ňr��R��ₑO �D��]�+k�a�c��_��nP�;�C�Erѱ�P@͢a3���Ye
��s}� J�3>�NCkB��	��;��K �}4��^���u�k�qeՖ�S�g�!P;1�@m>����y���f�����z	6�!���\9�D��a�D�H]�$����u����+�6��fE�.��x��Ͱ���N�߅���Q:2��L�YٙԤ�J���˓��oh1��]ͥ@�����	�B�:y�����ba5�Ry"x_�/w׊_�z�^��{4�mI��BN�4��[B��= ����6��L�3�NC��	��j��ٵ-�2,� �\@5�*��.��il�JWY��P�؟%^�bȤ����^&�o��E?Tl^t���O�Cu�
�\�b���~ HC�����+n&�]�LT�3�N���+����:�j��Z��Fآ�]@��hHaE%o��/���T�;7ABC�y�b�_qk������;����}��y���/�R�y��'�2z�rݪMNKΠ�[�O�zH׌C��'u����(+�B������X���C{ ¢�� h���'�G�IMC[�/��=��JX�9��|q�Ƨ0b2�ztW\����kb[F���������Z̖q �w�M�J"���B���XL]�B址�>E�L��]����� �e�x:4�g�v:ۇ�<����ݤ���p	��l&v��m����Ҩ�g�0�_K����Ms���WҢ����q�Nnv���g}ȫ���2��q���
�e�q�kf�w��ň=��K��J�Ϫ>}h=��<����'��u>ㆰ���y*��p��:��;�0q��U��}k�uaSI���
n��0����S^����j���ֈ�dal��y�+�!�����Ӿ�6�e�"|���))��/�dD>'V�N�'��e��2HHj⟑[���J �r`���U���},�q=�
@��υ�4_u��)g$~%p8�&�����_r9��8�`�96)�K�T�9�%��4Ҵ�ѯ�Ҵw0��4��t���!�������%.����]݃�_��-:&8b������2�%q��ш5p$ͣ˘D/O��� Q=�_̜�JW8B��r3�vzf��6+�˳bzc���Z��F��\�R�3��kb�a�����nt�_Ƚ�#����c'��`�５���� h<%�1JLUЄ������n=�0��<f_?I�ة�e���]�C덈U��H��;rD�����n_�1��Ű�dćl��N�����(��}��v����F�}�|u�`��������Y�"'����*�i	����P!��.��g�'�LZ��jBn����&�����s
���őb�+�s�
0�6�>�����IqD8�Չ����1k� ���I*�zp� �_�I8?�e����Γ
��CeDQ_F�����r�;�B�h��M+2��%Bt7찋�2��ݷh-��v?/9\H�&�y-���>I�<[����򒼮=4#5Z�3�N�]�(��֚mw�D3��f.CI�Ģ\��?�y؟)�K���,��Y� =���W�7����pO����gD�&n��R�����U/l�����oU��\`rb߀�A�L�o.$��n~�����P�"]�X�\r&V{�{L?2�'�j3�iM�d�\��7��j�W�-��K4�*N�J�*��Ȼ�B���z\���y�1�G[?cQ�Ж�q8_���)tV}����\g2�P��_:ŀ��/sQX�P�},?]dh�L�~S����v&�����q��B-���f=���[�TB<u�_/�b��L�؉����T<B<@)�� �y����Hс�����>��Qo�1�z�3�2���'#�ޑUg�Č�+�G2���P ��՟ج �b[ȷ��ASR�:��ry�\��ݗP?<�C�.��#��3�XrC�INr�/�� ��Q�;�ʉ�x�� �X�]A�*��< u��z��Q�����տe|�	_a�~���.���Ǌ]��<j�ݙ�C��/b��<$Fߗ���������Q���2�o��RF�W�`W6Wi����D��wR�w�A��S�� ߉��k�����ވ@Z�]��=��躡��_U���$]�����{.��r2Ȉ?��=�qe<��UK�I�����-����YۀP��;��%GѠhH)P�R7u�x_/C%���Ms���KZ�
o��q��)Z�	I(��I�Ҽ}�O�u���Q�q[L�_D��iJ�wQ�9���9���9�ꌵֽy��:{�%��2z�?U�HZ�KÈ�^[�����r����BB�h�C(q�{�����5;��	Y8/Ũ������T�2�1ROv�1��mۻ��[���%���ʾ�C^��=�j����q��o��b"+Rߝ�P^ic����Y����]�=H�5O<z��i�\S5�*����ـ�~1!	g�Fn,�1lB�ٴ5�F�|��@F�N|��K�_{۳�R��P�l�\�l���I[O��sm��N]�y�9lA,0�=d��qaJ ��$��F�d�=�����J�h����$��+�j�7)Hp^�f�?X$m8�1@Nf�u.çT���vY��Rm`+n�%�^�礪�T$k�x�\��vL��d����K��~	Ljp�[NҰ1�͆��,�鴰FÊz���OO�$`��MGy
�V^�;��{QCơC�Ώ����C�����Z�5�����!�ql`��o�4r[|�/h&�)D&d?�.c�Bl���������&�>�ο�9i|��*'|\��%4�-�X�
�.�������ϋ�*�h�B���P��r�FJ>x�k�&��*� *yp��6��Дʨ����о��\3�z� �ZE*�F�\��D�}�?�B�|�5�Ev��LQ��Z�� �N��������刊��?��o�d
��e�ѷ�BEZ.�ӳ�ȴ�h�k`�J��>l��
���2��ru���K��4S�=�=�5`�W�ev���z�E�	?��9�-�[���E��	&sw�eؘ׍� H�Z�<�&v#e>v���y�6)�r���t�� ��ݳ^�v�Z3ԉQ.E���{%'SRZPbu5����S�lf7��NE_���}���@�iG��l��Ӓ�>�g/S ��i�)�W��ݗs�sV�R�
s���;$�G��4��(����ڋ�V\^P=�:�^I��U`i��2U$ɐ�b�Y���s���݊z�fP12J�uB�����*��.����x*�X\k6��/)�e5�	����$U���T,�B�����a_��O�^P%-۽/\&Q�~����}3���/w�q�%��؃W���,�SM\⊄�nvٔ.�E��-|\ē�Є*%�&�i��Է��U�οQ8y?w�@"�H4��^���������c��5�;�87�9'��:��5�N�8X;3���,"	�)+BN;_����������P	�,�['!V�,�,��6��gg��%�A�d�*S��ChωP�kN&19gQ�\�S�F����#�`���.�I�4d� zJ���=�'��aFhً��4�7χ5N����SN���h�)��|�2�I�,�gOc��bz�)�jm�N��%�3�j8���� TۻG&E���~]C���ϸ���:Vmn�@bo�n��^�pӟ�q+F�wє��δ0�MÂ�?<BxA]���ٯC8x6x��HMHW�_/L����TN�$y���5=�)��R���?\}�?�x�1�u��@z|��� 'F3��:�|��y�߈b���86�[�E�u��R�c'w"�MV��a�7�z����*J��{����� #��?�/_5�e�?��#>U����5����Y��F��T?3t@���-˴(�o0�/�[�����Ssw�T5c�����{��x;�~A|�S͜���uci�-�Ex���,HWRq� Ԙ/˫���d��M�RU!*q��5�ەI|��$�!���kI��?f���mலP�O�
�H`�kUG��
�_�S�R��� 3/�)��CkM��g���R�i&h'�J�vw��+' |��H#ym�>��uM����&$%��"z��d�>\��PW�>.t.�A9���-7ݱX$.��[�*�C3�p��]�Z��1 �k���]R�j�x�3��Hd C��k/s𩬞��s�Z�*P'�et�|�!DH!Α����x{�$.�� wTE��{�����;s)S�{̍"ġ��%q�i��о���}X��{I	ml�9����{=�w�T��a��i�S�����U����O}�]hMY�q7�����ga�nn��ax���r�r�d43��!�uޠ_(�B�ѷ'8~�Wd��p̃�y6���߼��l�����J~�
?5�a,f!���Nb?y٦�ӿ����<����<=h��Um�8)-��B8�U~��wUL��[���(ޣ�-����Ԯ|9��6Ν۲�7��o�4#� ��@�-����"�/�~W�H>a8?�;�tIZ�=J�0p��tW'׻��z~)�1j&�IL�����v`k����>:���f*n�CF��^�
J{)凉�m�@�RtnBm1gb#�몄��P:u<}�%;U�r`9&C
O%r4X8����r��5��a�<� �꺏��Q�s5��>
C�����7��7��j�?SPz��\�v��9r��Sš�5���X�G�%��K�?Sr�]�k�$s���zMz1��S#������w���#�r��*�ک����o���
9�a���� ����q�4\�+��A�*AN��#��N[����i��$_�ɲ�#���ϊ%�Vo��c/R�3���L 3������;�~]$�G�1t.����6O l�U�p�i�@<�" ;�%`W�]J]�#?=v��QmOsq0=U1����ޕ����W�k>s%���K@H�0�\����h�27s�#X{�������nÓ��A���a?j=j�W��ow�>�7U�G���4���:������4Kv�"�r��P��)]q@Og�t�KR� ��C28�H��g��9}Y�L/�&u�Q�} �C@����c��Ա�$2H�" ��=:��7���ó_�u%���?�5�P�@a�f�%Ó������=�+?e�=x���F�8��Dڨ0<�)�jZ�c�{�'Ĝ`�0|�	GNcA��=�:�}��5�
0���``P�L���@Pc�~�:ݨˑX�V�����	�G�9���#b��E���~BBD�����Z�Ϭ�n�{����t]��;�����v��}�g����Ʈh]��o���<7܂w#/�0�ן�݅�9��N*S��S���J�F�v�\/u���pzb�Z-N�r��m
Yd�oƈ�='�S�yV�H�˰�y�R������)%@~�"����5�ؤ�ſ��g�6s]��o(o� +�6�s7��l�"]/�5 ad���梞D��CI���[Ç�31J[�����+h�lf2�e=Xu����o�~�џπ!8Ǹh8�|#0�Y�a��s*��/U�� taa����Y���=2��Cz$�5�	Nac`��OE�� ��Us����,	�@�վ�ﵯ��
�=!qO�pF�Xi��&�*�7�]H`�ǰ��V��"؎5#�*=�L�`X�2�Y+S���f��&C�U8�\���e�I����BϤ��}:+T�u$�X�q��q!��r0�N�0A�c��g�7_�=r7��P�4:�8�i��CP3�MfRJ�ca:\�|y�-�x���	�Ca���_��Q��n$F(:��3?���?L�[����CKO�X�Ë,	���托��N��%r�%D��`#V��5g���h����B���E)�G��ހpx����0��$Z���!��	�.�th��Sh����u���������o��yc:x|/�ah��$+�3�αOX�=$�~Rw���G�"�֣�G3fk�����4��墜�.�(ה�+m�64ڙX��d���$�c3�3�X(���:�(�/pF^����2u���!s3]8�&
�Xr�H�����f+�?�t��˔����זh6�Bk[n��6k�)$B�9��ݧt���t=#}8I�H��@|1v9�o��n����m��\
�I�S��>]#}�e�:��ǴD�����E@�@h0�Ic�F�IR���J���l��%p�G��.��l؞��"E� maQ�d�����L�hT92׏ϝ�p���B�PB0ѥ�;g~��E fW��Ʉv=�$h�m��7�>e��p��!�~�k��ҏw%��</�v	 �����뤇llw1Ԋ����s��h�J�d/'�o{6�_3�%�p�ѳ~��/Aاm,X��ȼ��.�5RaM�U�W��`�!�>mV�^��#�ma���5
4�e� ���g��O ����i�J�[jm+]1
�%'�pN���-Lb�|Ȉ�Z�0.�e�s8�g"H?|��K �H����m�vg�t�����������#��pB��n���DW(����b��`���!��@	ٚ��j���!�{��l�Z72����Fk1�T��w��g����{5�������/��9����N�W�����V�`B��W;��g���^�Q��P�������3�����Le�<q�=���>4>,�/���%�����@:�=��q�\�����M,[,�Ӈ�ﭦ@?�9���!,H=���?�ïp!�Q��������,��Z�.��Y����|I8���c�{`�h���!Z&{fT�;�w˭D�fLV63y����;�eRP�U u��{x�h�-j���	9�8�*_�`��� �z�!TV�|<�E�+��"�塆E=���4�k��Q̼=��9�����k#��!�!1�]����2�;J���p��1���,�a�=�|�*����=l�TFJ�S
%�h�R0I�<'�v;�r=)�(��|�u��ώ����D��Zl��=s8�ZO����D�G���I�&��;�A���Ǝz��G@|�z��:���s׿���){�Y�ol��;ۧ��Ru#B�������Ŭ�1/X���IQ�[�(K����o�ԭЌAӻL���qH���`�@`���b��"ɞ�i�0��Ӝ�,��$;S;#pV�}PA`�>�L&��@0:���3(lz=(����)� �)�{���������Z5[2W[���5!\�L����M�i��R�SU����J��H	V���B	x�布�BM*C�mxs�]u�	��q/e����uZ䥕bɊ�����4�*h�O��V��=Y#<��������7ػ�rx-ӭLL<s�Bi��@�7��#Cϫr���q;%�^D�**�Wbn;����ܐ�tbР^��k��YzV��YN=�3�C���`R�m��R&(M�����[��q[���1�r�\Do���s�Nw�7�cc��{�� i� _bm���D���V�<�m�\�E�vP�b~�	�{U��c��Iy1�Q����+r�@�5P��Y�����F7�N�j��x�J!&�ʃ�]�[��'�|$skj�0m�i�d ���'�e4O $kO+	�t�Z{t�]�����/�ǌ�Bۄ�TGi.t����LAz?P-�6���sCe(a�z����� �.V(���N�6��.� [�O�D�MQ��rͿ���D��S�d@�A'��w}�OL{g�5���>�n�iXF�Me�������z|Ca����d���-�W�Zm<���oi��F|�v�f��?�j3�
���f�_��`�.� w9�\��)W� -�Vˡ��Fj���G4���PX��̻�߹�4x�.Z�e���:��$�o�H�8�d J�kU]���z���H�[���e-���7X����B���/����Izc����v�^{�$��Ŏp�R��s��ʀ�?�i��@/_�`��=RF���tJ���9w�y}�w�MS���b�x���p��ƨ� �\�D����W#w$q�\�({m��H�,*��+�vMSa�ѐ)�5A���p1�� v��FO�vѰ�C.]\��
Ogxi/���1ƾ^��_��V����1���NR6���Lf����r��;8(��c�^�õuђ}�B�<��������X�/��m~92�J��3��s��P%~��`fX`*Ȱpm
�~�ͯv�VGU��m����҄dX��M�˦}8yd�x��k�L�8�f��]MM�A.�!x.���«�QA��?���s���JCS���$E]����F0a�3��@��׺�A���^F�D�
�8ρ��	�<�57�� �Qq�/&Tz��ƫ�[�� �{d{���z�7�7w jdH�hpj,/�8n>Ŗ����.d�7�m����<7�S��X�r�`R�<6�i�X6pۡ��
�#tc�1�e�K�B�g+�0�{B;`E6�����EM������L��}�s������#~�\�='.u��BC)g���ރ�SC}���	�r��P��yrv��b}@����]FN����uQ����P�	�ѹjW���'�[�m��Qy�7��w9ª^�S/�j�C�_t��qL��3��P��ŭ���k�\��eM;�������Z���O�eS�?Ü�B�[��$B�B���u��"�YO!� C$��}xP[C�E��yq��O]��`�ǜ�R%�� q;��"�m�k<��9��O6S�O����v�M*�����5&�/w�$�ԉ��5@����}!쉋݅)Tk�N������4.������þ���@��qrP�:B6����{O.� �y�E�V�NrYc"�ۄ;k����^O��Sl�ew�K��Y�+b�a(�y�!5L��w^�8�&:�5��L��%��������PY�����)�y�G����i����D��{�Z_8�D��Ĩ���y���@a�c�ٖM��!�g0$Q )�#���갨h:�R�2�%��5�F�=(v�h���y^��Dq!DM���������g��r�����:G���xL^;�Gz����VS�d��<�8?�}OxD��rhvX�S��V��}fr!�h���`ܰ^�ø����H	�AL'�^βk�clt6�)SNfw����w4�4��^;��+5в�%ym6��O�������y4f���W"(-����D�#9=�v=#b⦁�˞Z�8�(��Yd����`�+li����/���la �z5/%A����EQ"{�����7�r����0��@��<���qO�T[��^���z�8��.��K.���
_E��.*^A4v�� #'����$ V�p�l���S�Q�|'��lJ���֕h���2\�y�\��`�J^+�nk'�o-�xt����ڧ�Cӭ�h��v��pWn�b�x��}�1�"[�������'��ާ	1�Z]͛A�������d�d����z��i�	�zj��.1� b�W(d�c��k�#���ok��y�H��Ȑ>�b�H�+m� ��ק�k�U������>��Z1,���U�69��k�,��u=���岼��i�(~�'JX��-�!�Tv�Dv��r��V��Y�nl� �$����p���37rc�^�%=JL�W)���#D���U�ɨ����\b�07���/�;�:w�K��|������W4 ����W�%j��F����F$gO�#tu=\��E�$������ze �\	���خ!�9�ێ�%�w�1�Ǚ���f_7����C5H�3s읉�_����m����`m��'%;}�ȩJ*���˯���L��3Q�s������v��,���y_1�����ː,�y���gHgt0�d�l����C��ɓ8e�n�}:�hVL�����E�`^�S��z�1���B�%8�����P8)s;�&ռ�|��!��a�EЎ�mɏ�G|����"n^�SpXA�hR�Z�i�@Gih�CVJM�է�FR_���S���+�h�B䓽]59k>,���Kr���.ʟ3��[e~�#Z<ǚʚW��]ס���p7K����*N��6(��s3���Z���;��b&�(u	W|ޡ��Ykf#-g�[�a[�?mb������=��dF<�a�5Ϡ̙��Y����ɒ�����H��e,	d]{�U�-o�u0��/^X��H�X9��a����Ǿ�S퉻�@���nO���ܥ��̖��,:Ta�9�|�9�}��D��o��8��T,G� r',�/H��Ai��l�	��QBg��`�#�eM��H�j�0��eZe�@�|Hd0�6pE���~q<���	��솥2��+iۄ���E��Gv�|I�p���v�I"!Sp&�ZG*���,�ػ\�y�Q��,�^6�:�Y~l���o9Nb�G�+s��:�8�w�f9߹���^"s��V쫦��)e�̑�A��������P�P�)�*( ��$��aȑX�H���P^���<}�=xӫ�j�>wQ%v�W� �5p�ވ�rF.1����Dw����&�M�=-�r��gw�,�����H��\���̜U qh}�˰�����
 Y� �&��R��,���|\ν
e;�!�ȟ�/ 6X�K�Zv0��զIf�*�tN"6��]3)��tl�{z�V�0(�"�� �^^*�d�B�)��Z�Y輌�ɟ�B��,����b3��N^��-�B�
���]Ͱn��� ��Ut�BU���3�d`��ãH0�=䄦Xl����A]�@1���'9���ĝ6�`~s�4��vp�Z���_ѐDRS1�5�v���6p��-��IߎйN�+�;���[F��1���s !��k]A�M�}�HD9:^憐�����=��՘��F��e���h�]7y��߇��}�?����|���i쮘��gN�~�?^�:o��u�~���P�	�.�	�n�^��8ϕ��AP�U
)�˜X$�i9�IW���r�%��G*�A�z��uܫ.��>���
NN1'xS���/*�W�/F���q���s�⟂ �w��o-���f�	b���I�x�E��5�xr�Q����Pǥ>EߦG�T�{)����>Q3��u�3@] �V�!ř�˫3�6H�X;g�_�L[����*,� ���Ya�u%<���R�)�<����w�]������"~8i�K�*�9��H�;n@�����Sh��(��|�S�}����v=�F����n�橠� Z�7�������!g' ���dU'�:1m���+9�V���s�B�̓`
%�TT���Zc�+ٷ;����(����5�-�1*�B�<��R��/�3w���(�
Dۡ�UV׶B֝m�Tǖ�k��]��.}�H�X6����mC�mv'�q"7�`�!��
@�\�Ӄ\�A�~�M��K���R��y�ͦ� ��w�*�FA���#����f��=L{r���_�1L��N�`�M�n,q�5T���2K"a0RX��3���~;g�)�
6��w���d�ŭ�ҶS�cz��m�r2��XY����Jl2`���:.���q��&1Ķ#__�s������v���x�UV2)��o��i��c4�7�.ȼ{�$�%��uY��<��"X�K�B�~ܤpw�F���U�s���{;������[֡��O^�Y��#����I�P�''VZշa��'��[����X\�>I^��*l�(�^�ǁ 86�V���Ϡ��8H�|#�思�������{���pu�2Ѓ����I/��H7���K�$�vlxGA|�a` �BeH]-V��TXt�A$�rX�_A�M��#Q���� r����[b�E���T�˒��m���Q�#�1 c��L(} ���[$�W0L*��k��J*���iZ��y�c���;� ���Ӏ��g�n�<r����]�J��&��S�c�[�K��EQCƇk������oK Z����ʡ b+*�b���L��?~\�Nz8آ+v
�p�]szQ�<H56�����Bh��0[�^ 1�]�e�JG����%�O1�>T_���74��^\�O��b��DM^�G�[W�s�h{��[ϙ���"��|�6�H����}yj�r��N'\|D�}nW�~�P~	&_��Kx����!
��9O�R#��S��x�Q(��(D&@���b*���X��F����G���H��Lu�^�K�s��҃�i�WhOV�:�!=9��������Þ0ж�$en�R,a �;�V��(44E�z�����GZqp&Sì@@�������o��,)�
�.Q#xT�r��z�-��N�6z�{-oh���a���kB���o�c���3s������"�3#�K����8��u�����]��� �+�jE�����v�D�Q�щ
����q�hg�������s1T/"�*�����@󵷮���;|���7`�L�f����ĝw#�����^����~����Nͽ�L�p�X$��<�O���Fd"�$6��M��
?�)X@J�J�Y����-������2iOc���Z!�8~����V]$Zr��������׉9Lߍ�s�za�(���C�MF2x%|8G�P�Ѿ����T�b�d�3M1����vό����[(nK�Q��
lϡ���8���s=8$��X4�4���*D8�L�,KC����;�9}�D�49dۗ�:��;3�EPJ�����V���H�Ǐ �*}<<*1;�� v�[��?+E`�"^��WN;.ϝ},�X�Vu�	�P薵��m�p�a���4ަ�B��H�ݾ�l/ë�GA^��6�s�͆���پT˘����QI���x��p�9�mI	/���Úң�	Q�(��5�����oaW�Xw���D�n�����F�	r�6��:Q��9T�7��րp\P�ڡ�ܢ�Z�
��3��ZA_�f���a���u��y��OĜ��}u9��H�	ٌ�`R�-B�T��T��������d�SDp���������&����󝽟Ӌ�o�/s9H�M�*�/\�u�5���5vO+2����K�&��F�}�����f�� ��G��{Xw��� �2)��f���*׵/y��n����%Y������?+Cn����2*�+�?A��g,_�0������'Y��}�x�QQ#��O	�CHy�5��ß��wX�y%>�V��yd����V��_�0o񇮍��$�m]��z{�C��K_���ݭ��=f|�=�{�Ak����@߶�R�t-=`%B�X�bk��EW�� s�4|}�>ȚTB����b<,�m�K'�!%�:��c��(���~>��`K��i\�]U�����Q]���R�jC�X⿻{��)��"ǳwȸ���wk	f�+D"��b��R������VA���+��nU�3�u
����А�98}� ϗ�}�a�sީ����ڧ�n�e�G\��5�^�eboC�>��q+Td�U�G����/�B�<��ȵ-]"bm�.���qe%�M�G���(�>�$�!;]�}���̟��ݘ�.��e�9|K|Kpz�9�ƛx�r�X�?݊ᒛX$n�(1Z9���@c�d�tY_E鯈�(� �fO`���8�7#9d~���!��KƏ��d��9�n2vK��%�v�Tʁ�z��y����K���H�����y��d3�qr{�ZBU5�C1b���?�Qz��:�m���<�O�� n�(�]f�[��Ϧ�	��~}R��#gC�w�i��w32G8:���|\+�-Hd�`D~�2�+��:�^N���t����8̂@ �JIBz��7,����CgΑ�k�>+h�+���d�y�$�6������ ����z��z���&�� A4)�sU���;�%(�TO��Y6�Fd?��~כ�h	+��:.Ż��x��W���+q�����SS�qBq]`&? ��G�|e�v���;�ʓ���	���`[����~�� ]����m�##u/��l �-��*�6�F�2m�����.< �����w'
W������%��!�~U��=~�l�3jg_x��谧�
���Muzy�,���<���bM�2�u���L�'��%���wF�E%ͅ���:�[�A���nI�����/E�兝޽V��U�K��W���aC#�;j�B�Z�yI\�s���<��2ߌQ���]U�
<
|6��sLm�XE9#+l0�p����p2�t:pbp"�HC˾�*Y�S�Q¥�c���}h-��Qo]��L�9�Y6�e7w%dZeQfg��/�-�꜑RAz�h�ѷ��t�-� կ��툥i��@?�z���v�����|f����4�2'es
���6;��!E(�F�Badtpl�#�����N�C�*�,�jv+��FEU�Fe�T���̥R��˖�uWK~7�W�����v�S}nɠڡTO���Ϧ[`��N9���������A�RQZ4ߍ<�����R�~M1�����UI���#i3
�X#��w�8��C]ןڃ����Q� a+T���Xf�/����'�\��_l+�:f<���r"pkۛ�nz�q>z1Б���t���;�O�ky}���c�c0��x��	���n���p�.�{���pp0�GH�a�\��s@N�4������QS�V`�sd��1�W�Ubw @QD�ult���;����"ڸz�%}����W"8D̃ΩA&"���� t b��T��b0�%M_�B4|>u�2�$;I�-��J���j�w��<�oiz5��|�.�"��6uOjr���}�k[d[����L���T�]��+��rҜ#b��j��D����_��e��|C�K;۴�D�n\�Q|����N."�ŧ��m����u	�j�����jr���Z��s�P������K���δ������`=����;�B���j��U�ms>Σ�G���8�~�S9�|@2ؖz ��:H��9!eb��.�V��k�#^C%�<�U mGY�\̛��H���ўɝ&GdH��.��(��u��,V���D1���".�zڝ��I*ܛ�5P�)�������H^�������I�-�C��/�>�
 }�Ќ7�����B`M9�%��~�%��~�I�O=���Y�����[1�B\�'����%\V+�j�?�W��5E��@5�!�wF:|<��0tk��$�`�âG�p�D*Nn�{�-��$�`��Ο�� �b}�f������4(�fYB�4E��8DOm���t&gĮ�E��]��mV�r䩬������P3����D��Z���_�NA(�ӗ���ri�d$��K�UP���!}�SXW*,��9^����0Kg��yp��vUǫ��m����<G�H���C���|���m:� w����=b茾g�ph(�u[��!+PcQ*s*�$��:��W��׼��6��:[��� ��d���
:߇pL��4�OQ�۽�ГZLT5]Q�}�8�N����U��S�O��Ik������(�� +�V��9�'�Gh�q���"����cj��AM\j'�*�Z�������=��1�`�!�µݦ�h�mVϤ�I����ex�<���f�������sB���� ne����	cr}�=�z�"�Z�}�ed���4�3��nI?���_��V��J��5ma�� 9A�6)��x�t�؁��>������\��I���인��Jq%�\48Y��.�jZ	%P���CME��Ӽ��;��{A�	$�?�@�Ҋڐ��j
H@��ޛ �7���a�N&eb�@��2n.y�l;|�]@ԣ/�-2����Y�֓6̢�1����]}0j���3"���BI&5|_=���H�� �6��_� ���*�ߟ�B��ѫ��[����V��5���#o��pS����v��m^1up�o2�Q�N�=�Z
1��S������`X|i[ٵ\�<��9G�@��)3HZ��?�:���� -���N�a�ܪ��x�LM��y��� &|��S���'�˼'Ũ`���	y�;�=���>���ᄐ��@醛����ߘ����*�X2�m�'6��b�ύ��;!��^ʑp�w[G lC�#�{�7=�:�!p���rۍ�\�����W���j�st�q��tAד���Ţ�A�ϊ[�#�n��*��_���@���D�#e�@��R˳)�����{(��*��i<�a�'�m��.S8+����Z�4�R�C��Oq):w��}�2���h���[���>�܁��fK�m��E��;h���|T��ph7`/7�rk����V����){�R��?��ɘ�G�HXM�-ˎ��<~MK1��z�+����g�L.Ĥ�	�u�{�	3�w��X�����=�M+��+$d�k �g*�t˳�Mz(�n�6j�L�Y&$Y�:�ݠ���G�_[�Y: �!�욁�>C��	��F_� ���.mY��nJ�mJO�>�eK#)��`���Mj{�����JzL!Z���!��c��5Uc�U�
M~��]�����Z��M��p���is�i�]ـNNF��'
ѝ��HU+�Y��s�9mXk�=��m�K�:��Ua�"A�`u���*m�|�S`)��p�0�t�����m8h<l��VB������P�ϧ����Y.�/b����7t4��<���!��7�yc�QD�V��ɢ(�v��Dtd�厊|�[0��pq:��Ô9�k��rv��>۞s��_(ʢ�=ZR�Dֱ_G+��ڰ"G~�����H��A�O��@��K/��V~Qv��fo��g�������|��+���ۓS[�<9NA\`9\�@�׏2`��v���r}�)�����:p�z;R�-��}2e���$QF�l�r3�TK�/��tv��[
�k��{Q�߹�Em���.��L�=3����ٝ ���sK�>V���_7�ց���21��٪�:�N��$�(Z�
D�2�N}V���g����][��ħ~c�K����}!�3��J7A8G��\c�6.�����uҨ=�u���|��h��*x$g :#�a��*f�-]���%�/�? nG2s&���k��rX{{�%�^/��:�W�"��_�w��R�Ӂ-�+�����:�c�UU�I�4�$�@�2#�wk]:�B� �m�:Sѷ��^X��n�8z>�U�Z�2>��0�M�0j��������_zo@��l�6�{���F`G���H	9n�	���.O)W0��d�{�D�N�}PM}�)6�,�����r�:O��X;��~f~��V��:�][��Ӹ7 ����Z�k�wn�D�>}Un���Ð4����-����O���Uv���4 6G8cY�(�o���v��&��
W��v�.x%CCG(B�iT̡��SF`YQ��]4!IwH�x�O���'³��*�bK�]�["�JS1F�3!���w$���>QC�7��p��3����O<M(��s�K�O��·����K�nX�z�m�Ɩ
��A��ȭ"���&S�fz�xz�ؐ��E����g�$��:w�U:.�4�0�UH÷��@���N�8}3c�N���F�͍�����5�zP[�	}N\pe�Dj$[�Y�z"�"x�2�{���1a5>�~� 
���9�ib@��mc�G���)�v���at�,_q��:Ջ��4L>ק?�!b���oҥ�Y0��=,g*��\��/���4y_���O6Q�KI���88{1�7��~�����Lێ�Iʩ���׆=D+���RE6߅F�f/;��+!���ʂ � �k"�r1x 7L����=$ԁ��$��Z�F��-�s����[b#�i���]86 ���l�ؔ�T{_:�e�vﶪX�~j�i���(�u�X����/,�7 Gk�G����� ���eʨ!v��~�q�L��.nU����~p�G"T���2T(�$#��B;?9�nh��j��u����۬��n�U'��k����9S��n?VJpRA���m��Fs�>���N۾����|9�d ��Q�-^h��"5�j�ʍ�^`�}i(�BQ]��͌�r�B��#�m�,h������}����� :���[����DsAϪĎ�~e���K2Πڕi޴��^���NХ|痳�I"�3�;�Ёnf�T��ih"�U�����=x+��F��w�~���W��&�59��1Ȫ]nQʎ�ĮUh�<:�׵��dls��W��ح?��4�J	�-���@���=]�S���L o��L�T ��������g�����1�*Zk�y۪�����Lɿt{lS�Uɝ,Ȧ�ئ�� ϭ+B��I��ˡ��^\6�|{�a�7Y���0,
��|�f�&�s��Y�-	~Q�B��=22�%5�K��Q�n��y�'�/�H�0ĉDy̹ck��Nw��jb���'�kn���H�+z�t��[�$���1�y�5!��#�C"WՐ�
S{��"*����y�'��b��͛y�����|��m�10w�#����b��j�eO �����}\e2����fE;�fL��7�q#~��6��	
�A�k�3pa�VA�>��3Aڑ"�JS7L���S{ J�%x��M����$���ҁnk�w_�˵#WVq�$�"sqa���۶Ő���n$����5Y��M^��r4��t
I�˓�GQc|Y����h,����,�E�3�sn�'������x���J�I��z�[�0���U���$�̢����N~��<^aU�'���<O�fef�Ϥ����m�����QY�N�Zj
����'�
f/��
�g�H���+�+ �`	�J�L5�<����`8��M����"�	�P���3���Ut|����?��-�'�z{�����&�o�'9��7˵]O ���<�[��rK[}����^$��J��`2��Ԝ8wҐ��SWq���-\C�N��u�U�j�4���~W"[���c 0�;i��SeK^�Z�o��I.I�"?�̎����>du��HB#���9<��-wN�ׅ{i.O���M)��~�ʩ����kC�7
���ީ�����E�����P���O"a�1�v����s�[s }���OO5���qU��l�5�m7`8���G	�����6�V�9|��rؓϯ���q�Gu���'����x��ڴ�Ho5�cP���*�녤�����!��<R� �>�-�Var�L�����B<��7Й�����C� ���WI�D��=�nW1�
҆i��f��1qG��� P��cQ����2�"�@Չ7Ͳ�L_�N�6�i.@��>��}e�ѽ�4��7>�F ɯ�\-���(�TM��G�9L�y[�":3��;�)�#�Wx��Ϋ�RU(g)���*]��Ϳ�������Nؾ�	P&�R7?���k�OR ��˿P�cMe���3v������K��(�r��8p�ډe�0D���s�V�%�,)G�I�NWz7%o�/b��?��gb�Z?�:�Z���!+mM�V���݉�U��gCi�g�ԊX��j����~�T�װ�!&�w߫�%
��?���������hh�歫KO�	]u��[s�����Ŭ��!9����X�y�O?�8���TF�8e T?2H�#u���2g�i5�mz ���V�������QM}[��J��4��.z�`�Uf���h�M!��˽�����X�iR=�9����A��T�QB���`'48�G=;��tl��ATpq ����n\#CjQo�8��ƧK���<�/-J؊�b*�~#I+K���w�����G�Y��@�9}l�5� f����/Ea�l�.Q<b����DJ��y+�Z�p�#�Y�=�l&t�<�����f�ɷb	���F!�Zx!{9s�=����S�ʧf�r��!�A�4��]I,���fB�+J���\�Ten�}�����KT�<d���*zRYCe�gVߵ(���|I{"��&�ϓ�A�/�f�O��A=���1��m���oe�.�ۉ�l%�cu���`�����
� �yb�kV��zf?�b�2�TSP��;/#ݠ۳����^�3���HZZ˙�464`Q>r-Y�Ϭ�W���I�k�ҵ�T�+��&,���S;'Ea��΁:ͫ(s/�j���2���j��㖥1XN�L�E"T�"�<�+��+��C��!^%;���Ƃ��me�{�J���`m>�[��]Ɏ�v��37{��u&�l*��x�l���ӺU�����e>ۯ��&t�S��;<D�c�Ih��znK��׷E5�a?��2���]H���'��8��<nM�MQ��s�Oa����x{ ��;��N�e�$^������U�`Z��u��BS�՘.ݗ�TI�OPShN��0��C�Q.��f# �]2��HhbkĈ�e�}X��5��F�̬�g��"3�&;Cď梅?�6N�����ƀ�C�=�_�~e��'$�K9��-��c�Kr�4��ە�;�$�+`�3� ܧ�Mz
�,6K���{==Nm)M��Y�`r���&��ybV��qxj���v,���A��,��f�4Kg�Wym�<h|��7�b�_׳����`쬫���L�i�������B�j`�7YD"���TDPˍ��<G}��UY
׍!��醳i�� v#���Q�h�L����-ONZo���GU$UL@t�0c���pT�NZ��t�����h�b�o3e�UqȦ�I�D��Ƴ���w͕�vv.ݝ��C(�03F���1�	��)c�@��%�Kԩ�>��ypÜbِ�).|���� �ף��K�a�<w�>��K�0��6r<�x5ϧ��u�t�ɚ8���`��G��;s��Q>V\�K���(3�0y1a*�W����mD�*�{�;��J�n�Tzb�O:70K��Afp ;�2�UWHˬ�E3"]�,?���ZR�M��T�{E��Xp<�>��h̏D���=B�BЊU �
!�g�e7}�L���ܛ�)J���\�G���B�
���Ⱥ��(<��g�.n����9�a�΅�0�[�����=��OrB�ZD%����\F*�T	P,��C�]�R"������_�cL8ڮ��y*Ie�Z��S��h�TW�%Э ��t#S���ʼ� q���"��c5����ӊ�
+;E/e!��q�f�Se^��,t�u�(�PO�73�vec��3�N��aS����a*R���a%W�X�a��wY�re�$W�e�c���<i��+�	*�T+B��~�c��B�8_�E��/���qs�ߙ۰!�Ca۪r4Vy��\y��l�ą�u���f�}����p-�v�N�[���?׷N�մ��^�u���>�E�
ʌcl}�C��`�c����t7����P<փMv�����كbEΩ�*�-�5D?v�.�р��0&0z�ŔS�V%*3^�q� h�N�!m��	��_��y���� ����:��b�A��jBɹ�P.���g�'�
S7��ڠ�¯F9�C^Za�~��/ں;�Beof�^�S��d��SyU�+��>�����wZS�^ Z�_C�y������ٳ �}W�+���I�I�Dܦt�m@>�;&Wv����w�Y��0�ѐ�7Cid�ۉuP-'��'t�l�����Jc׏W��r�&.X��"�=�\@��5O�����V��C��ꬳ�C<�b� �u~ni�N=w�_4��a��W�U<����^<�����߲��4	�MB]Om8y�ޯ��5�ي|`b�k�&�Z��� �U�o��մD��J!�;Ȭ[�d����P}�䘦4��K�i�p��ʧ�S���#.��es�t|N���I�2b�����*&�6�)W�?�,����Ph�c�Cu/e+�f\$'=Y��=�P����ܡ�ͦh͂��Ɓ��R��'���V�"��«d��;��]G*p��J�Ĵna�
~[�l�4�|�z#�"!�Y����N�W�R��f��S��cV�J
�8
@W���S��� � חT��4_)�D-��L�j>�x��������[�Η���bN1LQ�/�A�v|���	9���ـ�}�i���[�.<Ȼj\(x��E�$�nӝ}~����ASK2��n�쑕#�5J�M1�=Cb������	*�C�7��P߈��U�baz�CE�EA!/.����
�%X&9��Y���P�X*�"��T\k�
�D:an�N�˝�B� W9*4��=�H[ i�����w)���8ю 5��c�4�[��d��;(2��	É}������JHtc���ϕ����3 �x�Eㅿ��>[[D����:?NzxA� Z�?�������у��ާ�u�� .��8-� ԍs?*�FŚ� �s R~���P�H���5z1s�!��y��f"s<��}?��[I'�s�������x�s���Rc��9=c9��@���Sk��)�ܟN�u�~��V��
�C;��ܦ����"Pt���\C�h/юavHB5Դ����s��SC;y�d��yxm(%��Z_Z�~ܿ���.�X�L�hr73i�G;9zވr8�b�� ��w�,�,���FA��f@�jS�ȼ��Pm	z9�!�=}if���&�BP�'m���5C�S�����ȝʜ�YJ��)�����׽f�剎秋*� �x&L�����a
�g1h[��d���rŐ���@��9@�%�����`8 ���9è����N � ?熞���nZ`V��Y��HN
�����B;��j�t�i��\��&Z�}|�;���|1�3�WР����AZ�A!D��}B[���x���G6������A>(!R�clF�`�gz�A4u����0�<:�?/1�EwC��ΐ���q�V$a��`� �`ʮ>�<ޚ���cV�hv�Zh��Y���j��X�����ݰb��BsN��G\;��/88=^u�:��^+-��ܬ��QUTYKyk�9b�P��p�U��scD��x ���e�1ʛ8#�1fZ���2���R��X�]�l���q~�q3�CTL���O��B�8n"h��e؋�+�un��GW��ؤm�' ��u��Vg�<�cо��*!uc�W�f�4'���a#K�է�FV�M:)ߦ2�3j��Z{�����|%�Q��+1���7�	�B�y�gRr�a<�iڵ�F�j9�o�Y�����h=k��\}��p9�B&~���>���O%g��M��:,)���",3X=�S�N*q�C!��8Έ��j�]��S��RCQ���!-n��aSxI�ݎ��4,!)��ұX�z��OH��%vŜp�/���=ڤZ;o����3��ۉV=E�l�hVg�y"�V3|w,:������G�s)�7T螶+-x'�U�����E��s�����_D
�N��F�C��c�����w:7峅.���/Gc=��F�#�O��� ���N�M>Q���K�ӬTΝ�a����<@`����x�@p�n���φ]���V���zwt��6��Ի�.b�o�&�0�6�s2}Z�6#���{������j�{�hqo{q���l8�^O_��E�g�l%K�'�D�޳�x���ІIاk�u�ԗeb?ITu5[Ҫ�@{��fNJTZ��O(�:>��y'<�y���e�S���H̝�d�݄6I� X�sJ�dc߄��ቛ5v`��l�V�^zV�6sB���1^�37f�/r��V�3�?T���W��"���TLX���JC`�jp꿝c�y}������6�6��ב7�m3���K�V�EO�8�xl�Os���l��%�e%X��/t��`����Wi��U� ��o��ҝ����aYr޺�UXn;q�:|,�4?���}��m�Qw�k����ʝٲ�ݗ. TB�2Eh"���8����Ņ���)��D�s��P����x��h��x)�ULsR��^L�o�YDY�x��ߠ�:͹����C��,�&ⶏ�Dg���%���C���\�l�o<JĭUi�%�7���~H�8W�%��Tx��l-^�gE����*4����g�Iw�R�}�w԰y��8�LaCM�v�ǫ/���ۿ#�HwK i�:��Y�wCr��D-F}sU�kj�ZU�?��e��
R~�}M�щ�x\JH�J'2��\p�~8�@��N�j�𯽭Y3B�K�P���1�d��uMoT{<�ɺ	�	��[O,q6����T����'��8��"��.�z���l�޴�Q��Պ�I�꾥�uo�Ł�B���2��m餶���:�(�������9�S��*�qO*IܬAhEbl���)Ik�C	�mjj��ȷxE���j���+�D��@��y��M�}u�e����^�֫h��yːld�Rȳ��ӵsr1'��l�Y�^l���mN
lU,:%��IAʧ�e-J��r�&��Q��g��A'�v))U�0l^�^����ȁP��E7("�!���夡���J��'3mA�`#r�ّu�HN�#&��ܮ��7���l�	Qi�x�p=#��"=�}���������Yq<@l�W��ǥ���ܹ���ǳ���~Wߒ;��},�[fQE����˝y=#�-}{��hlC�N6��jMPm��:-�);��6�A�x�p��^�����u�%��'֬��������)dж�FSrΟHH�����*P	t�O��pʽ��\�����ŽS���xv�<zܓ9�����+֊�}c��	���m[�Ѕ)�&���{z���������D��P�>g�99ɇ�6�,G����/��#�QV˕���zqp�Ydo�d�%��� �d�W�or9l�)��F9�����KX�'���b,�=��#G�	��'c��fة�d$��y�*03�e%��Q�08�t\�m{����\$�r废��͗O)u�T��K#�Ȣj���ڐ��-�-M��1}��#	�ha�|�֌8E8���2���1�)ԋ��ޑ$�rd�=����ѳô�xL˷�k���\�F����CEBw�~�ۢ�V�q��R[G,Bs���]-CF��H�M�e+>����ś�R���Q�����Kc��Ў�,LB8:%���j(��:6�����h�׺5!2V�Z:%a��QGd���Ε��3������ 5w���yc���+e���x_�y���)n)��,���|@�d�#"�b�tU����}E����"��]��?)m2vs.?���	�	�?������]����+��Spj磕'��Qw��|���W����?P<-��NUy_�$��\Җ�q�+����t��E�@[[8a\ ]���T����w�v�r���`��l�n�?���i���'��8F4�b]A�MG/��u���SZ�uѤ��m���E8��Ʉv���k���៨/����iH"�u�Y�[n��s�����$N�_B1���vX��y��Aq�Q��B�"M�B���E�.v\�����'e�py�`l�M��1q�*)K�
��k�OG��pG�20�g���N}�杠�&�F�3�m����!�(X��U�o������z佯�kk�7�sL>�(
������P��	��� ��&���Jm}1��鰰D�V�s�j���aת���cS7a����_Xo�I.��*e�:���=0�e Zm�����i�]�0������F�v�*U�X����m��H��r��ӷ�ÌD������:��<	~
U%�,M���:�箝��t�)Lc߂���r��mto�zϾ4��ΙL�2P�����BH������8VI�?l]���B�3�9/F���AiGN
���)D�*HJ�j��w�e�c�_o2�u3�,U�e�M����?�H��DB9�T�����Ȳ"db��݅�Oꘝq��.�5&�S��/ռ�7Z�1�A�������%�&y�l��n���x��=�|��&J��4.ss�ᚁ0F_M�u��d�~�:ƾ�?���w�W�>+�.����!*j�I���U:����A��ZAخ6DI#��=��)�����
}�3E$���H¬<v��ЁW�,%����@ƭ(�g	�
�rz23�>i��C�(}�����_��ؽ�y��*TQR�Bt:4##�N��~50�>�U����o&��˻���Y���P۶깬zu=F F���O\��D.<A47�#@C9雉�,�Y�=Tl4��G���1��f��_��<�:t��e}����eK��|y����&�����D���� �!Ʈ!	�����NJ�t�M��-�/A�9@��,tdF8�OO�h��'��u����Aw�SA�����}{�x���_��S �M2Z�r"'�¶0��d6wP�܎�?>�	$���h~��b��D�����s�ntU5�TP����/�j��-1�`�9Isjc��w�C�������P:h>`�T�_0����Mc�.
�i�Cƾ��hR�?P��a��Μ��)�n�����v3^�(�]BCyj�{��Սl��;�
���Ske�YA�X�e��gD:j�X�	���i8�l~�V�u�s�&�` ��7�"똕�*���l��<�{K��3�笂�'�
K�{ٚ��Έ���z2W[��=���뫯�A�݆}�}��t<��ϊԘ�*l���3 x~����c�0g��r.�ז6�H��g��ZZ�N�TUT?gQ��&���V�������b����;c���[U�����(�sQV�q�b�
̣�̔W��:q��t�\8��|�82����\�X|�<Q'p/B;���1+:\ ��àrsF֤w���Zy�R^�w���Bm���o�q[s��xs�(��_Z�}H^�L:H*���:�#Ҭ�@�)ڼ�H�y�w���}�+9��P�I�菧�,]�;��������.~@7_�9-�H��J�t߼��}��& �}�xrP:m<D�u��{	c%�p��ܠ���-d��8�d�;Y�'��v�
+o����6��h"h���o���T��-�z�M�=��e�֤c�7x3��z����.��� 2�@� sV�����
�TM˂�N��i}��}a���P�r�L�+���(�X�i���ЖJ��D�u��@�E�B�?)�c`,��DA���;��|��嬂�:+	�(T���=���M?����Q�.W�F�9j�b2�'�ع�M|��c,�����m�]�W�"G@_�ǲ�	9�Ǵ����\Wi3^%����X���b�)]S�3��B*��T�E�!�̴�<;��a@y����Q�"?��JLr�Y`=�3�;.2�ߔ�1���8��_�u�����Ɇh*XC_�4ޢ%p�Y~��/-�L�/��Vxa��|hb��
)̀�0�81D&g�
a��G����%784�d解�![a�0i��� �H^y	����97��Cg2%QRi��ŕ]����2s|L���[=���_/�tL�����P�\� ��E���!L����i�~s��?3�N|-I�\�/(Qt�e�=�����:	���Q_�!�J��B�=G��:qL����>Q��X5�;q)s��7���W�Cߔښi�R���bcX�����+9���WUX��s����n6�0{نF�Sߠ�����`�`��h��5�A�]q1O����'|��)vf�r�T����ӥ����r��wI��Ѵ�E�;�Æy�`�;�Xҡ哇���N�A<,eSV���S>#S^V�L�����5�tUؚDϣ������a�8&��J_H�Y�*:�AF�`2����G՚�R7,;�E�0�����b�<;��S��Iǰ���F�~gPY*픚���C	[������x�vu��ӥ�|���2��q���;�x����h5�Cڢ�{�0����c�ֲ��c^�'^��i@��f`�B��Q�#�Slr䇲�in�B%|U��1�jEO��7���N�:8�_J᥵ڙ��>�j����P�Oz�)�N���桊[�I���,�Q%Y�07S�u���Q`:ro����
]�鹷Mčܹ�n��8��+��xz ,VSk0̀��%~�yr�[
����T�=��rxV�8�wh���xݷ�.����p�����\R�"��+M8��Ww#G�&mn��d���^��֑)�W��-%�Z�/X}�8'h7t���C��[+ABR��3���n)UN��̐� iO����1�2�/#�6~�I�	c����xC��\�L�YLR��[,|�qV�SX�ѵ`�4�<�@���>�D�<.1�ı[T�(Hi�y�x p�)W=g����E3D?|+����ɉ�ܛK��Qq���[�y��淡#�E�Eq�_ַ���M�Z�AAF�>zH����-�;,�^b���_�F�9�ie�X� ���x+��Y��ji���<f9����3i����y�Ilీ U���S������h�6�M�W�����@
J�e|IǃK_�^g�-��~�ܓ�!�/f����:U�`�9T����I�%��;�'���>��J�?��Oh��ο4���Sf]Ã�G��"�Ѳ�M��G��g�W�Ʈ���=��(%O8�kġ�']���6i�sĬ�6�g �厀���1_�������6Ikc�|����͒
�n�٪�b��/g���v�9O�n��a���w����vȶpV�Bb��������Jr�2T@B�Y�`���N�|�Ae�h�� c'��,�e��R剪�3y���)��,�[���	���#U:Ig�j�<u��Q�ڰ? w����72�H�h�(�ǅ�4~6�N���A�#��.!Q�_t�Q��8��� ��s�4{�&�r����|�C��.s��s��S�v��7�@�F�|acZ����v���C��&C�'��6F���P4��ƙrQ
 ݣ'qo-QL(h�M(C�iZ�dYn��R�V�M��ː�G�Q�2O 1��"nW�B6f��T���
h�Y��m�
�(Xe=��p�/��7��.Nن��5�\IkT3����}�`��]_�����e"�Sl'ԣ�nP��ﲉ[��w��<U�(��E�=>V4!hx��&[����.�+R���D|7�} Uj�f��H ������dF.>ed��'@4,#���)Q��1�+��쫙�؛��Z�j�׍Ufn��Mq3���2�d�;��bF�y�P]-���^��/�G肮�B�K6�y֘/�\�^����w*6u:˜q�^7>{���/a��&F���3V�t"���3�3A;$>��[�0�=r��?Fm�?�Jʂ,G�Onz�g3�������Vw����f����J����p}dr�� �O��.H�'��z��� !�._�@��E&�.�ZP�^H��� 5ӂ/�Y88 %�:��s'���d��sks$���WA�1�Nz�]L��kv#\��Q�ۊF�����0S�180Ib���&)�L�Y˽�yC�9���"@�fA;)�x���t�"8�\��T��n�K�RdW��4�(�6gC�_袪�S�ki���6�A�X7B8���C�ȋ����I�ҧ�FX
o�ҤoZ7��gV�����kz>��T��ܵ[Œ`4�A�{��8]ML�<��o~�����ퟡb�2�৲�us�E2�"^��.��G�<��s����$�:dޟh���(�����@�^�yc��h��^;�"}9�ΧH\Ng����� \_��i
����{�8�Ûn���`f�韙��<�H�Z:^&��7wkA��&�(\W*t>rA% D���:_����a�1�i:�A�x��z��b�֦���UsE0���I�N,����J��~����$��N��?E|pǿ��2��������;����P�)��M�HHՍ/��Y��e��O7�����Qtj%e�hY���Ii:�H�i�����[��.m�?N|6 ��D_��ij%pX Qq�M�orWi(8nk8�"���] �J�_�6�	o# �\!��:��\2Z�y���� 1�7`E������H�+��|��:�+Fi洃Bk���t�U~����K�#�\�u�a�^&���ͭ����(WI��f��s�f��fg["��~�e�)?Kh��	3���v[�`�p���JT��	���7�IC��
�dcL�70��f�W�o)���$'� p{*��������j���,�v�wDm�[8j%X3h�t14��� e�a��Cݣ*�M�[_���Z�Ծ �����qV�� ��@<*��m��/?ޟCJ H(ȔW}^�@���SA�]ˁ_��]�>�w�Iqa�T�@7�إ8�^�����S��b��Tn�]�E
�H�&|�7�9w!���<���p,�-�U��a��4q�[�Jߔ����FJ�J���6������9���b���o���h��f�,��gl7��|�UT�#l�v_���`�f�a�V�:I�{�d.ϒe����(5�.+s�}�|�	�_���-JK��2�Qﮑ>\�:\L�)� �c��l�8����e����+{��L�J�����B�w\|�DsZy�՗����M�+m~Z���|�h�H�+� IY���3$�C+��h���!j1������Z#�O��&0��h�n~C�0�(�Zf�>=���5��/k�uo9�T�m���J�M����3=��g,٧�6�<��2������TȌ4����]ֆ&��m�q?���><���K��bur&f���&u�L���I�.M��Q� ��F��ϓ|�s�v<�"�l���D9�J@�H/��@�)/��N^s�b���A�;��%�>�Wb����r6�U��r9���R#F��#�W���*����?��x�#�����-U3�06����!q���ʙ���1~�yh,TA��.a?Z[߼Z�Gx6@�vG_��7\�)(L�7{�(P�\YU>s�XE����d:+ F�(�P�Z�������$�#G79��<�W��;�{$�����t.g�� ��9'�D=��w�	�2O$�_CQz����xrs?3���y�Ly)$gF���
^*1�{�@a���^%��G&d�6�X.;��}�*g��#Ɠ��p_���p�G�<!(/ ���y�JVQ��'e�!�K��z�y�W����I���s1|X6��@�^@#θ����&�9���	Fi��T$}+K�H���a�>/rx�ߨ�ɡ�}���/�i�Y���zGTy��"h>`�&�o���vWpb��q��(����#"��=��ܳXa~~zH\�a:G��s��ڝbޱ��)
�k��$s���
���T�Bh�N���<G��}���l"�ϙ�&{! Db���![R���˦ X��<��f�������ܤ +��7�-	r���\�-%ԣF�d�:D2�(�����33�i�@��z֍}[{:����G[`D��(@��;�ϓ���Z�W�v��T����T�������7Au���D���n��h1Z�*����7���=���ɳ��_��+9��M�w$�"�u�:GE�.d�X��!�k<!L���:?�|�'��z=4i�E'��J{�3��k�̏��7���rh���o*p�9F���)��Ńr�	C�^غ���0|�\��,,��$Ї+�z�l��G�0��Lh��x�w�/�<.*�����F1�Чm߁��Z,���A�Zb��Ǐ��DruA ��b�5��؉�(��ݚ��s�*M�0�4$���&j�F���C�	OA��[A��!|*�B�!����)xAwzD��;<b�����:㱝�����7q�M�
Z֥8Ot���-��
�$�8�L��C���*W��t<�����o��"�s�'�9E�E��IR��##���AQ��j8v�y�"�S�iV�狛�#��kH����8��!2o,|	���9GKdɝM��r������~�MM������K~Z�R`%`�$n�W<�2���$��z%������X���TcL9����-C�k_ �$Lr5@�i��b��3���:8|3�X�>������H2b�>�� U ���q�%�[!�\B h.
_&;r�q��G,0�U��:8i��,�q@�b@�o���,��(25n|`��ܬ9�G���i�T��R��q�ЬX���?�z5+#�����D��j%�_Б�W���N�T��?BZ�/�>ڂq��)EuP@�X�D��@Pg�%��ly8Q�`a�� z�f������bbn�����P�G!C	��I<���W[�V"JO�5�ݢ���*�[5��\O%��-'�-T���O\S�t�I�0|�;l�\��u��~�����B�u��|(e<DJ��;���G��N��r}�5<&�a1��P���'̄)·P���E���xZc Q��n���ZO�r[g�Ej���fe���ƶ/y�n�X�V�P�w�ٯ�fӳ���n�IP�]�x3���ӑ��L!<2Ј{�U�I��N�5�*���%�~��|J8�S��Phk~Yƕ��zg�cΏ@ ��YN
��A9�E�=H�3��TGWu�y�:J�*�!���,��dѹ�����]�GZ'lfJ��w�����Z��b�$I �����qut)�]{|��)��lC�!�.����k��q~��'T��j��h���}W�ϊ�H�S;�{���E�˽�~��r�r�wpX�9Z�΍��!+s�����W҈����+1�ϛ�)OJ�7&d��'�E�X�- wx�������e{8�BX�������Ssʢ���֗+��p�o*�s���N�{��e7O�h^���sdnGI��k+vK���X�Bs�e���|��3���>DI%�^�*�ɮa��7�*��$.�TL���g�w���$�.I��*6yu�ϼ�B���%Y��Ϗ\ �/��n�
,{M���X�O�.GXc�v�nK}�U����zH-�2:�&/|�.A u�(�{I�p�����[M-yYx�tD�0o-����Gmk�.�{��Ojޤ�Qr�w쾊H�&T�}4����Z>�|��(�I�C�u«A�U�Y\͉��H���CE��s�5Q`�v����T �i�����j\u[���P����~�h˨>��*)��p���mXK��Dz����\M�h�H���<˨@��9�fH�r�fsn�'�P�q'�z��y(�8��#��*lu�s����+{⒙��c�Pyɋ���SDک����}kQEJi���������Kx9�A3��ެ��/W(]m���L�v�҈IU���mf��Y�ޔ���ͩ�S��tb��e/�Px��j%nE��6Eos�C�]���c�ޙ)��,� P64�xN4NIuA|(p:�"T#X���I�׿�d�
�?��8���1֫��R���
�J5�Ev��H��U�QV�Q{�lel��őI�ըi���y����P�3Y��5^�{D4a.�C�G��oM7j�)M��ࡕ����Z�Ʉ���?�1�˿�@!�%.�+_,�����q���И�
�o(+W���S�)-煢#^��W�lyt�"������I2(�0�r6�#�V��ĂN"ӿ����}�	� ���xE3l=<e1�6�M$tsilimȔq�)~���P�#�>��+B$�|��+�^A
G<�ja����K�PD%�e��;ː�|����ޠJ�\zR�"�i�M �S��>�<ʺF6EiT��(��#�}��h1����]c�̗ 8=F:Nk�5&��p���hT�!`�f=By��!(��̦j���X� ���	����?���w�c�7�uQ����&�r�!�_&6h��Q��ЗK,���k���������}F}���c^�SG�������kd�
뀊/J ���Rf���s�X�����^������mW>��/� h��P�:��=,��o;X؀�;�ُ�ϴ@z����6��f>���x([�����#���$B+��|�g����-��xo��u�!���?,{�O��hj�|����Έw��"�ˈ�)� ��"m�]�����������&#ې�Y,`g]��1���[;2��9�@�/��g���Z�ʎR�Y`6A�t��z��y9�0�/.B�\�⋠��hñ�������h�&��!�Q�vFdg ٞ=�<��,�#���4\��	�}.#1�r��GpI�=���Yfݧp������h��v��vӺK`.1|�K���)�ܰ��Ə{��p��p0Q�K+51^/�(�^���Wݨ/�\q��M#��	�\�að���iD��c�Ԩĭ��$\���ai�Ǵ�*�ާm_渟7�5L��jٰ��qt�h꺄�Mya$��j�i���[,��� �����9W_�����?��JxQZ2��s-e�T��h(��?y����a��V�ł�
���$`Pm*����i?���^|��2�=�$�@�RU��R���h7a[�K�,�z��(�c{,��������zs~� P��X� ��k�7���|]6�幠)kf4R�pZ\�j@�*�̈>����}k�pB�
��Q�2cO�'��X
�~pQ��4�����B�>c-�j�Z�tߊ͗6�{K �-M��`)��yKcr�mJk��!��(���U��c�_�?�CQ��x	��
M�<����5�q'.K�-��٤�^���)w� �!"xM��)���gq�kJeH�3rh�iq�������D�#������>�)�%���2��hY��}�E��/8$� �M��Kq��|��Oq1��7����%���'�19MAiR�I��Y��\��q�� O6 s��n���Nl�wC�^~����j(�w�M���L�LF"h2J�P+�3�{@J�[7VP[~A��3{�a)���f&4�ˤ���P���m#{�����F�w�����	�4�1�[@�4��?!�	c.d�K�@o�����ɒ�$���<����(=�Us�v�xc�7��]	��b�������&��� cc�>��֊y��u2�{�E7�tCGA�@2d�k������J_N�QO`��?s�3K�����+1W�����Ϗ�Dd��GcX޵}�˃�ȓ��H�I���y߷�� ��
��|��:�)w�);���Gmu'����
�b�uR�3�ߡ�8�aU�&���xB	�����6�g��bFF�ZP�k�3+�D��gø����2�4�����K �#�)���Q�����\r-z�d-��zo}��NR�C��z/��ŉ"ьz�/����$O�gu�ٚ{I$�q�4������xE��_��{�.��6h�����h�ŤC�:��5���OZj���Cfu��:[bD�7Wݡ�aȂ��qG�/)'����y�A��H��sşvծK��y�2/`T�Hl��#�m�����o���s�N���^$���9�b��ޔ�a��-��}!Ǌ(���w��%e�U�5'9��
v*��؅������3 q6��<�_*�;�`���`q����-��SP'4�wNn���BPc��Cle�0d1�R�]n��7*����'K�03D�
�<|]\O�M��dK`��%J�J��y�|�A"����	���Zq�&��ϟ��J��`���Gt���Hy[0&�I�)��830ާ�� NH̋�~�H�R &udh^�#mK�����Iy{�7}U&W|�R��)hɕM1��+O���� ���<����Y��մۅ���"�L?L?���/m#ļ���n����Q��2.mC�	��ԎLݤP�׹���тyD(��w	$�h��\�.0�NL�ZF���+CU�z7���=���U��-�℆�-y����n��T���A1N�M���P$�
�x�=Ή�Ό��(��~Y�'��1y��nB���1��=�L=I�(E�rk�4pHQ�j)����X�b���۵�\����$ 	�,��Ԑ�mG{r�7���š.����k���H�Z�����6ߐ��C���I�6����G�$\�phR�X��Wm��=�'�<��5]Cs0�!T�{��舕�8�tp��s��+04�>���KWk����֥�$�����_f���Ʃ�'˻#DD��0t�[����9W��Y��]t�;�8>�KW/A
�AQ�t+!r�2p��[��M5F���.Z� Ƅ�iQ�(zZ�i������븩���MT�W�e���u��#)�I��3��a3�R�<#�}K%���S����t�ÿC���I��j~��v�h�P�s�R���!q�B:���>��4x��Хjo}'�M����"[q�T��x&Q���1����y���O�=ɺ��@��tp�E�x!����``�s�P$���&��j��Z@+�L��~������{iKF���NTR<��8����Δ�ᏽ�21�}W�����'S��������"�V5�f4��i�*ΏSud��܇q�LL��2:�${��4Q��n�*�%��jL:V����=�b�2ٟ���r^Q找�tg_������?D%#"�ԟ��n�K��G;�J !�[�]���RLLX&mHG#��C�-�����*���qwGӐ_�ē��ܸ�s���/P��W�K�������Ъ�*ϮR�e�s<;r#ܜz(���9�sr�Tq�YVooM�Q�'b�SZ���_Q8g*�����#V�;�ny���e�mܼ�vgc���kC���^��۝�BM�h9ہ�CQ�(�E�p�XTIp�n�p�n^WMR��v�M��i��o]t'#��M���Rb���?>�y؁k�+-�(�Ɉk��#U�����:���K^��;�@�?�� &gL+V��RFu@��K�:F��t�I��vM��~�C0n	`uIf�9>��Ωb>�ܫH���eU�"����N�t�@��W�u��w$���'�:��Џ�3�@Y��डJ�5�&M��~�f~&۾���h��'	��&��使>?���]��=ƥ���4����D�Ok�		㉙���c�(3�2�7�vv�z0�^2��b�����+�t���M=?�m���F=�8�Q!�@��>"�0�Z���9����g���Ӗ�"�O�+�xx돘e�X&ܻ�::�����G��bq����������,+RUX�eyG�U2.�[ˉ�@���7���s$��a�"���|*U�8����{m�]~xO M�_T?�/@��]�N>E��`��i�zl�r�f��x��k<��[�H�L�%��|A���SK�{�ǒH��);���:-cu�ԅa�j(&�`
��|�a��e%R���/�B�~���D��yO"JDB�K�|R��˻寮9%�K޵�j��~���/H�vd�X]}�;��[h
c�N�L��	���C�3�26kY�~?��0�}\#x��s\���҈[5G�m�:/XP{j��C��z������Zq�8��v4��)/2$xF����w�k4�ڌ:�����g�b"%!�n���ٍ&U仧�qB���o��n��,�H~4џ=��C'�&q4��p��C����I\IT|��W���$�(�$
�.��፨[�<t����l��-C%Q0�uH.py��%�2$�� j_K��KF7ʽQM"2���6�����_g����S���1LxY��Y�j��m�$V�F|��%��b��v�m c?eVw��Q8�þg`N�3U���"wF����i�"��*	���Voa�EƕV{�������ΎLY��葉es�~}|��U���k�� ���Z�qZn�(�G�� �ʑ&e1���� ��	�es��{�.�@�`_2;za��I�k����N��S��=N{t�w�[���f�J�I`䏥��Z��A&U���п�-�����T,�r���q��Dv;��M�>[���gW&¶կ���Ud���%��4�y���|��!�����!^�6j"Be��{UC�+X��7�r��MJ�$�3Qdp<\��W*ޗ���Ў�����|��B�;{`�KJ�>�O�8�.#"��S��F�����G����r��x����l��I�޲�~�� �ǔ_��[G6!nBr��s��@�t�?Kur�D�����H
"�����9��@	 yuk��c��mB��$}IؤZ#	����q��Uy���W��� �Nh�v�i�
�ٗgT_�F�¿'ܱJM�	�=�G�<���2�8�i1��o����1Y A���t�}�u��|�,����J�;��7�a��H���9wO�Fˈ"�Dl� �\��7j���?]��^pNVz	#K�;���T	�fT*��<]�{�ڐ�$*��X�<�C_�����e=��r·�&b�	��Q���_�.q�T��6z�}�g��+c
2�0CS�N
���l�̽�v��������5&C�윜v��?�"�ӻ"ꑧ���u�)ʡ�Sc����w�I���?(�~����S�V�����*9�Ƒ¦�y}r<=�Ar�qev�/����Z�܌�ŷ~��"���;�;e��0]Y9����,U�&��Fu�h���s9��o���}r	k���D�_��G�)���Jx��}��#1�����`A?w�&�b,�F����F�e�h3A�踁���K�i�BdޗS4��S���f3kOw�J�΅��H�;뷴Gӻ��������}
1:.E��Z�zTDy�\��1�m�޿��g/� �M��x̤�jn4[����ǅC,�<+%�;�Rت[��㽽,)����t'#�+�)�'Ɩd����fP��1��Y@�\��3ϋ��#��Ҁ;����7���f�ɚy���bTSŀ��k)��x���h~1lE���k,<�Bkx���P�924jAv0w�RO�CM�8��-��i!��ѩ�l)T{�
|��dL�UG�a�'t+2��uA�eH���80�2T��y$ ���t�iz��2��ak�Bh�-`�߸����+� �K�Yހ�f���!b�ٍu�Cl�qd��a��/zv΄����U3&�x?6F��[�J��gE7�,V���-V�.}��"S���#�#���6"؞�H�2�H�1�?��5B*4H�'1�ۖ�9�z��DJ��Ѩ|{#���jY��(d�_#�1��t��C�Y��T��I��]ĂU�ϩ�Y�ڈ��%q��0���a���˶3P+ 4�O"t.i�5��}mm�O��(N׃�*]�B�O�e $�I ��J��E����s�[�pD�B٣�^C���06�!8J���t\$�z��|P��̱/]�&��.��^UJ�3�)�����ln�!��B�w�>�����i�)��pl�{���ۋ?�H���������}�M�̨�,��&O����\A�2K��t�|Q�����mj��E���U�F���V�7��:��4�j=w}Z�'�'7�0d��J	 F������q��){2Ok�ċuU.9�P6�-��?/�t���"[�&���;sbq{���]I�}�6S�s�
#8�pI<����lZ6����9@��j<�ӛc�Ջ�B��{�X~�I�ǘn9���"!G��3�t!��]���(ɿ�p�bQ���1UV����[� )�>�i%g��a��s)�<����m����;��sII]�R�I���>������޵��	�Ø!����-���\a��.�j-�t���i�Cnn�Ö��WY�%~��QX�P�ΰW�_���-���𱀣PE�ʱ�+v�u��Pİ�QLh����.���%N��%�f�H�Z���Y�Ώ!��-�����:Jgf��xx�(z4v�t���é��F�g�gJ�҃�l0��8- ��R��a�O�S���A�Jq�h鵣�ZML[2�L,�a4��W��3�dHx�5�X->�L};<	݊��d�=y��똪n��
£o+'�L�s}/Q�n�yC��%{�O�P��u�ƙmh�
��ʖ��/���b��cG<ln�C��%���Hd���a�Oo�޴�;�a����{;#>������j;����u��f�3�\�ֵ��?�f�ew�'2\Jb�־�}���[��V�f��?3�sh�*H5��k�f�^�P���� >N2YΕ�N:I�� \]�E�6#�V�O�7� ��p`���I>���5�bM���wmJ�R����D*	�˺���[�8�.���׎�QN\B>���1Wf������k|�%D^b�}e0���]�%�J1x��*.��4E�njں��My8��,����`@"[�&`�������H�U�k+d��p�t���~�Χ��(	��j�g�G�w�)%��?�#`����&77N�]��?��B>��σLp��"D��L��s^�UO�$�t|��i��В�'k&�����~�2�e��@鏶Q�����X�)-�\k�-��T�$E��[4��e 1�n;��"�
j����p*��xd�~��}�Nw�'���O0<�b%w��>�;�J��v���	<�C����,ݬ��|Cl\�{=.�
�"�}����`<��c4<C?@���7o��O�=�'J��˖�� �>��z������_�	�/�&:l�f�BN�K��|�N��9��|&2����R<'��^j��)�rD���S�^������ˉt���M�=;޾��-#��%'?5)�i�<o��������ֹ�y�sؖ��+k+�����������I�+��Ӽ�Լ߭�#��[۝��ʱ�	�"�&q�ɯr�J��Ϸ��`���Z�����tI���	AE�R�g��^��.l������4y��8+$�pϒ�pbwas�g�>�}OF`Wi�>��e�؊��΁�߆��C�^�Z\���AJ��m�C�ɼG�Q�,���刯>��J��>�Đ��ּ��~%o\Y�m�x����''���[�Q���ݕ�Wмe�u�W��2I23Uq�R�{��3e-����3M��O��ˠ�e3U�����v�(|h�g*-��I�����8N���nk1���Ȭn�f������!�������s�d��T�J�3S `�3�L��"�k�-�wht,��P�ڄ��l�dn7-ja1�4��]ཥ�&����:�����lM�}D�/0P���"ׂHG����愌���Eu��"��~�ND��o�{NC�,L;"v�s�L��5C^�b��h���w��gcO�&�Պ�9�lH?�fWN�n�s�\�Jʈ�#��J�\t�3��ic?����Xʗ��ܑ}�?G��^^���iB"`��)�
�
��l�Ec�FX��3gɝ.�=z�}�����ՠ��W��ҽ�-�����1(�`jwbZ�B��E ��V��$ۚ>fsۘ�R��
��W��G��J,f�V����K��blj������(�����"�l�p��Z2ky�W��Wj����r ��؟�0Ru����j��8����'�ᫀ��{Sٹ;�d��R�P�/�_3=w4�}�z����_]��:��n�y<q���W�5��<uӠ}��ڎ�]� Za�FV�GJ�đ��Rs��Q��WW#�Yrr�u�EQ�ր�n"���E�d�utzZ�}�`иGy��Y��K7g��|�Cyw<;�,�0���0!��@;2/8o}_�2��b���Pd�J�m̒��WO��Uk>؇��@.m��Ek�$:�F�D�ED&�RL�`��g"8i�;�7�e�ٓ�@�6yR�~��Ӆ����0Q#)�����It�'��{� �H�������GWp<�r7A�z���=����}C|%�;hBA4�*�J��r8�-V��O#����D�ݸ��ԁ,^�h�Q5���+MUZ�b�6)�X&>w����I�u�h��"�8�����&=e�}`�����y(��;�ؒ�P����Bߙ��VQ��wH+����y�Ņ�Oz E�z�h����N���/�Zt��U�*��*�rw��A%�f�����ЮN�,%�*�m(���X��Ϟ�=��N���'d��a��7�l5ۂ�I7����0�zuF҅�k9A����+��4	i��߶��V�ʪ��["=�^J�
����ܚZ2p��Je��oi_��f^�um2N�M�m3��g��,�Igk��6JL��=����x�Iz�nb��>�t��c�=[ɖS��K�^n٘S���
/�έ�(Q�H�dY@���\:�n�~���==�M�.te��@X&����~�*��Hb��� ڞ���p�����xs<��\�3>���(���} ��g�[!��K�s��F~]����_�ཻ5��Zݲ�AM�%�hC��ߵ���Vx����C9Le-|�ܙ��W�(����{�>L��74�5���������Vp��]���;�~ub
3��{|+	@ځp%69a�1��(�q6������a�x�T3E�z������EZ�U�A�S.tR�D��: u�܈�DK� ݫ�o���-�r <���t)�fuї�8kRQG�L�"���wPw�n��?e4�d�D�-&`�,�����'�X\|a@=�o�\��)��$S ��wC��$e��ҏ����W����8��<x<Z\8Om��"��&DI��r<�y��'?(��t�a,��Z�D���M�����+U!b�j�����# �]	��T��SVq��`��G_�jC�����1)�����
H�G��1q��J�<%u���@5�/7>���!V��s�,����P+�}�#�1�|�W��^/u�O�^������ON故wRdbWu��hPMNyםp�`.�Մ3�x�J͜��Jmud)(z�d7 t-%�l7 �.���Ks���	�L!�#{j}�.��e�/-�;���d@�V���V��O-Mu?j-F�m�7D-�3�آ��d�=*"�h��������,T篵:�ǭ�Hr�׮�@2}��\��A�Ԡn'iu���w�AW�;��$�zn����s��*΀��i�A�~�n
v�i�{/�Ĳ�

��Pd�������"���=lH��l��C[�|X���̸ �ݺ$��r*��p���I�s�p�:�L97�SE����>�tKn������J<�X�g�ة�\J<��I&�Pd«�i=Tw��MD捩�ᗉ]@ݿFڂ����������R�L��|s�Y�r{7�O$��2��Q�鱋P���&���u.�Z�l�����F¦I�F�q4�v�#�a�3_U����\�a������n5]�˩X�z�?0sK��fv�9�<�����Q79Tki9�撄X�e��7$�/!-S�b�YA��G-�\����Ö��@��yaMw�*���Ȭ*�]��j�l\�����pr������@���65Hz0��l|�a y_��Պ�'�ڐ�8�Kby>Fi�13�R��t���#/+ٵ%#�3��VC��9�2~�|4�D���#�
x�fX�R�)&�����GO]� As܏J���вc���(�K�I�d�B���:�0'�9
C}�E�K��,5��f]e�	/�uu���נ:��4���[-q���4@PI��9@�yߊZ�&����m�P�M~T�ت�*U�Gnξal!�ID�:�;CP/�S*�g�'2Y{*
'7��=�~"t���6�hK묘��؇X=��A�TK�D0���G����yX�#��ߏ�d,��!K~:�=�Dw�>�\��x��"Ӛ.�a���z��ouUɕ��i�k�i��?���)���}���O���N��]�c<Y/�7,#b���E�ࠖ;�	Tc�Q���PE;��*yKu���9� ������\���GtI�]i�i�7<}�*���b�`E��H���[l��S�}�L/d���ddʯ�
|�'����ťЋ�w�rd�	�a��AS�䉹s�a6����#�֦�Z�-VL]�ߢ� 
���*l�9do�J����z�s�>���2w1���=�-��U�����k�!э�_���y���	�|6E=�}y4Ӧ���B�ٖS?���|��?�O�i�$'�Ms����(>�w�s��?5�fɮߪ(z>���R�f�Qj��Q��Y�-i��u0�!�?d��X�wں����/:*���L��,���4� �m:��6����AB=�S8#LF��s)�Q��܌�J,+Ɋޘr�EA.v4"�j���n��mN�t��4#:y�m6�²���:K
i���Pc��~b
�W+�XEώ��?9)-aŬ�Äc
��_�)?��?L���ne����Z��J˰��%-�xT�:���űFy�	�W!(��f1M�������K�����C����t4|��/�l�̀){1<@N�����dw�[�;���=e��rݙ��I��
4�_�^�q�l~�b��[�E;̽��H#�f>�9���c7�̶Rc�d5�,	�.{��}^�䤮D�&Ǎ���tl����=�Gw�Ȓ���f5?{v�Z���'�!
��U�f��F���&�~���s�qS�W��;`bÍ�MKQZ�F��5eFR�"���0��r$������W�4uY���|�B������P�g�a��(��#,�L�0��7#���Z�������8K4fF�&=��8����b���?���0U=̶f��l�R���㕱PE�"� ���JXz�I��]Fc���7���0-P�Z]�{�h0�t�tq�A�JH�D����KL@=d�b|�H����0(�QCP�+=��|��Q�������#'K^�Ok�W�Ұll>�N��ż<�[�D���2l�����#���Tl��U��=)��~&͝�Mi�2H:�u)�AB���y���
�~>M!��m2^+�qL�Ʉ ����@����JW�n+( tdx$�n��eE�Cy��V�U�>OGg���Ϙ��x�Xz@��;�LT�m�|�O��7N�;L�$�؝h�_����&�'o��:�u�������!�6$�S,}��_uѲ?ͻ�V0f�g�Ů�y�=ط�q�#�p0�M��ZARM��� χ�%a"����ڞ??5A$�Y�<EB��i�MIj���ņ�(�|�Y��p��ý9�����o%��ؽ�C����tM�&�dB�%U��!�����`|v֤���I�'�DR��M⴪���z_-EzF@7�Y�&��^�j���Kx��utd���]�e��e���=�"]�l�M�;t�8g��&�îQ�!�����=��_y�Ă����4e����	�X�X5:fE��p�\�nt����F�Q��]���a9:�.M0�'���3����,�K���S&�<N#����ׄ?��d슼*C�$�:muZ�����ָ�ǧ�.d(�>��WSǐ%B9��G��������*6��E��ϝ\�$�6ݍK�oD��bdF��s��$FJ�Z�ǫx$���U�t۽^Y����:��8�[��1;RT�W�s���P?�����6�@cS+���������~��j�;r�"|�����X�Q`ƛO⮗��3af'�����E����ᶁ�z�:�,l���2*����?�4/N���a��F�)57����"L���F[�ձ�&� ���^"���h�f4F�H��]��g�_1��eܼ��������r���pۙ��+��S�:#��
��xY�� z�J��;�}ɱm��#j�rkhh��=��� o>���p��Ķ1�~_�ښ%�RV4C��6k�i;�v��lj'�FK��͌z)�s��E��}C���9�Ҝ�~�4ֱv�':�VS��m*�b��s��v����!v,����� ߼�NpP�3�D��&�T!��_u�ͦ��k!�Fg&	ӧx�g?dZ�_:���_��^o�F�V�-���G�9��o��\$=79Z��fe���Զ�kt@���&�o.�b��&,�lP��"z<d:�(/k=�묗B�H����ս��p}�M�˗��	�|�i���1kQ!���I%�U�oN���Fp��@���2bXL1���RGtE!NZ�a�(��۫��ڡ����a�笼Ie�UH/�Ӧ���k��yr�8\�LW���t	�Spi���������l�٩��lU�tv�9��2��D,f׶!�d]\�`Ύ��.��#ʚ��g᪪o�r�-������c*|��q�v�dɬ^����T�9��N���Ԗ@i�ɕ�2�e���傘x����\��P-L,x�\�mY(�.%4v�ZY��*z����k�X[d�|X�������׺a�n��W�Qge#`X�I�hd�ARH��d��n��;����bo��o��!��핪�s g��<`�71�;_;[B�ˇ4#,��ò3�B�fA: ��6�[�(j���V���j�9*px���>s����*����\�A�p;V��OJu�ÏC�*~;�����'��R�Lp���T]`���ba���Ae�o�}Ũ��J�|(s+u[X�����.{E���:mq���E	�s_�[	 Ytc ��x6 ���ImmM6D�Ii@~֜� 1��8��t�r1�|���2d<�d�&��b�j~jsé�y��ćB�Y��:]MN��֧�����
��I���8��ka�/���ӆ�Blb��ch���u��cg1X�!�juۍI�rexW�#�Vyg� fFs-���G�<�1���+
$s�q�A�1�nB�h�"~Sx��y�~�V\Ys}h��0�u��&	��d6أ���2�6��Y�|{���.���՟���gK:�cz��2S���ޢ
��`%�R���cnIw5Ɛ�j�w5���d����b���O�?���z3��x&�M�L�ٕǍ����+�/�1��.~�Q�*�*�6c�G<P�����\����'S\_��g�����,��N�#��H��?���I�~7 &ĘH(���u =�t	���$?p3�*�o��p�DO���7�:t�L�^$"����N�v"2�m�q9KuPΒ��5��D;��]xͣ��c@�,�J��4v\�CCm�sl��B��1O1�8����'�%:��~O���{��V������@f6�]�$��0;��U�.�2,����aJ�Fn �� �AiG �a�m
w������-��jG�ڏ�-��!U�i[X�V:���� �$9������vj�|�_}.e��ku٠��D�K>�ZF�9��i4��˳��k*0�l����a�dٍf-7@;)
��7�'�S�Fo!U�^q><9�iEK.Y�H���S#��f�Z�4̴�
���:��i]4��yJ�1	�/��
ܙ����'@i@����HK�߲�
��O�O��n���=�%��wn��3��n>������+̀�4�葔���(<����T8�%��#L����9�C�����lNe�Ƈv���:2[�R��lY,!�Dwa�)��|*"�e��X#l����bg��o�E�
A����5\2�8��_��✤33����:D����|V��731��y��q-�MR%�(fߵ����}��y��b�~��P$o�{��@)*�;��q* �g!��ܯ�m�ƹ9���Ty��G��fr�y�N��o�r��&ֹe���ޓ�s���x�Gl�	�,ًqQD�w���KXyF��l�:d�/��V '�C�?Y�s;�֋
�.��I��(��6�N�xp��������]o��l�	�`>k9��BJ����Y"5K�޸�'�}ێ�}҄J�+�������or� )��X0 �>��k��P]�Є������Jo�M�d�	V�|.���TQ��EG�K��e���M>j�����e}2�Y
Y�v����:hw��o��.qJ��H��IŰ�\~|�.^o���k��K	�M�"ǹ��}J��{�#�!�!�_$���B�'Y�H{NW('c���ѳI���f�bW��k�>k|���`|��i�7��q�\���R�J�/p5|��`���ʸp]sE�
�S�z�,��Z������@I��}�?1+(�.��q��A:8*�}%U	�T���}���z�)dWg���fL_�V�ѝ�"u�1��"v6����=C�(�s�?�_SWk꾋�M�f�O�]2TR�V ]3jkE#��hkK���b�S�5>/S�񆦏�@*��lt���/j��9�i��XG�]H��]�
��D�9��έpo�����$��X5}.��״��x���5���1xX�Q�ĸ�����ɶ��hrt�V�Q��d}�L�o�f� �o��ܾ�e,���EZ�}�YD60<�$iRY@���4� ލ��A��a_U7"rV�@E�`�#�i�Lzn%6YN� tc�:�Z�:��Du�y������}��7�Y7��`����4�>ӔO�*�Ǐ�m������N�
~�Vq\�`�ws���-����=��րi�k����Q;���Ӱ�q���m�)h�Z#}t�|6�v:�'$U�/o��c@�8$�x��;JU;��Ӻ��a�x#�2��=��|T ݣ�?��+�(��:e#�M����q}�3	:L�I�-T��lA-ʋ�ꌰ�1�w61y�Wok06$�+Z���V���&�`�c?����#BL�Jw�2��c�~�exs�({�6/p�S�P��+�����Q������G!�?ώ��!p�L:m�x�Pw7��(^����r�#����{KL���:��K��
z[:,&�%)�9�lW��(q8�&%Z�J�S�
bU��t��l���wrՖ-�	�IF%�#�����M�s�'����&���y�lX}e�b�)�����,3�U��[�S*i���m��Q	�
�OdGD!���bEj��+wh]E�'&�w誥��lC�C�c��[���Y���:s� UW5tX��M^b�N�.~��ȉPj��j)+s��Ŗ׫ӅKpV�R���T,%뢧�������"�A��	��G�Ȁ�1��[�yfJ��Z�T���-X`z�dD<@�&�Ư���R_����$�iF��SQk��kT�*{$��E6�кgv��~�W��4EG=�oW�<CXl���1�xl��T�G��ADWC`���Q=n���i�*�&��'
=q�'�霡�w@Zw+�x��^��6gl"jSh�e�q����i���eՑ%�¶WA*W6�a�"ȵ�bХ4�h��fy�溽��X��ĴTZ���6�`�Z�q��<�Ś@�Te~+�2�͘0���^��S"����S�;
�t����t.�87���p���X�e����²�;/|��t��t�#&�F;���
�nJ��O�IX��J�2��9����o�_�L��E`��8�1�aq1���?rF�}$(+=��\�W���9t�@�O��A���̓|��2�@Jd��&�Y�����4����IwI�t���gҢ��-<o�16�Q&�P����d�<k��~H��*o͕�8O�+�V! ��1�ʼ#w����3����ʽ���O-�R��1�]��h����ڣٺ� Z��L�ˍ�~��2V�?�b��-�T��{��~�A����z��(^�������g��[�q7P���;꡽l�� �F�t���) �GIz��h?�S%��&�q��SU}��ȞMA-C�l,��� ��F�y�|�9$(�Ћa���(柸2 3)���1B�4H�H�$��=���3�{�`���/�f�QS)��9�N�'�Y�@/����T�����cY���ipfEA8�(\�n̻6]H�O/��q�.k<{C���@�&�����ݎM��GTPy:���st��ߗ�s��b�j{��g�[�+3pcb���Yv��;kL��eH"�L�@H-�pqFU�5A�f��>LߎI ����� B��>��'�f7�7�y-5��^k����:��@؃�V��M��v�B���'��j�C���3����[�F��[o1�LZ�Ϳx/�L��y/���>���vܜg�ʎ���&:�[	gv�� >9N��!P���q�����A� ��~�i��aΆ��W��ˮ�G���{Vw��ÕD��g����-ݻs�N�6�1��=���h�%��F���3F��wz���<���"�e�g�g���:}��w`6��X��8����=)w4���j��9���a�:��=�K��n�]�ꝣ�]	���&7Q������=6RJ���%�!��O�q��Ku�R�!rUȟ�
:�s}W��;A��C?�7JD^����)F�=�]`3�:lW�\�?�b Ȣkemn��ҏ�`��a��tԏZ��-�� ��[�e��������3���G�d#�&�i�<v�U�bΕ���k:ɀ���cbf+�ӣ�G�(����߻�Y�Ȼ(����C0^%���E�TW�#w��A��[�ۭi_\a�`�}�Y���d����F�"������s��t�f~�ׁ�)L��o�{XU=�ڛ��A�r�����Х�m�M��x�/����Zg�g�S-�$u��5��{^µ1K���w�|a#d��	�߽�^$Or�y��+���W>m0N���}��e׉��pU�T�$K���X��i�j�I�o��?�F;n�o�R�}�m�5�ۣ��]:2���/eW�޵�Y��2��r��~�<�\��e�?�	ga�է�����(�;bۤ\(;gϟ��5F��YAM,��/�p�g.`YfХ<*��(���RT��㲃:��7��ܽS���o�s@�>T�Qg�EF���U�$'V��Q0~�d!��<��e��$ξ�?"o����)z��'�8�^��i�=�,:!�T�TrtP��!�PJ�d��]�^�V�������I�T�
��)�����N\>Hrr��5R�/�������T����,��_�P,�>��\�B ~P4���ct'�-o�1�c�𸜎 �����:�~�4�Be�G��^��@n�x�q�^�VRi	�R�u�X�Bx`]�>�%d���1 ����S��`4%hjʭ�e���g�hf^�D��.Ҝ(�A��]9����Ƌ�J5�_E`�����ξ.�������I���lLFC�rh�kS鄱��خ�/4?1O���Է��|�������5"؏#�o2>3b��8Ӕt`�G`Rdh�R	�O��ώ��Gj��M|g:+:-��85�8�ם+-`
����/�-��Okf�Y����M�ip��d�}�b{L�g����\`�"^NV�*�j�'^8Ѝ_�����|sX�Q%[5�E|�����2zVH �r1��DT�Cg4 6f���mv�) ��e�p<�d��E�zi�?���i2��r�.!���{2kG8?��K&�#��}<�Ƅ���$M`��U-w	� V��/��t��0d�!���E�s�6�J�s� � n�k�!�FnJB��CG�HQ׺#[�~=�)�	-cʆU*�?d�s+�f� �a2T�+j�l�r�|~@Lã��x���;�)�f��2��Q�wT��,L�L[9WH���Z��X+^�+P�	K��kE��%��i���M�L�FP|�h��D���u�<�?�Bt\ډvrW�.�z
k,]���?&�ϔ����{7�<�_�@\ɵ�+���S��o9��ڍa	Y���GF�9�o.�%9�fèzk1=�� ۨ�+�.Éd�[���j��	��M�rf���A����F��!W9|�G;�u�8s&�,��$ъ�tgs��Ъ2�Ks�|��p����G�|d���_r�?כݤ�x�� �2p�_��>��`��� �� ���C`���Cü�"t�<RA� ��gb<��za�tR1*&��=܆�'�ϓ�9�\p����o<9�H���o��hCE؆��u;��eh�-&z�Cd��Dܗ��^�X{i
�G7�1��ʵ�Pzˈ�Gܺ�Y�_Ľ`t�/w��A��'�<`�(�Ĥ�U'�2�� �E1#ܖM�ܒ}��D(�Y�9DU�L��	�p�X@���R�E7@N����\�Y3��iw�K�����Ά�67oL�ϑ�nw�w���@LD�qr��g�'mI�L�Ou��Dʍ��K�S=�뽵�ևn�qmL�A>jb�~-�
�g	�\���{K��=����0y�(���] ���N��u%�!*�{�Z�����"�GH�==�=������o=������H5ۅ/�&��H��@��rӈ�i"�~7���Jf6��>6�H����^f;a}��
��@��w���]܎ZBi�:��rי|���a*�o�T ��vz�aC��̻�A�a���2����\^o��?�*��>�_#����R��ГY�(��N�����9-�ؒ6ގ�
T���5���+���.x�6��>8����Ez�R4�*�J�Y
:t󔭡
x�MQ����Kt,�I�&°Q`���2�GB�K�Z1╟����xgk�[�8<^f�S9���=���K�=�84�KԚ���+�M�ax�0{Q���Ix���Se�N5�)�1R�zW�����]��xs+F�z"N��(c�ڛ��'�M6�����E�R�~��N�9��&@��hx@�A����)E���CK�E���6]���ɛ{���^�"l}�? �)������2�Q���I�}��MY���b<'U��"�Yܭn��!hN���kJ�v+�va*�Ȟ=n�E�:��t1=s�K��N7b�T4��7��W\N���w�=���s�&/�#��L��Iq3�ٕ�;<\�H�zI�?��p���h�͏�{)��!m�� ��!���ݝ�-���>�����F(�/Ij),�ߣ�R��	տ�����HQ��>ˀ�qB5LX��8E��5+[x��7���zy�ǀ�L��ښR؋IX�	��3�F+��z��S������i�+��ڳ���":�Us �����B��0�3�bB�����Q�����<�G=�0y�j�T}��[J�#zm�#��n*"'�X����t��_����>X o�~?���+X��|�n�>7Ɋ��n��<���4�MU�+'�P|�{�qg����qӘ(�ap����Cq|�f����'d�mQDIGc]��b�x��0����pQ40r��*+B��ܒ�!��"��U^H'?΄)2l�t�V]jUG׮c*�Ju�=|f�*�:P�@fj������TZ�j�T0�bv��3�:#l'�}����C!�)7�p���3�Jތ�}PE;�޳F	���p4g5��g���%�kA�Ee��5���������w_m���>.|y8X�d�31�<����8hX7��V�Fb���� ��7�г	9�M��%1ü���J`�A]h:� �S�~E�3ds.N��H�%���y�5(N�IP��B!���l)d�ɵ���E��*�S��J���qth��jV�	�=�U��@�R"n���;�� ����o}p࿋[�Pq����NFr�D����~��p��[�Em@h����e#c���,<Q\n�.���X���jO¼�
:Ŕo��A۬4/T�S��`�V�`}��c�vg�X�&�Ab4;�Y���>v��S�"�y�F����y���{�������ߐ$��;���@�����3pQ��2���3����_�$����Z�;�Q�l؛b�<EC��,�J��� %(*96�JM�ҥO�m	����21PK����G��p/�K�5�)�z��vݢ`C�]���n�[Ң�(��U��;�Zxz���B�8������F�t&C����
6�)����+�݁�+x��tG���R�.���s�Y?���%��a7�X<�b�7@V����9Q��d���}�Rݡ �M餲C��J	|����5�?ACH3��B��C�&� u���i�Ŷ��)�����4�[��pk�bX��8��0���@�`6�+����?:�K��r�ԧ/���Q�Ĉ}�O�Q�\dW�`�T�BȣO_8�SĽN3yAJ? ��m�|�)<��o��`�'��ݫ�uIgj8�<����tZ���1��S��	�ח�0c�_�]{_�lӚ�KCL�;?�&�2'!k�������wm���������q�3����5�^K_�t��#;jM(h����H�R��(�k��l<��B���ѤQ>�� r����(����Zo?��q�	ĪfW�Գ`��^�
��������tQ�I�s�b��p��Wr�2�����|����Oٟ<q;bu/N�������>׊��M���:;���*]�Z�LН��zg���$�B]�|�+���T�-hP��(��9�|�&�kc��06p���`Q�C9K���et�����T�[�X�STsS�͚'?�^/��2,�Ll�_�O<s�8���c��>_0��)���.�D�yrݪ���qq`��Y�r�" �?���ْӅ
1�ex�6�E`8��G��z����L�-M�cׄϬ��7�u�~�J�f������̙����M��\���iM Ex1��͝��A��9X�+*����5�e�G�8�р.P��$��	����^a9E b�Ұ*�-��͙��+u�
�&�s^�ӯ��7�
� 6V_�8�>�����`E�V��� DH�`Ip����y�����D!%`bV�lż�c��d��!;6�˟�K�W�wN��Rt��۶��A
t�
�#�G�\FM�.��O#<T�6f�0`���`9�����u/x�Q)�w�\kB���u&�, ���Ss�:t�#�7jg�����t�9t
������f;d�23T��<��L���L4#1����������3�"r%[�6aK i�ݻ�ʬ�Q��K��*�d��)�3g~�E��@�������h���T��٪w����odTP���;��s�n\`t8�x��bc�2�rm�DD����(�M抨M�8Y�f�r�߯��$\$����gvL��F�yi�e<�VTG]|��~ޱ���y�r>�����ɪ���T��X��]��+��!1x+���a��>_M�U=-i"�d�d2�a�9�!s^�L�d�ȩ&������r���˱.�C�"�N[����G9Ud���~�����Z���ba���扐ke�wc�o�?slC�� wI����GG��W��:�N�K$W����$f47�Q�k��K�i�+3Qha��~~bcR��Ga���fYR"���O���Z�(�q�K�Tߔ���K��y�Wh�^�Uġ�$i�ޚ�-T��7�\�s���ؑT�(-�S<d�/�%p�G���@_��vw��q���Q0�[�ߑ��
����	6<�������f�����|��>[�O��a�mH���-�pk$8ډ�0���rI3X�YV�ʴ�9��q���B��QK��I���o�ك9A���D�#��# ����k,B�×$AX}�P��ki�C- H�|��0s��S�q�/��{B$���Mj̎�؍���&�O1��;V^t�4���t�Q��IY��v�D({�wQ��Ct��J⥹l%�%%�#��x�g���)e1v2w���̓��E��G���Si���V���,}u:p�Y~�jM�k66=��T���W��<����KhӟPC��; ���D]�/t�j����"�%��EchSh���@�Iad؀��A@��Δh�TH����T�ZY�'���G\���������S,�*B.m��1��K�����N��oLq�A�W��e���S�-����)yeq�$��+�N0�_G&�n�	 �oGJ�X���e#��	+��p*����Q�'�uY桅������Z���9��������ʇ#�*�҆գQ�F+>c���X|��>��O�u��d�x�{.�#~��,'n0�YR?.��@��k�������]���pF���q)��=x�VpE��O��_f�,� �����#B�!^�K�A�I� {����h���J�e�]%�Ti��g]t@(��L�Ԥ�(��S$E��R��&�j+K�!0���
"�ٮ�����Gisu_~�w�� OO?��1���� �X
5��a�����{=76��o��}��bf����`T��a*K�`�_v��E�����M��ʄ�%�.̐wV�cC!�	f(����������=R�<)�7\�����_W!_�릭�K��6|T���]�@L�Ϧ�������ʍ�j %/'�ʮ�+Q�=�+f��c���-ѵNyX���
'p��Sl�5�ie0��@O����>$O�O���٧{rپy�nP�H56�u���3��&���5�i�O��DW�!��k�3<B	�[F`�-rw$�┠���o�Ƒ�^$���_X�}�LSAL]��އ{3���Gg��x\ �z�ҾീG���:�T�}c���R�[Ć1�ms��`�ԃ����?�}�vQF�^%LE%a��]A��pI�c٩SK��sFA�D�׍�>��b�T�Ps��˜;-e��}���4�.$����W;B${z�\{s��Ji���%������%��Лԁ�$=���]pH�@I\O��c6�S�s��]�(VǨ��� ɑ9��{~�oǆ�{?%>p��,�LZ���8�`�[.V�}�3#�IW�+V�>U�y��@����9[�Z�
�)z�ѥ/�ouq!҄.?��'���X���L�^P�y�]I}�k6�k
��;��I,�
 �dMq����vsd�O�L'�q	��Aj)E�-G�����e7�&ܮ��j7�CF�E��F������3dLt�S�e�'��z�$"��il7fY��bb%�C�EVx�$(��� S�:��Q���p��&YN���R����;B�9H��Y#�ȣj�ۻ۳�j� �����:r�B���Ϳm{ZЦ#���V�+|)qŊQ�#��S;B�쎜D��Ӊ]���O�6U%p.�m����S���x
��!zM	�Bv^)NIӹ����Q���H@~*'��t4b��s�E?��� ���[h���a��|]�����9�`we�^��햞�ܭ���7O8��
q�"�V4�|D{�n6y�������������̍�����W� 	��Pa���&s���|������ٕ���#�����Eey����Qox��_ a�0��@L'Q���F�ɕ�E^�c0H����h�{Y��c��<Ȋ�-he	f[I�u	N��_ts�@�/$������>�u~�u��������u)9p[���H���ﰤ9����b�o��&�`�%��C������dXA9��D��BP�t,�5��������o+'Y��f$�g��?>���?�q ��h�_ֻ�'�fZ�=Y�V���p0E��S6�F��t���NS����ɧ,�94g��>a%�:Ϛ�4���̙KP�(�F�13�~#��a�'�n���Ni;��	�8�v�ï�+��������6�ԟ����8��
���|W��"Yc���d� �N���q�'��<>��h`�M�:4��T���rh��;�NH=���#n��Cg�W�}G���K�hW�p��Ze��d��@<�;�F�����nZf��k�.ƛ�dp����+��Μr�VB�#zs���i��ϋ�B�����.{�v�nF�L�{��L�8��J]�ah�B�ʕze��2g\qdL�=RV�&���3t��b�mA�b���Hph|���8�F�py@Ct��^�Z�Y��#|a�M�����d��W-�ݵ��`U|:�E��������/4�	��$������ᤳhmJG?ݎ~q��m"���@8 ��K��x�N�(�e���4��F�������%�>�&:ٖ�g*��o�o3��2~�"�.$?E?#��	�*h��p2�t:�Də�����Ƒ����>�ļ�9��ю�tcuڔ��'u�����)W]� ���j�[����P��W���F��</�y�^`�.R 8�(��ǌ�P�^���M�<�8+�UK������ɂ*���j�[�.N�n6�:V�����a�'�(sȼ�x�9o\����K�Sm}���.��Ek��'���u�g,��j�,�Ψp%c��*�v�mM4n�`�Q#�n��+&4�!�uN9/���8A�숃��/)����i[��&)��40y�m|��% K���bo��Ϩ�W=�%�a��?ΝxW�DUX�5bݪR$�䊱��o.�j8�ӣ���/�#��SL#H�H���j�XH���u�e� "�e�E?)0�$���|Q�$��b��F(��I&�'jh+���q0��%�x�CM�^ 8��BϿw�l�u��-¤���v�ǧ�f�|N�&B����C�[��SU�[������uX�^؅���� �F���-���g�'�z� ;�%�;]����2�R�B�M�{p2j�ť��������jW�,�n��F�-��?��\cɲ����I9b�fbW��r~���N�I��kt	%X#ȫ��Fi��������[�k+GZ�f����A�ո��K�����~�!`

�8�(�b�'�W
�@$H�M!iV�Ҹ�Z�b��ʰF��|�	�A2��W���JQc-P<�ް����\�`?6W�T�����ǕM\�5+�O���pB�Ek�c&�;���fO�2�E���;�fpX�t]���7#�#�� ��SL��I�m��0�c^޹*����x�B��+�M��!YC⛆Bm(����M=�I#%���s��b�?9������/�r���g�٭����U�I��3�9uo���Cj�@݆ˬ}�2��	I��V�y�hV>��҆6����,Ì%sȋp��l�a�pۇ�v��*�."��<�][N.���O��>��ĝ����+�/�7�_$͚��_��w*�x�
�%v�~D.̬:e7��q$���*�lFpL��s��r��p#������͋��x^��������拳�"#�ÈS���F.SC�� �;�@�3�T��S�Ʌ
�9�7r�>)��X�SK׎q[������ �/�o(��=b;T�אu�Z���rv?���<����e�&��9 N`���/ԥ�V��I���j�^�4��}$�&��
�Ѫ�����1�{	�QL��w��z:��d*ct�\���gh��1^,�J���_Ǒ>���wsE���4��c2��CD˲��,)*ᩲ¯ #
��"Wb.����ᭋb��7ܜ�^I+$�E�nWv3�%F��	8G;�/C�B@9���J�B��������oXB��B�m�4�{��f�w(����N��3Z������820���+ތ��	��
HmL��׍`���ʤ�,����)w�0p3�j]v�lI���2qv��;�	\g�5�U->�[�M�*O��>U�L�j�ۜƯ��Q$�3���È[�W�&���J�|��hmi��w��64��oexY�ʹ)e<�NZ�C��b�-�1��m��.A�Oσ�����DY�8�z@��ˠ��}0�<*��K�b���}uu���ä�acp��y"�k�>t���^��;'�@MG(-�j�ů\�y�.� u��}��UO�~�6;�Y�~<Yr ����a���l�p����ey�+v{�1m�3Fl[J�Pa��s�Y:��{%���g�=�f����k��,�%���,���&kl���Z���lvr���%�9�%Eי�o��JT�$~,��df�)��u��h,����"X���I�9���)r�~�{�/���J�w~5��S���+զ �+���)\�]^�~Y̤�x�ɦH��򸜟bm$��@D]H���Y2b��;��h�/}��d�X�h�+��3�9O�����0xL����D�^�'�m"����έy�A�B��ˀNV���
�����[֫BX��q�@\�T����h���,�a��o���d;��U%�=`�ߗ�>�������|�(L16Z!�=��S����/�	9K�%�Y٨Z����F/완�l�u�JHMW^�@掻�(��"lS�:؇2N76oV9���[q��p�@;��q)h�\œ>���!�Y@�&�o :<E��A��4���_��h�`�����-亡�MJ[J�c��s�c��zdݷ����"���r�7��0��Fa�ؒ��U����|�y���!$�8`���#(2�Z��$��3{Jp|���+����HA
����=O'��33��+q�4�OyD�A4!3����^a�:�ۦOLqD}�_eQ�/��zt=�d�i�y�测���_VeW.��M] Hs����}#"�����ڠ����Z�+���A^�i4E��a�g}W�XI�[!���Β��u��kan������3K�hR����_=#hP�����/Qt�vN�~7�W���P�� 1��v5QhǕ���P��`zTx�s��(�t�57��K�R�e�㫳V�����K�,v�g�l,k�>q�����WF����-�,��#q6��i�A��_*��%�B*R�r��T$��ڑY��6Q��e-�}L��*U8�?o��:�?��S`s}h.�� ��L�i�p��ˇ�e�nw��3z(���+"�o����2
JȲ��51��|p {��I�~�TJ�=��Հ1:�N��rt8�80�1����L(�=�8m; |��g\���x��e���{P�y��W�)x%����p��V>�la����蔶�z<X ��7������g�I�4J� h�Q��#�f�;���G�� ���b�y��ۍMKd=�h� �+��l�	��n �J��::^Z�)'�1Z^��e�5���ܔ���I1ё꺙��
I��k>`���q�l�ʌf���"�u�1�\��ji���Bd5�l���c�	�z��2'
;�S�2_1D@�s^9�
�����F�ZW4���v�U3���x�Dҍ���]�뇌��v�(�����&���=v96�:5hT���'1���_��@�_�2C�U6^����A���{�z��0� y�71��:���a�*l���
�*k���<�V��aT�����}�G�fᐗ]4�3��� %~��c�eG�{��Ȓz���G�؀"l�����?��P%S��N_ߺ�J�~�;~&,�,hI��� 0#v�G���������zɰk7xn���A
!��o���uR L��B)|v��G6i��h�4cd�i^.�열� S�̠�����r%��bmB`f%g��(�=��8��A1o]�ޑz<<8���V��za"%�:��XmQgw8}��/�,��T����<)�㽘�[�uE:� ����#�X�1}�%B�W�L�z�����?��P v=��2�?�9�zy����j�bl&��Fu0��'&�D���jں�b��
5wT��V^�	c��J��1NM7l���3	���H�g!�A ��#���	�p��!�E�E���{\�yj�8Kn�¢�ҙ�
\ĆE].�Ly~Mq���3��L��aZ����>4*�O;���3��k�À-�P�_��jkwyj���a@q���⺪e��ȱ��+�؅�-�)�N7;�pښ{eW}�pJ�s�+ȧu�?�@�j�M	�S�/&��K1_.�bx���-.$ �q§J����4'�ݵ����۹YP�"u����� @�hn�"��e�HE!��f�� c��\�i@&&]���W|��jY-���u�0�8,�h��i��D�^R����B1a��R��P!*w��E&3yB�9�)�n�q$##�t���\����
���7S�頡'��5!���&���D�q��@,�?3��:�y�V��"lˡP�v�+����V̵�z��y�´��2[s9i�Ï2��������ק�U��`]S�\�r~/�f�D�A����cS5������^��I��+xK;�m���b���/�C�+����U�6w8�m�<�1������P'.�k@1O;~���|�>C2]ε��Z_��z��ɹ/���C����7��9�`���1K�ϳ!=f��֚	-�
^�5Q��V��#C��Ȭ/ӌ!l<���pB�ۏ�d.�e�֮S�==L�]
� -4�����5rZ�ĩ{�j<�uh���t�#��c��)�GMŨ,��!��ITp'��8�x���,>�������X��N
��F�Z���I��4a+�I@���� �*>i�t���8IiVE�`O��{�\�c���V���CF'�&u-�� �y��#B�IN���s�� �QJ�o�к�jq��Zr4/h�E��P�`���X^3`�{h�se�Hb����|�{�rr�`���p��q?���"ۭѩ�g@3�x�t�lW<���<�&�/'�Y��J��vÁ���%?�lz� �%��� ��%�L?�!X
�ev%I�*,�ׂ$a��<1��Ԗ
C7]�n��i�p�������;�r�ȆO�i)/���5&��xy�/�v9���"�-6o�rT���#H�p)t�*e���s���<�M5m���������x������#�<@���6,�/JZ���P�}�۵MQ����Y�ͱ����,؊�P�o]���a5�c�o��S��&�Ei��aš��� ��2k�xþ1xk��]K|�I8��T��O�%��8ߎI:�?�e�C�9%ދ� z�rL9ϰF(�L84�,7�d��9|[�oR�u���>���8��h�[H_�L�i�_�I�,R�ޑȂ���A�=#�-���)qY^��j�Z�	p��⥤.������C���~�b  ��Rl���n�taGk��M #<��Ү� �'>ڂ�-�����ݳ��q��O��>�C
���:�ˎ��օ&"�z�q��O�tN�Z���}A�.���r����z���+T��M��D`3`��	�G��B�:EA�_NR�M��8�@�g�[({��&{���0Ne����k#�8!�+D�ܼۚ����%��z�=p�׻�H�C/�CP��"㬋/Z6���\J4�m>�Q������_ꍂ�N������b'^0r��t(�R��-ĪC�ǣ܃�{Z#�8qM)�^�)XH�����<���e3��|S�l6Ѯc����������h�B���^H�����{�H����o�����E���s�󫯻Q�'�s���_����z^�Cj#�luP����9K����6V���>H0���z=��윲W�s�h'e�4ī���L
���(W#M�ǖ�s�%;�j��Ӿ���:�n�p��������ᮈ�8v8C�^߽�{n�>�Σ.[�e0����K��0q��"�'d95=�:�v�)�-�H d�y��#V o���VyC̝V#��X#h(/T�7�#��%�L�`e��/�_��bIh����NZZiS&�"�VDY�-Ǳ�=�󝶛�@�@ ����<c��
�d ��������/���|^e[�% �L���6��F�}��@�nc�[�0��;�W���q�+0*pd<��~�^�DՎ��v6~uS}�i��f��5)�~�~$R�p�-�:^dX0���X9�ZW�Q�c�B��g߽\��d�Oy�"�u��gi����:~)�ز��8�Y�1��^dNbkC���~Zz�se��C��E�[[�^� ����4�|�'$]N�/6x�1���� 8�Ins�PN�o
���t����G�\v�z|U��.E�[�^�*���-�J�Ʒ�}$�*�>&���
հ;#Ob��Xࣿ`�E�Y�Ğ�vx	�Q Z�wE��4��rf�Peʕ|%��:�����F��'N�ׅժX��	H C	X��G�ʐ�}5!X�!�B��[7m��Vg�n�[��A˳��(@iX���;rx�i�4v<d�"��o
A/y��+�m/�#٬�|�����7��z����7Ɏ���ڜjT����e3��RtZ{��ɥB�챖�be��Gd!R	����g��Qr���FY����u�]�{Դ��(���̺a�P��"@��^5���\*)�ƐvW� �^h��,���u��E�㍎Ѓ�&-ha5�_�C�8�K���N�h��=��3�=æ�MےӤԬ?�	��]��tc�;~��CE"o���T�K�I���L_��66EDZ	5�^]Y�F8�įb�9uJ��%��d%���?�\�{+bYX:����r�1�8[���
�?�Zu�ME�~֬M�"!�%(��xD�̽�L��p ť��Sq*��G��]�Q%����I�GF���>W����"0Y��^����S��ޔ瓂]��r��g�I�ɅvW�� ^M��z�ZL���0d�5��
;jӤ:,$$F�X�c��<	=�|��Y[7�.lu*>����k�L���VQF�K [Ԭ ��{��y��Q�{����YP� @� �#�o�f��r��7#]�B��t�ҧ�b#ׂ��Ĩ���]H��HY��Q>�f�LF�`�6i�] �g��M%!���5;V���0�5��*r��M"m]6�0(�q6�Ÿv����oܦ��io�Mw�5�R+�Yc�����o�,�p���U��R�ӷ�#H���~�:�l�j��R:V��-����c�V���l�b�!�*�=a��<|hk��Q���(�{i���=�e�``眧��^<9���<R�UՏ�������h�!��<�UQԜ�����]d_��7.��|�i%��?e��Œ�|IU�9jh\I?���$W5�
�1<K��f�3Y"��M��1��"Wbkiy?����Հ���,
�٨LzK5�q쎁�+��������k�Z���6�1�uϖ~���Y�ƹ~yF��8�FC䓧��̙�:���i��|�����a%�ҙ���3z,�j=�"TK���O<Wp�fit���;$�&Ԩ*r�:�u0B4�F&$���-�
ݦM�Я\��%-ud �50O�l}���XZ�Q�����jƓs]馌��L�}M�"N|�[�s���Lu���P���oɧ#���R+�x0�|t���"����L�c�wʦ�ܼ L7��@#�x�{zL�������Mʬ�o @"7�Y�Q��+��V���]+��?�w���f�O���.s��.�v��)s�2SrR^�xP�/mVƥ|��5~��Ѿ�%�"b�;+���Q�<�|fd!ϟ��m�#��/���Y�����'[ؔx�$v����Ò���C��EseK~_��s�m5�u�F�[�G�ݢ�+$Y"a�d��獉��?n���X�Fr��6O������ZL��u��֕������0�����/��-�3�тl_��^�{�f����J�W	X�������}%(�]Ԛ�����9���N�r�.m�*�p6DR{<� (ͪt�9)Nr�am��9�ko���Š�x�31��k�,���CW�!�H�;��g�8H���̪8A�~�߮2R�:=Jx���%tpP+���<C�)��0cK�:S4�3�#���Np�n��'�`ї��J�w|�t��g
]� 31dTÍ�h!�Y���3��h���W�:<���6w����?V�O��������f[f�.V�9�s��K���>���Q݃� �+%�;�{X^��>B�wJ��G�hT�`�4��9�j(�m#����3ʚJjso�᧢���a�I�kݳO��i�%�T^��sK�s&V �ڴAo$��'�� �����h��Gf]��ڄ�\J:}���rA���?#����/�/�11��*:qG�m�������>��O����Qw�[OhQ��С$̏��l|[�.�o��h Vsϧ�͘�6
r��j��`����W:"�H5��t}ud^�1����ߩ���&6��*÷�@��К����1��M4s�_?���Bז�}��t�����n�;֊���Lhߘ�� ��Y�"�����%��,d&jl��~+U�����+P\�q�@>��I�\.�L�F�%���;i+QZ8���mjO�YjB���4��R	����(%�HB%0װm m�~Ie$X>��)#19��O�Z��O.�����JqL���zѕ-���H8f55<:ݬ�p2w��06���2�����1���Eak�܊7ȘL1R[�ܿ[R�V�tY�j;�F�d+5�S�l�z׹�Ku9�����M��E�
�p-�i���#��5�Hѩ�j�4�_�!jt�����th��Cs�=�FiyL,�ӯ�Q�T6���~HI����D>S��Ն7��]YAn  gk-��/�i���c����/���@s���l4t�f'��6�_���UM��'��Pt'���U���79��=4�9a5�$.S `	Wwh�uf�?��/ܙ�!�z}��/�����%��R�_�F'�m<�^��N�����J*�I�;]� �/��1+ˊo���\���-��<��`[�h�Ӧ�F�sl>���,��a]��{�����@����cp�>9�E��c��_��iPGD���q�D�M��SR�����Y}u��hW�b{4�5��S	Dᅈ&Ze���]�M��n.��n�Ч�X?�I1�4?��ׅ	���*͡����������v�����}���,��靺���Q�AG3���x_���
J�Emm�n�E����3�X<ePL4��Nmt�u�8��rO������o��o������u�Ǳ'�	�� b�Fd���>�9��K�I�>4�Ҡ`o��
:Z׊�nQK��/Ϭ�r"����$��h�����s��[�o�o'�*�.]�j���b>'CJ�C���dJ�u%�9,C���d<jc�-9֍�3�l��[�yk���x�Lu�$c>�[t7��+���=�˭�w�O�S	��P�x1B��ć��8� R������w�f�������ggX�$�
�OŇo�,Rr���FH�+ω�\��M�,N�Cߛ��ۈP�0cQ�	
��YL%�ἵ픬��z�9PzS�n�>t���n2fV����4���^���\��]ldZ�U�f'�4 1(�sػ|��\JO�e�v$!��`�y�e��ƿ�h��ɯ�G2ߍ	����W�����z�	�4�f%�9�U�٥t@�UǮ��ܓ��Z!i�Vy:6�_��Wh�_4��*K��� �.��.Nc�S�~�±C�lw,�� �
1B��)J]5{9��}�~��ɟ�-t��Uߥ�}/\�@%���i�֫9����z��3�[���2�����t7�;����(���ЄM1�՜G��x�X���x�]�z�|?L��2 �����*�v�0��3k)��&�wq�f+t�n"SO�ʪ&�J���HӾ�3xTW�� �X�˞Ӕܦ�>�����u1R ��������:߂S��y>U<�6�mT�9n�'r��Ot	<:d������JYT,�&��~^M���e0Ѱ�C@� ��-0bc~dS�Yf�\~4�#:+Fp�]F��xۗc̣��z/����߂�T" �ϙ�n�����D��
ytp�����G�ESy��#A؛x/g�e�@2�Þ�A�	���5]���j�"��]��'ۖ��9_�'�0�)'�<���p
N��T��0�(��t���_xt���YZ��N���f�-'hǍ����_���R�W����z��ڻ�0���Y���c�>Tv`ė�	�����
�������m��P����{��U+̓v�T��9��2<�N�