��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��)sZtYzѦ�#����������^{���f����@,�B���ul@k�"T�z-��0��{�oQU�<cM i��CV��Ǣ���j*��>3���B��1����ݿGi�b�2g��8��H�2m��@�}
�G%�p���.�x�T$X�v
��;�b$C����f$����D�j����+���DM�#��k/��|�S��p�k�ҘMw�����t���3��	�ΆLww���LG�\��*B/qR�n�d�"O��
���<�[�ٮ<��?^�+�#�����\`2Y�Ϗ�cR�W�G���	@oU�z%�� �˗�#�fŪx��>��1=��&��mErc��ϿY>g#d����WQ��Q��h�.�8� {J��=}�17=E-�挴ە&0�3HFq���F�W]E:ń�{�B:�(��=Y��َ�o5qxE�~�4 %te���s�6cܮu_�b+�K�s�_H��м����-�]�Ô9s���f�Y�5@�(�:Fl���t�����"���s,*�D|�ޝ�'/J���v5�������n���4��>� W����� ��驣�֢�7]�DÚ�\�y-DӢr�X��5����}'�E3c�j��6�۫�����0D>��Tf�G3�>�~�0e� ��d'ɔl�GP�j0d�S�T@|�;�'���t�C����K�j������E��n1�$b9��z��!��o��1V��%��xh�Xy�����B"�u����hk-)���7�b�ψ�V�*�㿓M�}0K���.��"����6�4�yjᔌ �a�o��������6�1s���S��.��j9��;�;��|K��Z�n�>-�����o~�ɪ�`^����9����/I�g�j��x���Щ�7�&��]�2[�y�T��س�� ������<4�X��-j�p�E �|�
��Y�_����}'�,���Q�NW^���w����U >0QU�Oc�>���6>6��7W���tU�*a�ֺ���C����
2�9S����9���~ �`���ko�s������` �$�jN���ӧP]c'�I�H�9�Y�����ܒK�c�S��fp���4�h&ig�����&V�X��Lh��V�J)c�M���K�!����TS]�4�"���i�y�Ŧ��"Z�P�����^u�8i	��-Xx�O� �B�T���4���Jc��J�B�[L���%�Q��Ms{�������Q�-7�E�6���, ��=q�^2,�#y�%��$D��
�/�	��=��e9����nrV����F%�d�3��/px�3��Y�n��B�y�|���+�#r�{��3������uqޔ����J�7d[���jL�s=�N�B�;-~U���f�<��5�64�,E��O=�B�8�uR��:+�ӂ��H�h��H}R����E�Sf��~юr�n��*�_�������X��AӪ��#xhH��dKj�E�(��q�E�k�W�]T ��
'UZk n�,C'��J�7�G�I�	�^.��3�LA�$uB0�i��Q��pj�w��#��wկB
�ӊ���*����1M�髾My��O�vp�������m������֗;� ׅщ%�zH'�śs�q/�M6��wT	ũ�'���t��:��5bkq�'I�o���"S�A!%pQ�8f�O*d\������FT����.p>�^+�ї��^EY�=5dޯo���V�BV�"4�N;�P�ָά.�.gl���kkq�L�t�v����$����6^E>.G�wL���+:�	K\-�.��֡�ԁu�u]j�#&Rt8��b^�hP�_�p�g.���`s�ѭq��)9�m��8�W���m��v4��\sz�,6�>h��-�a>�2��7�������ɽi� �).�o��0��kÌY�ؙ�`����,|�=�n��Ղ��J����tdk2��Ih������8��(=d"h�l
9��~�[�H���<b}~_��z�By �<׿��b���	�̷O�^R�wg'�N6�%O���)����rJ�#��߻]�[�1��Cgy�cƢ%E�M�����qe�ǽ�å~&�:c���sj��fY�?�7��|v�i���㽊o��pgk)`>	۫�����lL���[��ƃط:g���7��"��<��̤�~�Q]s=$��M�㞧�ݳ��I�f�Zh��iܭp���Wυ~�i���_	��eЮ�?�/4bl	��Jf�5W2
7vD,¸��Le�e#�c�FrK�=²a���}�zv�N[��h��<k�	��v�2��ʺ0]�<�z��$�%��<7ӂ5��o���$�.8�IO����l��3P�Q�be����9�<���+ܜ٧����"O��ǣ�T[�K�N�3M��(�1��m�����e����up��������?�#��h:CU^:$5��w�I�h���:]ֳ̼֯�+P�����R���k�D�%�B{���좳8ڧY"�ˎ��r|1/�2������Y(�y�̭�c#�㈋����AKQ�_y^q���l�U��ٜr�љ<U�&,�[���}y@{�b���D`6��)�P���/�~bрW�%�u����>G�� E�V�>�Q�������wC��
0r�@xdp������4j��(�� |z�c�w��	5w�V^dHKu"�d�h?#�X3$�eb�&ϖ�aV�nT�)�O��o��iXn�H��
Ҟ���`�T��{=H���έ�#�[�_ZҦ	)b���PґH����n!g(���M^]"
�t=�t�s�AV]�Ner�´��1{�HcPJ
3<���~-�}��m|�Ky���NO��v!�C����eH�J��s��}�t�Ƹ���A�S�JE�:T1��Еn��t(a
���ɨd��͋��*���Gra�C#=!5U���&o�<{&�	����m�3MbN}�6��I, J�j��Lf���y�GZS�a�����$��,x���D��3��O�<������|<���#��m0���)O6%)�����&q�ɊBr]�5vh�hɋ-X(��d��M@����0���Zh;�7]i�*�iu�@���Ĳ��3a(Oѕ��L��+HIP���EU55h^p`(���G8	��x5���Ȟ�M��6���~�gF;����9�i�QL
�dؐ�Ou�A���A�ʘ!s�:b���\���Ge�����!
}fy�1+����Qm��q=������U��C��6{���3]��<E�}K�V���	B����>b�QM4Xq����@Sy�y�mVڏS�Um�L�K���b �kF�KՉg	5�$�*f$G�BKސ�U�P6�j�8`bݥn:$�ӹ��!3�9K�V�6�x(��I}
,th�����l�H��^�hʒ0�� B�Xx(�r�L�x���@�#<w�8+���ܣ��o�ˉ|�߱�/I���5cOwv��\�>N���5���%�n�~�n}�{������Y	����Hi6��"��p����_r�7=y>x'��|h�c)�4촖�˯�닕��=%#t�jm�[.�`䑲��մ�J��O�� �_�L��!ϝ�<(�J��Uω��O����</�6�������0�G�ba��'!g�
����X߫O�����oU�x