��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^������U�#R��y�G�g[}eZ��n�G;�ieY≘�`{�{�E)2���9:q��e��:V0���	�};�o�h��#[NOD_�ZڅI� g8���+3�@˕�򷧤0�d*A��	�;un�l� �cQ�i�w���ii=��<K�iI��� z[��b&�(V��h�|'4�^J	�ó��+�K%�̸F�7�6/�:���	�m��#)��K��ӯP�]��J�N��5��X�����2���HG���~������걺� @��FjbZ���闾Js���pu�W�ZFC�1��[��W#z���o�x����g�ƟM�уg#ד���2��둬_aIC���6cöyc�g�Qy��;5�
M"��r�Ţ�,Y�S�?TҁI���������t�\���N����Bɢ��;y�_<�u�98�uq����e�������S[j�>�>�t����W��}���-�͋��W��&�(�:��������� �������¥�P���I��f�%�c>�/]#����;�Z�O�ڴV�����C���]�̒mh��"oI(�Y]����>������p:35e��I�U�r�8r�X��Fj x�%e���t���BT�s�f�(�V�QH���f��h�ud-IϏ�-�Օf�Cq^�w��ˤ)!�2K@�E_�0-�hq<L�$~��i�ÁƄ����|���A�����D�Y���	���Hh���QW�eW�b"�O�#P�~��ۏ�,� ���,���hHF��0�?0�"V�~�f��x�C�a����M�"��f��TO��z5�FJ�@X��V�����|֢�H���'E�Ğ
V���	�%Ȯ&ĥߜ����B[?��6�B&ƳT���R8;�fHoM��*����f+n&B#�1o��ʅ�!�e2��q�cM/���x:���RRt1�5�|
�i���-{ǿ��`�����a�[b�{�����®L$߲�����5O�B���x��ك@����A%�s��6�3�EU�����6G����8��v�.S�t;f�������>I��O4(-y|���`b-.�;�f��e�a��*�?��f2�����%A���\a��n%��?MGא
���h���L=�������,���p��T���j�6�����E�3�̻��	$u)o��~;��k�ع6,����G*v��� �P+�e�^2�&���­�YFt	"�$��P�����o�K9�=�C�/ˍ�_��@.�b[d���S_���Oi���IfH;������W�-�0?L_��0�S�& T#Q�QX;�<�6,�}H���+p3�c'��	�+��Z1=b��)OK��<�M�}B�HuYg���Ƣ�E��Bd�Jo%�?������ߡZ_-A�/�^��qP�e`��t�D)Xt�����x˭�����`f ��(^� Fz0���j���{��U��պ�kP:U-̤l�ޕU��(�#�MwIӣڵV˒�0,9t����P�ȃ�ݤ��0ĭQl��Ꝯ=Eo�+/0��8���p��5����ж0�Dfkq̮������aD�R�R-��7e	=�$����ծ!o�1����B�75�0s������Vq\+�1��)|٘���܇�8#��i_0���]���E���!�D&�S/%�8T�Rd���ƉAaM
�^����O�\
O \�AN�ڣ�=ᵭr	�#�V���q^�*�7�]uB-��A4ʓn&��$���$[�_6^�����'1��0,�[UwYE	b*<O杷�C��>ٔ���%n����_Lk[�����b"r%��JZ���w\K'�b�$A�i|�"o���"-I�W~�O?�5�]�f�q�a"(��-���58�����V�����8�xQ�Q��r*���#|������[Q���IM) ۫y�c(Ѭ���۫�(���J�7AD�)d	]T����*�u��"�<,�Jdun=����o� �a�-WgJ��h�s�,8A���s��3�۱nެ_��Un�z��
Ӌ+&����)!�X>KH�D��woDMr �ߖ�D=l(v
ٞ"������ұz���.��x��"[�1��ou��v,���P�cr�4�A�JRӅ������h�r��䪅��tw�*�<�#`
��b�oi�,*�XH�9l�E	�^��},�C��G#�m)`�@2��&�1�mN�Z�& ��bɓ����\�A��R,�7#��J
xC�L�eʪr�҅z��N���8;Zm|���˦\l���a�ج�*V&��L=�cn���[KE�;�
U���1$�̀�|��S�0+@[����Z3��l)I��&s�Ζ���&t���e:�x �|?6�<�t�?
$X&1�� �Vې1;�9�� 8^����ƀ�����,|]9��^����s�Y����D�I�Fw�
��z��cd!?�=B#]쉥%�}��zwm��j^����1����ʠ<0�h׾�ď�ٷ�)�c���n��Gܼ��T{Y���RD�\ő\�	+/�K$1��ϕm���O�j��8�%\.�{�SN��/��k��~NH�����[z���#��vj�H�z{'"m�X�N�K@P��4�8��c>��I���h]�_?>KSTEk�o�i���T"���zé�m����*_=�۲;�z��,���÷�d��@����{)!� $\F��ժ���;ID�1�K�w2]�.sp3,N;���ߜ/�Ȝ�x���aΥ�j��駞
/�\�(9��T>g�V�ai�\�	��;t�Fcl��yc���!�cn�k��e�bZG�gy:�3��)*�I��"G���8�����t�G����2L���·Y�R�g�LA������5��S�C�$笤$�}���w�\~K�3f������ӟ�p��ID��>C���@lV��ᷴ� ���l	��g߲.VȖ���2����A.$��*p�.|$�ab��I �l:C�Wc�??����Y���O+�I�Y޿:I�|H��t�vg\z�{�e�q����
�̧M�W=v)�z�(�~������1�Zf��jrf�ڹ��C�Z��BdT}��(����$����c��@�s��\�몑xU��yB6؞�4���ޤ�V�:<^��A�jՐX��Ske~)��#jn[d��:�j��-,�#��Y~�x�M��ʷ�J}���<��տud����|��/���Cq@1����l�����sӿ	��}�5���v6�=;�^���]/2�y1�jի�\�iӌj�M�~�V)1^[�fg�X�f�n�t�R<�����VMG� k�ʺ���}<%g�*�h������u#����c�����ka@���}��j����{��d�t:?pC��	؀槆1/d��Ah\c��9b��$�ʄ�53��g\�r���F���k�ﳕ�Yש�.�U(�f���2��gDVeAE<�ŉu��vEk�%>C�P���p��k�]����o��h��Z�r#T���ށ>�QS6M
���6��z�jhܯJ6ѐbT!ǅdT�.jW;�j4H�L4��ӽ�h�Ӊ�4��5�4�����]d~u-A��Re�h��3�T{���ʀ;�Zֈbf�ؽ���ȫ�Ul�޷w2xP#g_N�
T��|3�	��h���v]$4V87L}�p)�S�j!�`\]�̭5J�5A��Ս��$?�b�Jt(Fk��U����~�bP�2�ރ�]1�+�1����YwA���>3oՅ��mZ����2k��yӻ�Z�`D[փY'������2����+i?O��#v��~`�=�MWrr�a�d`��w��%{���W�:^��޸������|(D�_�Y�>8��,<�:�&r ���ؔ���Գ����Ё�a��8�);���q�&1M�'�����%�x�_�J�i�x�'�m��	us�։u�*�2���IPD��g�D�|,y�#��x�4Ԥ��t-_i�+���~_i�NU����ȋ�y��4�e������BF�����p�C@g��*�8" ���@,H�M!&����	 p�X�C��i�bmz�}"Ѡ3��L���4SU��#�/�4��E깝M| �33C�Af�c�,]��Y� �q�$S�t4�����6�	�T�WHL�jUUo'x�F�W'��P*3�r���`K�كy�S�JY�Pڪ~I���땼������\oq�����g���i.�[��'˭��@�*�hDۚ�T"<��lC���\-���փn�>�F:�jL	������ \h�yp�:V��t�z��="3Z;�~p�y�)�jңo?�S�-�������NF��a�yg~�V�t����&9,͠�	u�Ra���!�u������-CE���\�
��D�w	��NDx��p56px�XX�@<���h��
nVJAG���@r3Qdb��Fa8kE�I���	�I������R���rvj��W�ķǣt�Rڗh�
Ǜp}`m���LT�H �:�r�����AT���0�#3$�iΗM��� ��j�0SND�K̬l1O!m�PS!
��~*@����ޤ�Z/z�{v_O�,~��+��N�N����{=�j8Bu'�D��;�˦n�'k��um�>W�e��mRZ����
�:�2��ՃW@�I�|G���k t�-�݊���C��Hx�h�Pd�	p��xI�RA�5�ay�O��k���M�jǭ��/�7d~G����虻]���YP߹Z-��Ĩ	�Wޓ���t�:���57<����R�D��A���S��!��g���K����z|�,򛇅�k�_>� Q��y�C�8	a59\fi^�����rtu��H�[�v��s_0^[~��F�� ���3ß#�0+�K~Q/�p���!@�Y��Z�7��M�ze�n���,��:3�]��Ʃq�7J�ݝ��7\�Vb�ON�_����Ѵ����tpL5Vu�!!�p
O�Ư�?�N+X߭���k�Y�1��N/����Tn�[�(������:	Gl������x�����pKH�o]&�'ja��Kk�Bo�&��� �il��U����gܜ"C+������1�ڝ��ܿ����]�1W����Q`0!"���z��)
0�AN*o��[�#�uz�+)�n��71��,�\&�@%$���oB^���Φ�C� ��ɂ4ʿ�O[���������YT��2I��X��;��m>��j�L�'����q���b�M6�|��ʺkc1<�i���˂�W!���p�/+¯'c�Ǡi6B���"�*��]�4b��9��rR�v�m@#�|RXπ\~���Vb�"��]�.
g�w�S\.f��xj��;�6��$#�7`��Jg:�T�CI����ԑ� �I��5��q6^ƫ��ˍ~�@n"��ǲ�C[�[�����롐�oJ�V����O��|=�	���n�]:(&��\&C���7B�d0	3�����<��z=*���� �u}��Z|X���j�Ro�'~i�����2#���n�JLol�X�����iHEϳ0�w+9��&���^�;4>WE:����eJ�?��^���� ���ky篫�k'ڨ�	@V�ο�G�
��mƷ�CN�WZf=���3C��7��?H��G�ͮ���x��z�t�f�5��=����U �����6�c5�#$y�-a������f����O����#!�r~H�d�ը�ҺhU���ߝm�����*�,�z���3H�Z���s=G(��B�ᰗ�s֏<�t)�e���,�, X�.c�<9TQo!x�+�Vc���]�8Gᣮ���C6����K���r�m}�9t߿��=������m��E��.��5�K٭��|W���ك=�����^�/�����a���zn�Z��J�n��0��fX�Q����սu��i�?��1����`#�%x�o��b�-Խ#���3i�ⱘ,�q!��/��Χ�/�  �~~e�X�dKD.���G��Fܭ�,�������sќ����f�u�e�3�̕���(����G�E=v�-�u�� �F�2jD�\��� 6p~dXS���<S�b$gq����?`#?`������ԡ�\�5&�i�Γ;��ז�^e�;{��!�&I®�9_r��p$CS���(�	JV[��g��Ë��ᘒ>{�f�%�y�}d�� }7�.��{WU�&��Ø�t��܋&�r�s��I2���6z�p�K>m��ߝ�؁.|�T� ��?JO}M@�K���cf!Z^77�;���$�q������j�6�<��jio�����=�Y�T�XB`�͋+'Vw�T��YN��#��~퟽��H1����\�8�z�h����"=m=tJ+�7�$�9�-B�SpW`P�]j���{�W(D�WM��L�5��������q �J�0_'s�6��bW�j!�Xj�c'�K	�3.���!���s�+�ۮ)|6��t�	&� ӑ��.@z_H�7�n�.��(���͘w!�K�o�L`x�x�����f�pğ���HHv/3_|j�!=FS�uZ�f��ʭ!�Q���?8��9d�8P��o��5ˀFr�w��U���p���~S�|��b�M�Y��G8��[J4A��bar�ͺ�rT�ŀR��fC�&��/��OTOq.�3��R����PI�{��u�b��>@-RZ|� �Z�T����I?���嚭.���f҈x�����/�+��:IXv� $�D<=M���XhP�8�eNsM���Q���*��JyC�I��>W���v5�8���Kc�$��#B�
?lP|�A_ �SP�O/ ���q=J���J槱�Q�n�C�l��U]��B �T�Cq�x��Ć��ҕX7q��;�P��2s�q��_QJHx4��A-
Ce�Uo�OѯF�ġb��dc4[M��A*��9NU[Zat�5l`|,��)�8���SL��%�iw��d�/R������e�e��^�av�Fd���WO�c��V� �ۧ*�+)��
*��A,ӊ��&(E~2r�V�̹9�R�����OY�c�j�QX]͞nsk��t1M�!"����	�-@���?�_C��?8fΩ����bѐ.�B@lJg�aFɡ�=�4ؔ��Ng�$Zۨx���R��em�jLM���_ ᣵ&��L���G!��CL�P��Ps��K_�ؖ��<F3����������� ���S�a�����1e����ܒ��*s庙�W���)'ӝ$y�r	�q�Ѽ��� [*�l�H���!�Iy�p��815%��Q�0��.��TK&��s����Ҫ�G&8��0"H���l\�;�ʸ���誼�X�P����AS�C\�I�uZ${���mK�c!�͔_O�����,���D�V����Y@��k��R����y���7��R$UR=�5n`@"��a���hp5��8�8�����6�P��u���s +CHǡ&),䙯Ed\~d���E-�շ��dt�F���HO�N� }T}  �� �H'�F�4�c��oK��R蚥�\/�07,\�ӄ�}v{Ӆ�S�y��F��mü� 2EJ�i���F40����ھ�:$箜� tjS�6�)E��e3К�,`A֑G��>��>����o �AY0ӃLkf+��^�0P+8�Z1!��aG�����{"�f*��17�:A��܏)ʎ�J�j��L�%��~)�oK󨘀+�떲�9��K�	��8�J�x�Ԥ�<�!�����R����T�.6��:��J��KR��2V�x�f�� NO��uj[ߞ�7q
nӤ�^�G�ih��D10@��\6����7��pҍ~����@��O��G�7±̯��gU��X0!���Eҡ��5qO}���9"��,(׍Ӎ�])M�����#����f�k��0[e�y,��"�tx��J��}�#��D��|���郥� &#l�N������+�Q�X�`c��>fҲKՈ
b�����3u)�h��}�G2#D�������}��,������"�<�٠��3�6���X�M��0P#��}<��؟��P|��NI��n�`r�lW˪�{��b��e0t����岿l��(*۟?��.�j������Q�b���]�b T%r�;IOb�K;���A���]��7j�(c�qdI�6d��xɭ�+�ɗ(Z�����dxv��� (;�eb9��9�uA������y"��V�#t?=7.k-�'�t��f��)gX�&�{;�<Pq%-�h�=��x5�{1%���cu:�S^�M"��{���}!E���[��el7(U��>�u��#���1�	����C&~�M��n	��L<8�k#���E�S����ʚ $J���$�bK��6�w��r*��9�u��Dl���e3d��WF�oN���l��i�i?1�^CAHj����i��ai?����G�3x�PN
���A�=}����V�0S��ujg�v-��$��/��W�����jD&	N�kn�O0�x(����Fqde�#(�F(�@6o-��<�1�i���z������� [�O	��h}�M��&_��M(d���i�\=u����A�@�����݀�<�w��&{*YE�'K��œ��
��J�aR+�q�{7�E����c�K�.V�6\��Ie��@9�4�1�-�~����z
�4���V2�z�0��96�r�Lp]�+a濡׉����b�d�ؤ�t��ǌ�~NZ��<��?���=���L�#����4s�
�{�h74�B ���ט�*���X�D�p �9��e5Q� P1�>�:������'H�5���!�K����?�B!�|�rŃ_ ʣL�@�;�B�;L���BV"�v�˃S�V1�a�p�Z�x8g�z�3���&����]zN�{ټ��k�c�	U�o�l՟{��|�����V/�������۰�YZ*�eF�d�8���}��{��}R��b[z�O�/h,s��e��!�r�+���9���&��->&�|`�b:"��#K�0:��U�혽��W�ǽD���󗕅&��n>RC�Y?$L�4/L�̭��3��V
���!�j�g���j�;Z$�آs�?�;p\�h�mJ7Vuluʇ�P�е�(C/��ne��s��x���ARi��G_�N�8���*��	( �WR�R�H��Dĉe�!�2K1��Zh���IE���Nh�đE�<�!4KBߺ3��d�͆�O�^��%�m���P�>t��"\�ײ2��_\DV^��� �Ize=��|$���l�Q�5��9����AiM+
��A�I>_�v�[�sTǺAW�3���V�W��wr��^��w�u�H���R�9�B,aX�
�p���nLW�ޝ��|��c|W�Gw����n��07�N�
q�����a�y�
s��#ͼ��<��û��>5��(27Ţ*�Ҿ#���Q�7%�r����K���]k��E������U43��K;�
�Me5�*V[�43�
謒(`un��n���I�,�T���~�Xe��Ƃ�bGKE�q�Hp�=�Ah��-K� �vm�Z�,V�!"��W��3� ��z)<fN�+�g`w�T�n4�3�H�pqyN��Ze}���B���7��eT��P:�^&�����^Vox!PGt�FQ�R)ϑ�Nܡ��Y6�VvD�
���Cr�V���-ݑr�{�e6<�6�sR���ɵ���PϹi�o8�M�>i�(g{���fG:�!���^Jq�ݗؐ��f��P\�;7��*�z��U.N�t-���^Ȍ�mG����N0�L���L�v�s��l�<m�0����[����R	�h��MgC0$� C�b�%�`<�d��Oj�N��G�Г�Z�@�={Q���9%##䃣 ��Ec�r��*�YWu�e�w������Xh}0�>�}�+a?pA��ѭ=Ȧ+�q0J��ʍSQT�Zl��P-@���S�5����ِ�.�{	ڱ�
������;��y�Om�1�nC���V�Q�q�8?�5<�+�����]J��=����n$x��Xw�)�ҟW�K�Fsr�|��K��