��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����F��':�ޜ�2̼ߵ2D�c�k	�?��lK���ګ�6�6K���}^��xF�u��hkp;���j�n���WVܫ� ����c������jɭ�L�5}��>��<L�=l{��	�Q�D�\V�d�s�囏���Qz��
2W6�ol��hX�| �/������¾7�z)�5���KUo$��bv̛�EQ��e������Q,L��d�tӬ�7���Y��]7�9�MD�vD��g:����rz}�|��x2��8R��X}&}R���)XGn��l���LUK�3�s��,<NqǬ�l�ٿ8D���qd]_�#�c){\�-�э�dK��N1����y�~�.�ߘ�c�� �]ئ��(�����Fq���-���F�e*9������
B��1���}ͳ[��y�?�,c����}��O�sW�Ɛ�ö�i K�lĪ��&ެz����Ò��$hP�?e�=���D���>+�`9��_Vs����͎�/'��I����_���s��A6#�3���h�<��J����v�F�8�2�Y�h�vhm(&��N��c`i�#��+�4�6'�q��0���	�x �Y��c?�g,�?���^3��HŬ���������o���5������x]�9�[���q��)Qp`�R,�ʳi����}�����Yz��r��ʉ�#\��-���l����g�CF����g�uLx��f�K�jk��Xs�ǽR0��Ub����� ;*C�ٲ��^�0�X^&I0O�8�h�V��M~q��J��(����4M�
�Qa"��`H˦���)�vtť��1��t��ʭ�F]��-�ƴ@�k!�o�ܞZi"ٵh��P[ę���t<7��Z̵+Kmߦ1��%#����M/դk� wp�V�*�~ZF禞g�-71&7���:8�e��z�8^0/~"e�`F��fBE8:���d��_!}�/����ݽ@o�Su���GJ|>�����kԵ�.��e�c�V ���� ���JH�I��g�l�D�y��v6�h��}Г�����y|=�MZwO�{�wI��O#�.㴤?��L��k��Pxx�4����E�=T�Ӂ|f{4���:�ܱ�?"��E���<,��[�]���t�tN��l�J�:�q��%!xg�C/�ݯ��b�~�w����%텟�WIQ��)dB�3��H�{#�~�*���j?��H��y@|J��۟"�r�R� ��>�r��*~}u��*�$�K�o�؛"�u戂u%��8d��*	'�u�u��&��?���)�NZd�in6(�P�+RQ�KVm�rN�G��3�sj8����^�H�
W{}iR��
4aE�F_�������\�%'�q{g|�F^lI�Za��W)
���10/��OAm.D�HB�+��V:�������޾F�C�	�Pyn�f�m����9Y%�ELː1C
*�F�~�"�<_�vR�ј����~?1����3*;���M^F�£��x����h[�E�'zJ��(��	�
)�P��N.���^MHԸ�ƛp ?>�p�8Ѩ��
meVHi��2l����~Pg����;:�����|!K�=F���F���b�GZK���塨��4lo>+e7J�Rx����񎉤ߒ��:Tݺ���i���ݍyY� ��؀H��m��)���q�ԢV�?��`{��	��c1�Fz�.z4���-N�q��]�, �'y�~�M���v��-�L(ۑ]��"o�=l|��Σ�G�j�	��Mn�0Ƈ�?r���x�\�Ƚ-��J�*��]Hlu�I�}�[�U��:y�X�O�ں���&�=g�,�6��X*�P�gy��=��˔�E[��\i���I����wR�pèAW."v�y�ءR��C�-������3������,��#��Ğ�32�q0��E,ܠ�[ �/���K�ݳ���2 *uk�O�'���"b=��c���<S�;.n��"�,:�{@g��?�pK�y�P�my�[&��=\%Kd�i8[�:�-��v�8����[�����t ex�c����D�N���Mr#���@��NzI�w��J�  ���ҰlLCM��d���]S[ӽq�k�H����ܦ��y��`�z����j��3�ȭ;R��q��&\!J,B��X��k��|M����\t#��RN�\3�J�~AA����
�/�ňy�zɾ;8%#��0S+@x0nҴ��T^鷙�g��fVGd��"�O�8V���Ih�#f����+z 7������W������9K�*��U��;���.�b�|fv�++lr���CY�,GV�:~�pF����%߮LmX�[�[<VQ�:�&<3�F.�����!��W��Q� ��2\_H���r�2!�JNY)����T��T�IJ�����9��?�J��'?�G�# A���&�-u;(�a{=��V�<u���ELf������ϗ��T8w�J�����;.��q���b^mT^Q1��m�W5VlG�^˯�v�.��\#~Y�����&b? �dHY����`⯛`�>	I��88	f�.u�
�l`�d��n����s"�@�r�����h˻Ά/����	��YAI������2I�~�� �P���Q@9�҇��!K��@͏�%L��6�DNr�j+��+m�_$8r���v+Ewr	��?�Q�j�$&�ۨ�>X~��Y�TS�C�tO���\7{�2���E�$��)��6#a��&�l����cNLU;3�s�I���HD/��uG!��u���9h��1V��;�3!���
�?���o#98t�`�)�����9�r�ج�R�ꖛ���,Q+���w��.���(�"�vAK��a���H��϶�7�0B �7al��p"Y�m#�*M�Wc���}j�nD��e�7�U%ã\Z���� n��
��%��Ĭ�.��ئ�{0	D芎�b �KlׁE4w�e\�p��9@����ޫ�ZP&I�'�z�UQ��-��/u��m��O�}�p�-�6p��Jh�A�kk!����(�� �Ҟ��>�$�Wʟ
q�__��6Y9���4ʩ[���+������1�Y�Eϖ&� �~��Ճ)�)��qU�y��
�K٨AQ�F�{��rl[+H�5kڃ�3ť�Dv�ø�4'�@��fr	���}/�3�0>�?�Qx�.6�Ab�W��#F��m�5�%���!�=Ӧ	�z0���-��!��f]0��ѰI�`������[2���)�_*{�_����78w�=Yŋ���be��>�$��)��n�} A�Q{����f9��^-PBS95�Ț���xh����Z�#���K���T����pᙞ�	�J���$�-4��KEw �����kټ0���i�*-�/�K�;lh�u�WF��ghj���PM4�Sx�������69J�����B�m��ErsG�
��t���BA���"{Q�wW�SI��D��4��QP�4��)!B��|
���z#���u�r�U�A!VT���W�ݜ�fCP��o��*z�\�5򒑬f��E̫ 	�����yMz5��_�����&�-�ޓ�);.Z7���� �����%I�u[h�Nd��̀���խ���R���޴Q>�{n2�9�l4jeǒ m�p��)���K^�V.K�@d�X��`�N��Z��B�eM��㣪�GI���P؈͞y6b��c6]�t؉pum��c�2�U*x�e^�K�	��ӫ �P_ve���#zF���1�� >U��ZYEO�f~~�y �'j/����QʿP�"����=����r�������������M�˶��N����9�۪N3!�~�,$�:>"4�)~�'V�R>*�C �F���?�B��������=�~�=��Ur��n�w&�kQX�ە�/�w_o�/��4'q#0�Ш�0	/�2��M>�W:�������<y���|��׃�o�7w�Zˀ>�#�!� p�Y�lw��n*��4�ޡ�ג�e�������݆�ȽTۄ+�Ad��fK%PTW�	��.�Xs�h2P1o+��zω���r4����;��`�$5ؗ���cȊ�!��ͧ���DG���,Ӷ��h�J�o7�;�e�A@j��m���Y՟'a�N�@"��t�h 1?	�95��b�1V��$u�Z��/ղkÖ�:��Tޮ#������_h���L+��MG��Urٽ�N[���n|]����e7����@��X�R�TI���1}F��t����,��5ć�/��R�/�tm�^�m�)��h��i��_%Lpo���h����V��9�J(@�|h"A(�u�s{��F���~W_�E��6w�ܥR�,X�d�=*�e��Ak�e&zP@RR��|*��C?���9��Z��Bbc1_	9+��l#M�١��@#�ԣ$�f�ݿ-3���'�����j��0�c?�k�v�3,�΍�څ��ʹY�{X�z�x���K�x����>O��os��jُ��v�!Ƚ�pS�b4=R
��Y��W.�%1����p�����k\�a&�P��R�#��{9�Mr��b�DE�$���<�
�6F,��84�'`xGYC�m�>[)��s�J�����x~���"���q`^�8ou����6��xQF���ȭ�c�-kr��.!�dC��Hz#l��nMO�[��D�KL~�<��e���V�/�����ѽ �S[�\f�D�+�-�e���sʛ:P�5��T;�zT�3Ӌ80������ƺ�I�f:��Oj�7p
>�y��٬	\cd�����>}��־7��fՎՁ
a���V��!B*�wl;haI�M��p�6��Q���OUq��ڕ���Va���q��@���nDJO��03�:���Ѭ�����ܰd-܎�_]�,�Uz��%����6�@ʃ��`�
1�Ujv�d�$�s�h#�"��iUl���NݎK�a__e�y����\� #`�j�ei�
��?�Kb�IQ���ꯕ	ŭC#6����_��	�x����Y3��lɜO1����N�+Dたds�`wx��g��#�eW��ҟ�3Z>��k����4r��"SU��U�c�k`�Χd�|P��h�8��|$�:W�L2Vj:@�.�,rq�j
Y�	-�4鞘�LG4��Ս+��6��k�F6�w���Sșg P\@2���,s]��҃'���H:����#1o'�o�>�W���^-��?OB���P����;Ìon����R��	d%7��:z�D��~0�}����=f�"O�~=Y�\�ե�9����S_ΘV�w >  GF��C�βYbM��=�o�H[$52�(А��ֵ����G�?�G@�T�H2]Of�v��)�\�o�8��E�k�vS�w7u�zR@O�������M��IQw�H���HN��Eyx�plF��nd��4Du��/@5�~a���hH�%A�W!y�H�x��x�y��"�B���<F�aʼ�[�6�h�>�%~6x�	��w�xks���dk��]\��"�A������ydb�I��gVHEn���*�K)x���*h�M4�l�����Oj�D�KȲXpŴ�w^�$1���p�ucR�d�*�sigm�(ͩo+�ΆO}ޅ��,V����0��/�~ԵPMd�-7[䒷�B�y:�a�vn��n%���J��b�΅ �I���Ix�&P->�%w��w>��8������j����	Ǹ��p����ʫ
�"e�E/�m��3�����t�o{N�0Os��� �V�)~3�C:���l�<��UPE�+p�_� v��{�9䙒~	j�;����;@��`�7���Z&��̩�Q����ÿf�D�Ѻ���/>�رL�"BY�Q"���jCl�om�Y�bc+]��xt���tX3�5�p��#t��xҬZ�]n/m'��@����тz���v{o�������I�/�l3xjɸ?3wD�J��������K3\�F�-͋��o1Yw�R�Xl|i?E�h�ȶ��[cP�����Sp�P�X�1����_oDI��\�|f!�F��6�Vb�vO����%|�sh*���u�iiq\k�g� V|
Iu�2Υ�0�_��]T�̶*GZ��6� ���%�'o�1�~�`ڵ�V׶rrB�6n�7�Vڗ&��Ά��H՟V���&���QP	���C�E2�{!}"}��`���[�rΌ���
��b9W˵��}��4��,{�nn�r��L�oCr���%0� eU��b���� b�y��Lt��b��p���@��ҨS*���=y�����*n��ϔ��vIUl�C�;q�S���;�����&����D�ai��=�X	꼆Y�I��!��?�,�A������mzS��$m�şz�Bx��+'R2a���9�l�d�?����i�r�����O�AV�7��+�8���̫�.X��I����
=��	�He�;�����@� �w���/tvpS�Vo�_Ό�u�4$�Ѭ7g����{��L�׻�x�������!0�8���d��3��xO|�<��٠���y�뚼w.Q#*�� u�B��+(�J4vu��1�-I��h�igj�J��<�p�t�8[	�f6�+��8I���{M���eJ�"dq!���%)��ȺV������:�%�UB?�@%���)�.ќ"�|�ҕbP�}K1+&�u㩢��Z��`�S�"��I��:`,s�ڬ�Bd�Bѓ�|\�/S�hĉ�΅܁f�C�|��Ea�^a��z��}yˍ] rf�ˀ��Qy�H����W� �>`�׻妲kA�s-�sp�oq������;$p�H^��ni��`O��D%�7���t��=��6����`}�LM]��r'\[��ɺm��+_�|/C}j-'�:}_���T^�/��g;��东ez>�vzhj�lzuG��lv�X�^����Ĕ� f���Ĝ������0��]��4�d�n��PB�\Q��Ԟ��.db�����׭��|V���+O�4p�xh|O����V�D���ee)��*�B�o	v.,Th���:���W��kF��ʳv��C->}�v�gբF�������_+m�r��@F葪��3��t�k9jQiY�R�sbTs�Z/P�0ģrY���"����E�HR?n��A�Q �깹<vb�,��;�0���?�����S�y�ZP����?�/�:�Or�yd�M�p��S�@�f�|M�ќ��{��៬nM����锤i� /"cRI�T��a'5nY@��Δ�&�Mw~Mx��0]�� v��*L����tjG�T��dxq���6`vP���"�xp���:��O�; �.�뜳����.'�dV�:=L�F� Nu�NjT=�}`��)C�_w�%��L*�~������d@4s�µ�@�!��,ch���hK���Eꘉ���ܯ��i�bw1�ٹ��+Ȱ�ǍAh�r���.���b\)�=�6�k*q������O�g@�w�m��T���GZ�0�S?3����E\��p[��y��H L��g��5!�5���6�� ��w.�	g{�o��@$��[,!F��瞹`mDs6M(rp��q�	HQGO�J�<� ���L���~G@�|�ͪV��0j�؋��� 9x	�N���f����v�4"T����&3x��0׹t�����~N���뛾�����9��Yz��3HPG�BX�_v��'d5�NYe�.=ZZ����j'��C{wG��5߽Y�2~|kV���lpm:�������ײ��݌�03U���6�R��ì�l�ߗvs`�<�����G�՚����h.'*�-J���[���Ґe��IL�C-$]/	���.`��d#�GQ:�=�;7:����j�Z�6=�����ba��^VO��U���S��$[��V��6�@�h��Z��-�y��Pm�x_��Iہ�^�m�����	/`���K��
�
��%Ύ���>�E=tx��R�z��ͬ���'h�o���=�d��//�SBzܴ���I��U�꣍2}����S��YyZ�S�_�<{"^���ϋ��q���Ǝ�8�#������maz����=�"��Ԏ��<E��3E��N�
������티Hmҿ�e��.��4	@̺.���8ڗF��ŧISs0�uґq^�.#��z���<��I/\"t
1�O'�1@N3��'���G���%��`;a����}�#/xJE�V�Y7F�>�m��N'��{lь��A*M0�صEB�Ҙ�>��ž�U��:z���V�}gYI��2�����N�a�T1/�:���
HT�c�=�?�Y��5��{�h�lp�8�Ð"#y�ݣ��\'ΰ��I�to"z��5�д�i���9���:B1$U*	�k����c{ P$��浟*J]��r)�w
V�T�4דu�}�{�-CX<LNM��!Ŧ�7�x�>O
�\��b�t@�.`��\�zC߃�wj"I5ͬ�����:��2HUT�^�,�O�*�ܚ!sN.�}̹�X���]����}mJ@x(i�0j�s$u;��-�т�JP�����zc��9���V�wd�fst�{NgpA�S0!/:ŷ9�h
�b$jK
��0ؓI�lXѐ1.�_�B�J�j���GĢ"���&y?ۓL%� ��_�e��P(m�t�\H�AS�$e
�9<��=A4�ˎ�LW�ǍJ݊�Gb�5�H��]����y��q�gB
J��G�v|�1�F����7pyhj2�ۍ�7�y�>RF�6@�t`�I�?W'W�f4Ѳҙ_x;T��'0А�&��J��=�q,�;26�f����As�k��/j��n���4Щ�Dj*5y7�X��l���W��%Ox'�[`%��f�V��p�[+\l�0(���f��`�i?�ڝ��N�Cq;L��1=��u�p�Q2뛰_
����-�Ƚ� �Ԡ8?6���M��׷�o��4�?��ᙘE�s��m�m�8J�)=��cS v/h1?�|WfQcr��1�$`��a�A��i���_"7�x�O^"x�1'b���w%~��2�] �ޜ�eH��޳�|�?��Q�g��[C�gW���u�|��@xe�"�wߗ#�Cc4`j���i����Od�a���b`"����N���P��;�vX�`G��1e�W�6I���}#�����
��A�+�'J���|���;1��*v��ྑ\w	ۉ��Z2H�Ee���0T�����f��R�HH���hH�zr	7��������V4|d�%�"��zz=��:�d

�萅���b(0������M$�M3�p!�����#sF'��n{l���<�V��4n4Ԃ�Z����ڦ�����˱�~J'�b'~�	�Ÿ*R$�L���h��v���b^�K/|��O�%3�@)��U��,�������KԻ ��m� Hpb5��$���o$�|�̧�F��:��-��*�!?.P�'Q!�nN�`�ȏqѰY���(��j��b��������р#�L�u���<�\?煕@餾�r���L�޺�{Jd��aDŋ� �pՍ9������&)g������ �)�	���4V�k���onQR��� �MY-;b�m��d�dT�b����,nw��*�ـտ:�'s%�O����
z/	JK���	����N~��m�yC�me�+�\�?7b��zW��4�x���F��"�A�d�c2N�q~��X�e71� �tP��n+)�ʋ�([J�� ���R�5�<��&W0����\���5�8oB <��������vq�Ƹ��m��w�d�|CD#*_��jRM�wD�?���fVG� c*ğ�b"D7��=���[�Uf��a�R�-����ψ�j�u�;Y�i�]��@hk&��]��H�  ���26z��0����G���?���^M
ߓ��N%�M�ês�쭜��$�f����ùS��5�W`�Ws�����F;"�>���a��Xa _l2�׮���~���Qd,�a�A�X>l��\ �oc�f�mg�ٷ��b�	`���� ���a���bz��鎰����?�Q��*�W�&knZ��x�k������=�C��|�o��i��|�*/��i����tC�o�ug��k�9�$G��K�\�x��!����_�=��T����;�-n�ћt��1�(odR��*�ܺ�E�z:%�)��Z������َ(>�@K���Z�'�G������ǫ6��o��*Pnr=�Z�H�c?{����/�l��98!>���-�{�Pb�)ej�9�  ��	���m�Q�^m��R����Κ��O�8э*���c�NP<EϏ�udi�ʅ�7�v����V�k�ΊSN�U����i_�˸GU@t���<-"�$���?���{7�����6�"�;���økGkF"�y$Ê�%DX,����B� K��Ii�*��M�lJ�T��
�i��!�B���$���ԡ�T1�&e�E���p�G$������ŗ�
*b�E[0l�