��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We����S��$tF���e�}�Ꮇ
	����ÀǙ��<�f�Vģp3�&�O��E^6����
� ���%ap�W�֘��Ib:�������ф�h"���I	�JD]�K�A�/�#���K}񃒂�Ib���v��'c�s8�����vվ�9�Z���ݦ�=�8��A���8*�]��ϳ���N�#4_=�Udg�bIp��BS�u�<���.��G�]�xc����d�e��ʞq*Ee���)0�C֗.�R�����%��@�B�i?� �����~�h���S�sW��s-�0|�����͘v�\0����P�S]�cR���O�=��l|���b�0h��@����F/=w����E�ȣ��1Wz���t��N�Et��`8�O�����[%RC7�^`I�Q��t2��v���[毁� ����Mˀ2*�*�C�f0	suМz��d\��vʵ]��Q�Z�Sԣ
9$ad�@R�������t��X��o�����,�����dcב����D��|��p��������5����u��p��C��/�U	�x�����'(�oֆůuާ5	�R�eQ��%��4'�3u�R�J2�E{��c����L���j��J�- ��_�௃��^�i�W��L��Hڳ�Kc��^Ee�,Sy���[Э?��.灍���TI`]	L��ց5S!�e'�@��(<�a�Sl�pH'-Mc�asi��V���Qnm�v������?w�q=o��T=�d��@=$��8�2���ۃ����~�y\t�G�	�$Xx�w������.B� v4� ���d8M�+Tedf�o{g����CeXO�B�V5�q�
CX��*
)���e��q@!X�(e�:;!Fr
vM�������~>�?nj��-sB�(��A�XV䭔��V�nlwjA�&P ����~�ȟ�P������2/i�]Y��O#T'�/
+5H9�?6Y���nƿ�$��z�@
�Wo����ђ>��:AL��b�����+�Ŵ���p���F,R�.`��n�s	�	�Έ�m	��R��C1~p7K��qXB��4��~2
��i�SW��XMYTB&�zxj-4��9����/��IgE��X�8���������K��q����~�ہ��O������}O����Ӏ�tDB!,�=xm�G/��	����w����h�*;*��i���SW�4nQ�ҫ�|�?��o¼�gy�-�1�kJy!�H�Ġ��_�� %G4�2n�Yw�)�oD_����)�._�Puc��4b"�V]���Oz��$����k��n2���*�Ro\��dy��7,��/�DkBȅ�&Y3�ʩw��V��iЪ���jy3Ҝ�-�JB�O&y�c�^�g�f��c2
��^��qc���ZL�K���O:��]�vS/�%3e�$����킁]��\x�u�1}衚�Q+��Lh|*�ɚYw����m���]���!��Ie��x�6��o7�V��o��\��nZ�8�12 � ��k �{)4�_��-6	!|�����sժX�¢�I�cJ
 |��i���I�Y5�����_ESOK�"�d9��A�OГ�/s/D`�)�Q�)�%�͔}��;.�5��	eUZK�z��ላ��MH��v�KmX�����SiV�f{����Jc��b�&ˌ���ɷ	g�Vg�~>�iQB��_-��NiTIh�X���W� ��/	����Ւx!�X�_/x���-�Jp_aQ�~�\�HbT�X(e���8oLAgf���qYg5'3����I�Y�Z�T�i���������Bڊe�xT��	���Nx�Y�����x�K�$����+~B%_��V� ?lRrB�I��y>Eɸ̦�r�_����Ǯ���ٻ%tt���������D��ؚ�Fመ���5���[��j1����կ5�h�<���G*�$?���=J�!s~���������>�|��M��j�+
�.qڑ:�/�>�I���+��"��Ԑ
TbU20*^��8!!%$�	i�t\��,笠M��o�Z��ռ����h$M22";�8q$�(�L�e���6�/�ҡ����(׶�R��Y8�%1��o�!�A� Xš+Mqol���K�T]��JĠ3�_�@v�-���Ч��u��ғ���!��Z񜲺���7P���P�G���%����l���B����2�jJ�v˙���6]c�ٚU*̪��x��k?����"���W�eB	������`��%�_Lc��	G��hUc�0��^�h�%h&�`Xg)�@�S�%�_�MIآ<��el6�l�V��B%���=d�R^�G�q���o�ݚoJT{U�{��y�]7uh��*�%(�����!P�%(���0;�S�q��>QR�!���R��׃3��
4��3��R�.֛O9�t*=O퇹>Ä�d�p���W,<@����z�eD�����uYf�/:�3S�t�z1�vk2����7�K����$�-;H���V����eнy�9lgn�ob���O��b�5mk�k'����7�m�L���&���Eft���.F׃�� %3w����~��;�;p�6f�"���g	
��%#n���xyWi�n��N����`-�E�K9�#�25��Y������ѧx�F�MI;�KڿM!���/���;�Z��z�� h��O��@]＝	�F�Y�i�N��N��͐�7�}��O���h�>�����~�Q��Ď���tV���W��~P!I���M�
��o7M+��;iT��/=��w�Ͼ�~'�b����D��o�C��s|9��vf+�=_g�jk��v��U��#���,s�8�vAh�~6h֮#k7���\��;_Чg)Շ�$�Uǳ,�<�ԇ�J�7�oF.F�+�%�(&P�o]IfOM@���TM�����
S�W}����d��7^��
���F�����>Ϣ�prh�.m�ճ�5��{�um[�&<�Γ�c{(�~��7��7 ���Ng����aML{��s�()Q-���Z��:e�<k"�)�ٺN���
���$�a��[d皺q'{6RC	��m.���Kih�LɅu>�|f��&�Y��ұ�6޺e�A*B��<]%�:-QzH%@�[��+���3t�ҩ�����>L�L��-�*"?��{=G@3������g}�����k�@5_R��GMI�"<*��
'�N�M#�
�.㇋��z�Ν�����B�tTK���Z��ն�h�_�=K���yz1�=L;�Ի�!*c�M$�&�r4�L�b��F��dPR����p�҆��0j�Zzw���Y�]�|3�7 ���,Q�Щ��G}���v�P��Х<��}�����e�#d�羚�y��yǲ���m��c'r8�?)��ܩ�EEiS���5���0Q@��Sa��0rk�`�4���3)���>xR�ţL���nc�摽��+w���f�-�}������C����[-f�;I���`��j�S����;����hr�5ӿk��E��tf��Ij-��E3���/��Phz���R�|ĵj�!W�z��:�s�	�/�
z���*1O��H[5#��d��QN�|���±{{*��Fׁ�]��z�����_hJtJN�>L�� R���V�����o&���<o��k��z�i^ܒL��0w̵�����[z�8�p'������J��(�%O��5+�$�d�YA�D>��
y�~�Y��'7rEW��k��6�N��m��Q��Z- 1M>e��1	l����D��$�ު�b�S���)�$�M�6h�*�^�׾#H��*>p�g�<���_q5�Y
S��m�0��>M�9"���|��Zs$���V0ă�He�"m���pS���߮>a��4�7\TQ=�K��R��1S�_�	��KV=nەY�eA�%FٙI���.�Cٞsf��%�8x��?�צ��7��͍D�����1mҷ�[#�v���u�y�����qȊ*�1���9_�N���b6�*�yW��^8�̰�$_�]��:�	!t`�����U��;����#�6t;�T�jJ�Tb��}1Ng叏���@��k%�{dy��R��3
�H��v��p�e�V������4�9�f�P�)���S�A�lA�=PT<}�Lr�c\�̕#�����Il+/%��l�<j��Ԍ�ߘ��R��~�~S��6z`�5�y�Ȕ���Iz�Lde�2(i�۬'��w�,�q�HW�[�丩;2
�1���vx��hJ[������z���O�p��LW�Mw��uk ]|�HFDB�ҵ(]���Ĳ�$�nZ��s��i�VF�
s@�Fa(?�C���%b�"p�6+�>ǹ���O=h�3��ɬK�A����W�m���ǣ���<����4p�dm�Z�3
���n/}s{�e�Y�P�i`\����,
�y��< �:E��K	�v�ֈ��ߑ'�����Ǹ�F��^��Y�g�'�|�i��U�eg�D%�n�!6"�<�������<�����K���FQX"يl��f[~!.>o�
��Sc3� ��j�~�%l�Z�PJR��x��+Q�)���0h�҈��A�}�W�8���g0e>7���eGM�0��J�-Xm���mFf�
&��p+��� R<�)�Z�ʐ7r�o�}��X�
�	r�$6-WW��ڠI��IP� ���{ �-a�c����9XV���I>	&�	�tp�!�������I����^mF��J�rn�?02N�L�[V�\X�HL�ۤ�\j?}_X��'� }<�+�X?Q�	<�8DEcߡR��_���"�昔6�T�e;���@Ǯ��зU&��a=�{����w�B�>�*e��1/��eg䳬'T2;�Y����Q[4�~2��rw�E�r&��p�m9�S� 1B=�33�-�_~cV�!�2�M��Fih���o��Z�=�t^�X$��z|~6��ū�
Yl�	o��JF������ko�1/���c[�eKL�+L_�Q�0�4����m�f}���_
LE�B��b�ۋ;�p6Ȏ���L|��,�V�����t:{-�U�H�W�N�J1E0�S�q|�vxd��W%��s���u��E=�>B
�_���)�^׆3�� ��<�N�NRȸ�4���A%�g���!�o0L+�]k��e�)}N���!���r�hO�n����K�7I"g��Yf�v�.�6d���C�S'�_��e�'T�!"��x�4�C���3s���6 HU���x�i&��,(�9F�)-��fs�?��_hO�ݖ~ߊ������|�ۈ�7�)��Rqt�R�g;B�����i�j���K����{|k^h�!��-�Ȗ&�3٠z8b\u�+�j��:��c�L���@؎����=>z�,G�R��S�$E�[�a{Z�Z��+����؃u�sbj�����WtO�\f?�����P�'5LvP��Ba�_b�����F1����'�1�0e���웖��M���E�5�2�[}�*_����+�?!M�ᡴ5�&�GGBG�ƨ�/���=-w��U3dk; ���@�xw$
���_*
�	j���&'�&�7��~8"L�'�_��HI{�2��Md3#�o���TgCQ��4��uwƴh���K"��碲9ó/
����KR�ԛ`���&�5�LȔ�	+��QQ{WC��K�>�s\!E��9��;a����F[�@����\��$�"^)�v���q���]y\�	�f�<4؎�����%�5Q�޸����%IQub��`(�'����-���,�6R-�wk#��e����K�F}�^���]f��σ+c�uez@^[PX1����|��0������]w�7Y��+D=5Ŏ�tIˇ#�h{Q�ȫ\*Ϯ�~ZsI>��^R��˂VHPK���T|ךϵH�}>��ʁ�a�pD�f�]���2�Qy��O�Դ����>'Uմ��&4���)�>Gt^�Tm
԰�Z�]��^3y����f��3��bz���+w6!dD]�{Uۆo���)s�'g��!e9�%���=����_���E�r&d�#��8�5�>'����3)M�vf8��`�Ȥ�DP���#Q�u�՟��sr�Y݉o�ֈ6��1����v����Z�X!r��Eo����7+�sԅ3n�	7˘e��!�$<T��<}V/�W�U��|D
��b�XU���� �"���au�����҂e%�«�ƀ�>���DO"�ѥ���؁!�E�`�q;�XI��nO����0�ru4r 4Og�^�Ћ�;H�%��,�ɣ�jAe㶪.`bid~�?��Ǝ�Be�\3�@���+�2����J0i�(��oG�S�r52��0��Kf#G���^�
w$&˥�KU�6b?M��3�#z�~ �k��F�Z�ʜ/�~a��i���O��3��[m��7��7���A��[����d��%��V��_Sʒ�p{^�7L�D����d[D�6��_18�A�P��.���c\�~�A���p�8@����Jܺw��T�wݙD��K��d8E����J��v�h~Ψ6�􅢐Wё.��S��tTD4[>�� G�}&��*U�צ%w�r�?H��y��DW��:�sx?9ǧ��L�V��x`���M ,p6P2"��K>J��$���ƛ]��(���r`l�
�[(�mrK ���[�?�5����������F� oAg�BF�.���j�5m������%����f����x�}���OQ"���|�#���ig��@�	3#R^��/DZ}x���CX��W\��~�p�r�P;��'�%nu( ��ALC�z��@C�`�U��«Ί�ð�D|�B��?ky����lX���� '3��(�:�m��Ng4b�wb���O>�#L�a����g��%��:�b3���3���g6����k'��:���V�0;��Mg;���P�yJ�M���������ҏ���6�Zg*e?<�y��\���Y�;�j�����V5z�D��x�G����%H d[+9/�Vj�ٙyM��D�C>��{,K.nY�!,!O���kF2����*-��?��jS,���{A� 9Q�2����E+'���XQ^��w�L��U��m��u���S��$�f��,Qv�/%T[�\���On����y�Z�c]}7Y�5�8c��F����9>��}K�0r���6�jR�2�H'\����������d�5�7��vƩb�U�j+��[3e�7&�~���g����s���r�j,�E����p��d��;Gbz[g�Oƃ7D>6��^�L�W
���q��u�<0�T��_?�
��؇R]�T�7`�G�3�RQ▛+퐶o��1�28dm����73y6ɫ�0�phM�r&���ݩ`0.��\�pS �����t�GZ�u')���h;i�8��"\�xV�`e�/��'b##�HlV�8�\1���c��Pf�zy��8-fW�B
z���\�2y��(�3D>s�q�<�7�uYKe�h�X'��ĝ5�<��L�QW��>p�8�>Kf�䊙�ҩT��(�-���>�Ho<a좕�6y'����e�uW#�>3�'/:d�%��B�9��k����ODk'k����4�	¬ >�&��$�����7m_%1&�9�߲$���q.L��c�4f4O�l��J4Gm��~l`���^�ɻ�-8�B��㠊��>4��t.���5 v�Y��%��P@W��$���Ƨ��C��?pN�Y|�B)=���v��gc�Y8g7"}�b������z����R�4̵�M�xo��ƴ܀��S�w���.g���-�'}�=\qA��
e,��K��x#5E��@.A�5�=!$\L�_%�K[�|�:�^C��ð�KYUj����a�%C��<m�-��<|����BG�F�7��Zv�`Բr�b��R{��P#RUl�Z���qW?}C�*R���31��-�LT���W ��H�Š���[U��1���i�������3�^#_���j�q�fgi�;�F��0O�ɮ��R�U��?���e���&�r2�4a�Y�w��0ʘ�~*4�F��;�/�԰��4(�΋��&=����M�ԙ��#(�.|)/�Y�5-�N�}I�^�"@w�ע&�њ�J��d���>��X�w.�i* {zJ`�nkj��V27S�B�N��)��������H����%�������m`
��Efε"0��=��$��q%��Hs��YؕW$G[]�U�!ed��֓�����q�\��&��k��@�O�D8����>�Dˁ�1�83ɒ9��-F�ӥ	�]1?C�=����������wƏ�|H��yۯ>%�&V5���#�`�V�ō�s����^��(6b�4�1�����\����d��őT�	���a�n<kE���g�Lr��ǹ�h�A$l}�I�0�B��C��-ޘ�G���7.��W	�>R�J��1 o�Tdh-���ÇO,�xͶ����������n���G���~	��EI,����Jt�KV7wk����c@jnB��ZHn�Yŏe�/�v��z�-�`ʰ2.�zo�n���bU��DB.�<�WT�6&.����Gr��^0��a����̼�>��	��Z���Dd�/O�ROk�JÕ5��*�2�₉��6�a�?s�r��G�pg���፦�W���b���c����Ȁu���F@&W7R��tJr����t��V�_(Ԍy�� �('���8��p�y��'�6��ӵ�:gb�����'��WE��8z�t�����l,������3y[��%�{�d+��P!�������ڬ�U��k �Β�=���\ʜ��*�_\v��Ћ�>}������r�0>f�-���h���[O� y��,d�5a���!m�����\ҚL����mA#vFtB/VE�%�]1R_��/XY��8�l����v.j���[2��[?��c�ߖ����m�mV�����!n��h��މP��$�i��Q��cqC�Hkլ1��_O�dMͧbP�\��H�LY�2�f���U��wvb]�
�s�x)
���=�ۆ��oXGp���bE>�h���Ŀ�<,��b�
gE=T _�eS��>���2}'g-Q+r��{t��Ւ����.�v<{y�"������b[�	���qTv�\��̃]?#.6�_f���܃��&Z�����4T3�Ú�/#Ѿ�PL�FF^��Y�}=�Z��-)g�,]噌�:��0T��Qu$m!�;�$�>����Yq���1'��f-���I�����z��xi׆]�+4C+�,>q>���������f�k���I�ۋYbD����$��Ǌ*�V$	j^4�כ��$�o��{%/��x{����h��8뚊h� �J^]������PM	�؁g*��ɍ3�AȘ#�N�;_tc��s3�OO�x�J���nﱴ�|�ˊ� �LjV@�� '�,��^�� ۖ�����Ay3�>�n���渹1��+���`A�߉�O9J�+r���Uq,<�̟껥�3*���z��7�hn��t5}�H�F�! 3����S�������r�H��J�4���A�����iԤ}��E�\���l|���ׯ8_�8g$���c]���!�cK��nѢ��T��G���!fr��i/�d`d�Az������Ky�4� 5f�W�=��M��7��Ӣ�n��*g�r����K�i�$bO��ء�w!	�CMʹ��k)�6܅&)
e����T�jr�AXi���ĵ��v���C��ѱ��p������@�c�`�~���,?�g�=$Ƒ���IV�[kͅ��ѝ�W��>�*��}|+��7���t��`B[ ��%A	���bP���%Eb�|N+\�>�=}��*���'X&w�1x�[ ��R��H���(��S�����T,��iC�k��6��-�仾���|6�Bƻ��Q�8T��Br�.~�QI��'��qEJ\%&����m�j������^�uc�����N�3�ڧ�./�%o$�����q��e�ν�h�"��;p����^>@ˠf�%p��>)`TVغN�|ɓƕ���$rR��h�==c*^���'.ʄ+%���׶o5J�˸8������{`��Q�1v͢e�pj	�,,�l�ɱ��ʤ���<74����RW��xB�}����p���Y2Ţ�#�
��Z@O�mȠ4ș�)��h/ϟv`?^v�H<������qY��f����,�r�K����#f�jv|�}�S{�UjuF�,P�zb0��Y�O�
��s;�Y}x�����S�M ܽsud,�.�f���Z�3����A�O@[�������b_������E=b����\�
F���Zy�I�tc���l*&[Q���%�!~q`��Y�����G� G�9�RDT�8�*#�c�8<������G,�u��@��Z��}�����<�P7g�y���&y��߭e�g
�	v$&�� ��pU��nQq$��R�v�w�F�����P��u�V��@Ɉ|)�cE~%G�"��FI@m��J�Tɛi��l}�F+����: �lƲ�䯣�����{KV��bYB�Ϋ >�su���&H��t�eVV&�-2�9QvL3���$M=,������|�(�c�\G"Ѕf,뙮�:�oZӱ;Yiȼ��������?Z�i�S�v��M��a���sׅM?��$���&��×�ym�斤a�I���t���"�!���0�s�Tǲ��8.2�Eg-�z'�v@&�U%�����|T���"9����ޝ2�Ro��V���phl��v���U�G|��3Z���5g��*�f�`۔=��zq�&f����^p����W���qp�W���yv ;+JF�Dk�]�W�nn�s���HN*���c�R�䁪t�]��ɢ�L*�3��b�P�VJ��pl��M5O��+��<�V����w�k)��<U��KL�_��$M��q�q��0Ɓ����V�u�$Vt