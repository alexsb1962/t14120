��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�������ܣB��p�A/�=�S5@
�X�_�3!h�+�.A����G�{�@�L�{^8k��XD�"���]��~=����l��k��)�>2�2���������X���9�R���ݘ=K��Q��>�z��FM��W>��X�(4r������cl�H�_'�O�ַx����i��,��*��2��
)6�)hj��|nJ�ĄAAvFm'�=䂗9f�qC�N�gRbH��,�$J�~� 5GmZ��ڦ��^���Z�Ė�v������^�:�<�"�I�3��ЦF����>��8:�r���ϲj�tG�F^:��ыI,Ә����[�%U����U���$K���$�l���2�6��Cs�UwLZ�����9����?��7P�'<^:皇�^-�ۯA_��Yŭ%�k�� UYCB XzKj�mZ���~$���k@��W�*��=�#E�5�dY�OB��M�{��o��l&#���ay����1��Z�#��_p������XUɰ��Pm��
�zJV�`1c��FX�#P��j��s�g��v�N���B�R���t�PU٪�"�cm�0,vլ&�
�7!��_HB�/�7|��W: ���cλ��H�d=���Q�
�&������v_C�z1A�Y�!�z
d�n�rw�݋����Rk�b��bL��Hk.^P2a0Jr�w���>V�=J	](E���O�x���T:lU&l�e�T�QT�.�G_�Ĉ1���G��q'��J�5v�n��;��99.w/�x1b�|f�����Cڃ]�`�Gu�\x8V5cs�	��u���c��������+��e�w]H_#o�A2����g��:�"��٦v��%�]}<�BN��^؊���D�º����8��K���&:
����MILc��`���vx�伴n����]�ޭC� �D��m1|Ӳ�ge$rn�T�:�F!������-I�Y��<��  $j��sb�)X���})�E)c��䎄�|g �N�9Z0�VcV�^��|�T
�N����J N�/�fz�+�j��f���h�EY�K�^:^�h8Kc��j��^�'˂�h�{Ə� ��xfa�G���jZ��NX\ܙ��F"r�k]���r���V��Θ�1��8�Q�Po��6�¿7�ʎ�|�G���pI뢢��T�(��ۃHQ�W���?��Dp�72����=מG˭�8�Y��g:s7{���@����[�$�8w��=uဥ� ��	���e�3�(?�⟐]k�I�,�E5t�r�����i��'ô9,�*-�!}�CA�u�"�Dn5��E�Ʈ���>�s��ބ�v�=ݷveZ�OY9��IRbh�Ri�8%OZ��b��tc�m�!'p���Ұ�n��J�x*���E���Fέ�X<�!��#�����v(�@��`̚�e���V@��r��!ȟEr��5��k�y��X�u��h1��ڥ)C ��5���4,N�Bv��;�K�oG~c�8o	��#>���z�V�}%((�#�m��a��ȳ��M��!��#���8�c���3���$�#�Ю.�Q����&JwHh�l��i��b���������V�~����y.�1��ߘX?��}l�Α�����d�1�z�t��R�~�e/��`\2!��!��ࣺ��ˮF�+nct�i�:{���8�_�^&��|�!iϳ��]�k�Z)�mfMHy�1t3�=�\��Uq��֝�[E��O�z���w��Ү��q�MK�d��ϼ��|�)#eђ}�/b�mO���٬_�\13��+���l� �`q6sfK� {�I��wUB�K�������&�k�X�'��r��Ō�n�!��$-c��YM��GQc`�{�0�"H����*o�A0��g�V��W����]�@�G��V�ݰ�6�Y���:Y���\�>�y�YyV'���+���b�@j�iw�S��ҥj͂v�X|#�/x-�`���(5�$��i$,"4��@�M�$!���s�`Zeͪ�@���	%�S�YL�Q��T�}t9��'��G�!���ꐎ.�~ ��!�We%|�Q���)&p�����i�j	�&�g����4ҭ��ql��Rž�p�+s]�A˿'��RQ'����M��%�o먅��P˟��a�ms�ތ�,������L�.��_�� ���^Ā��.�{sN��Kh�i� `�J\t*�{L�pu�a{M�[�>�G�$�B�J�`� :%��el'�);U��+fqv!�i��j�����~�~��n��KGx]j-�#@Z�$��Ѕ}n��֤\��7�ø���"s�d����iL<�ʟ$��LA�Eh�ذ���Ø$���`U�7�r�C�rG�?�N��'j5�x�¥�d;b����t��4�Xomu`H�W��Ѡ�=�.>�&�V؏,�CM��IS~)s\��HAH�����r?ܷǜ1�x�G�yj�-k8O��2��J5�i����o}��/B�y��Ն�Ew����(&�Qvx����^��A�ꄕ�g�?��l�@Ϊa�/�J�&�C.R�����ς�;9^�������啬�r�"����̺��\����Q=��[����3J�aix�ԓ���9w"��t3	��sI�.x�mv��3<���|����D��#�
�~�Z���`ph�DS�9�+*��� ���:����=�ï�����m�-����RłG���ybuX��q~q���*�ҴÑBt΃C�YT7���kc!w�x_�(i�Tl��+L��oCp{+�Q֣d �� ��Ƥ�����ې�)��ii3�}<{JH(��?�ЂR���ąբ=�4��x�ᕔ�h���)�������E���{��iaq��M�.�b��t�l�˞q�Y�s�
d��R,��[9F���RCb�E��̉We����#R8%0�T�nU��H��n�۪�L=LKd]������p��b�_d�IF�
-y�2^�jkM�:i�����M�@�lOխ8��L��'Eb��d��nRfacڪHX�(�n�e p�X�o$$�3ލT�P��>� Y&�a�C�4��c�midk�M��T�ݛ~5l���J9XF	�a�T��]�S<a�q�����̇_ �8�Iy�q�K������U�]!f��"���(�k��U�&Ga_�gJ��� ��ǠP7@Uv ����/���\��U�#�o�fb�g%do7��20��+ד�C��C�D}�9�K��2R����+��o*߂:�cK�jn✅A��| $P��醉"m��RX���l%�ʺ��B�� ��ٺ;�0�9����62� 4��!YU@U>@�j����,������o�Tzm�{��\�j�Ș(���$8.@~�>���#|$�8!�4�I��N�ZX��ma��{�SSR8�4��&��e7�5�-��=\�/^07���M:xx����)��b��W]A��u܇^1�,��A�����iwn�I��5�'2��o��?R%�QYP;Ȭ`�gF������ �f�$�Dm'��yػ�@ḱ>�oX����s�a����솇�֪8"��FC���` z�4O�l�zz��>���X'��gC&y���tވ�%�v*o�.[�prp��}*���_H`HCҩ�i�N��R�&u�8R�u���g����v�m1����
��F����p9u��Щ|;��B�q�fv�8*�Xl�S�&]�<7�q��[��2J�-�R�O��aW\c,��V9�h�eK��Yw��%� ��&�m�/E�S�cW�x�D�$q�ˠ�Χ�'�C�24�>l�U��r2q�<[W���g�*z�6��D�u/,�ۙ�7��Fo�N~-O���y*��4=PB��B
g���K���Ȳr���\v,N������^�����}��r�[n,V����Wq�*>�I�h�Sz_��&¼O�ϐ���T@�㪌��Б��
y�rBE�d2��ϢĮ��2�&|�T]pG���qϝQ�F��@�H�C"t "G���VJ&[��R_A�;�-w|���V�a�c=�<����~?��Z�D�x��iT��bNS�'�?X>����m�Dq�3P���D�AR��L��!}窭�[��q���]"����#bYھ:렣�����|䕣z���k#W�c4+|ق�rq�B��uS�T�bd]��k��"8��Xzj��[C�����ƾ%