��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����aКJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå=�*����������~���A�#ea^�����߰f���%�w����Y�B�e���5r��/��΀O|1�t��$,�K��=�xx���S�n!|�{ o���#��o�(ů!P�Ōo�T�Z�mh���XĊ*`�����-H�T�=&&@-�6�8.�6xyv!���"�\��^��P��~�&�b������.,V����W��b�J+Y�\4M�x\s3�枫Ԥ/;'F_p���:vE)o�t��6�	�
_��,9����Gh`�z����T��u����mR��׀;>����p*�%�$ucC)	�ӏ�������8aQy!]8V�h;a�w�������Q�F��vǥ/�zy��p���ɝ�^E)����̵�s]M�L���XY����%�AZ�%h:��Z�e���(�h������#�pЧ����A[^�ub_��]����`�ड़�O����QM@�����d�e�'����9!*[�=���1�Bc��34#�T8����f#k���$xp��Z[J�Á��C;CU6�Q60���ۥ�����bzL��(�Qy�5k�ǵ��0��\Y����X���pY�:Wo_W_�wv]�D}jF/���9� ��^���V���ll��I�ЂA���\��;9�Jj"��^�� �e��X%^`�SZ����j�v<�E���Db�Vӥm�N�J#��C��'��o�3�ٮ����n-���c��>
��̪O��w�J>O�ɕ��{qNĄ�Z�3#h��G	�{M�QT(�t�Ǭ!ȝY��>W�@�5Q5���(Y���?`���)w��3v\k�7����=�[�PI���������mz0Ì�����Lև�L�m='Z�����&�Ba�ɋ�ǖs�������5�W���Y^�# �c-h�eg�j�U�6.�9��|g��(����"����(ɓ���*˵6x��)�?gĬ�!^�2��G�M+�Z�ڹP=u���Qı'ċ
N9+^O����V	6����Z�4����;��% �y����V��e Ӭ�i	����""N��3�Ld��A�I��`Q�F����Exf���}�C�p����ܧ�����}�n8W��]4��a��vݑ>?s����E(��/Io�ҳ,����V�F�S\�����6ZM��ם����Y���z1oN���u�cL��E}�����A��p��?��|1��!���>��x(j9&$�o���)�;�R�00���E����N)��4͏{���a���)�(��J�L��p>u$ _�] ]-�w`�Ct��Y-�ٞl��o{�����+�6 �:Ё�Z�ϰN�3���7X�b��V�z~��aìrc�	����CC���I=�*/hLؤ�O| �(4�,I`}TTkݎ���k
mȾO�;ln��r:C`Z�qV\�����4��`�"���=��7��P�Y&u=^�7H�a8�U2}�6��	;�K<�~�� ֲ�P\w�l�\�Gӿn�*�*RmR�Z-2K��i���nd��X�2�'�l�� c��`�k�u�6J�*
��by�ƹa���h
�Z�8�7�vљ�b�����J�7X�����|�"�߃�28�=mw-�B��?��>+�ka�`{�誖o�}�����f���J0 3�}���ͱI��dF7��ߓ�G}���"�ilo����-��� �����m<GE:Η����.����8M�xs��k������P�(rW(*���]x��%���ͱ�\q1��>��`�k����8:k`1����E��D8�Ї�����y���Z�&������� S��U�0�o�?��L��߹$������:��ˑ?�Px� �Ҍ"���[ �1�J�ށ�4�-����P�߃�����?߽﷛P� �rc�~H 6��UQ��a��E���r�b�	 �
N7�~X�����w�֡Q�)q�%s�E��8C�xE�kzL��Z���9 j��<����O�!�)щ�S�$�������;I�PPm�T� ���j�q<tƬ58\́�\���5w.�G�#������f�ȗ[���*8+�I��D\Uh3p"V<s�g�xn�YI�D�	���>r����r��4�GmD�#v�R��K�5Q}X.��+��nG�{��V�N�罳T�|�	@�j�I��f�oT��1јЪ��O�k�&�I��F"ܨ�[�a��CV� �Bf���?������°S`q�_-a��-��h���9&��I�,4�df��lQ��]�_�Y��7�Ck-��_xQ��U�yp.�v�kfY�|�h�|�h\��D%q=���\��uW`9�W�9M�9T`-�0�B�F�-�?ک���B�#�7UA:#?���Δ����?���"�p�%4���CYu��
�jF�9d�A����*���V�{���ČL�M�g�F�u�T�V.j���3�U�낮��k�oЊ��@щ��sTe��F�Ì*��h4���͒!���LC���{�N�a����@&�ؓ:AՒ�N�FT�=�B��Ē�"�ZD;7V�����ؠ�o`o%9㛗�:W�,��h����h������9,�)�q��6��VK��뺿��r�#�+�ځw�'Y��9&�,�b��`��h���Y�E�}6
YX3��
�N��H�j�R�*?��߁^V�N�����I5|�Gi��/	>�#���Aıp��j*n�`i�Ҽ����:�4ƃ[��¤Q�
������hV�h�='E�Ph�I�"|��X�rg����B`�U���;_�1.e��p^�NϞjt�T3��\|
n|�r� � ��*�I�L��"�}��j�X#$��O�R�X���
Gr����Ds��lX�9��,)��������C�N���6�N���W[yCRt4ĵV��^�tƹ�boY8���.<�ߝ�+����}�ָ�u�8�l�XU�3�E��R6��G�5o3�>y����)ɟ�ytոc��}��_��t3�\e������))�v��� �a��v2 ��sMU�iB�����J�QDjF�k�X꯵��:;P��^ы�a�X���/ⳤ�YIn?�|7~�.����؈�õ�N�]�,հ:
R����|T�q�p���������כJ�n�[��QƗ������j�tw=}�h�:��4����8�T�`��K�,���t?�3�Z�\R�T�ͅ�6�]����>-m~�'3s�8�_��ەS���*�b��!��r;"�5_�M�x�kʫa��F�C�X��'�b�,I��ſ���\n��Ž�X�u$.��ފ�I>�Ӻ��j����WUp��[�u̠��w���u9��u�a22�u�ڥ��V��gx�����Nt+5��PN�$���<�\	���	_��1DߛT;y&�b=aG3_�8V#�(��!D%b�W��&7��� ��U+	��
H?�E@�5�X����6@���
�4�bǙ�����CN�� I�۞�
�m���S�S~>���g:&�'E���@ ��1%�Ȱ������3,)M�8{���޻�H �0=62A�A~x�ze�K��x��N�&4�9Z*:{�.�X��S.��@q��q~
]��K�=Q�j�c~�޽ e�v$u�>-o�)�a�2�Œs�ٝ΃[������C��}�#M�:d��ԔɧF[�������R&�=��7��,ƽ81����K�c�U��ݖ�˼�b6�;=��쵟>���N�3 F�E����{�!�{7���K�A;��ږ�d�A�W�G��nM�I.��0�)t��q#m8�U'����P8���ZZ ��6q�K֕s?P�t
<
G.�/�~t~�$���1Z̬X��Io�<���IHR�o�=��`�]U�2IQM��,�T��nӑ�0G��i���a���u��4d�x�$K�K�2�vp񪟅q��E�sf7�<A��HX�uV$�Y�,^��iW!Cl_2�Q�ͤ�	|o�g���`J~�i�H��d�+S�M��ӊҰ鑈Ό��}�MV���[�8׸0��q�� ��h�ݾN�3� �ٽ8R�l�D��e�!/V�M���p~�!�:ݘ;<]Zf��h-EQ�0�T���&��t?�
�q�*��5�&�y�?F���@�!@���@t50L��v��T7'������X�X��P�K	�!I�!�fqԇ|Ly�����vi���׳>�|<�V��/�Cm��6˙��[�m�P�o�)^4 �>���z=����F�����J��,?����B�N�Az�O�n�VZ �E�)��;�)�if\��o����E;�R�����+}�U�̃�S�%]��+e�O�Sl�3�#a��4m��o�%2�����8ق��6�X |FH8EF�K41Zܱ�bvC��{~��<l��Z�0cґ���:fwkh��?��<[{�?<�`����!̴�D��o/��,����"{��5���ԟ.����&��@e�>���Y�W%t܍��y:j��d>P`��]�YM%�c�=�����<�z;f���J��k �?�GU3[��Ӻ/�_)0ڞ�.��_����WX?��gV�B@���\�q��C�C�8���Uz�w��c�QZ���?��t*?B����4�zm	_lo��|�����K�~p}B`4(ɼ���0��5n$�-��S����%���Eߔ̅����#Ib���o�F�^d%AEز�d��!�Q��G�$��8)�����Cm����^��Yg�F��8Nub�UC9L�~7�p����9f�!7�����_��y`��n�o~���k �U�F���*�wy!�9�"A�e�Ż�r�[=SKo�[�.-�
(`:�f��y9����~��-����M�N�Y߂��Jm�tI��x�v(��qH�~_V=�A�$�u�������>�,O�� �(��I�9O�Re�c�m��ҩ���3�x 9{�cG~�=���)p�/'�T<�߽^$���7mxRU�S���ї�)i% &��Kl��Խ�CZp��W�nFH"7=@�ΡV)y�ӗ�`҄�}�AK	��I������qZ�=]l|���׋�SUh���@u�ۈ����`زqيׄ��#������R���B�6�L���S!Qћ�c.�&:6�\���&W_�f��/���
�M-�唫���:;C�gMt�V��;?��+E�
�Z�������)\��ez'X���
L��`x rEzꖆ�����N����������+�h�:��#[C�ȵ�9�e���5��N���8V<|�����;m`LP)���]�M�y��w�S��V ����n��0����-p�Sk�wȓ5G`|<��tm���]2��/��v�q�r�� %���?��,�X�����쒱�����E;�����fQkR�ti\���<��񤭷�"��Xt�`~.��Q�Xxp���+0,�ѣ����������O0ޕv��w6#+X#��ٌM��Y�E�G�ʶ/�_��L8�����9'b�.��/��>�ʁ����4��gT&��т�~�:�������]��]]w�qԇ��/;�v���IJj��G��?zG5
 ����1��p����3tD,�������`y=����9��J�da=k8������Y�fI�Q��z�0�7� +Yϋi#��m�9 �����7&����z�5�u����Lv,a�/Ap�fŗ�-rmq��{��R:���^nkڸ^�K`��0B:�V�+]�
�Q�$+8��>?J�H���և,Bg�p�����G(�'y%.�6�NĨ��Xٱ�m��s������N���yX㖪��oA'x�ϯ�������79� �u��3��=�r�r�w�q�Z��f���r̂޿��z�d�8Yخ�9�!&y!�������x�����d��SՏ8������B� J�د����7�@�wM~�-��'��*�=��esC�O�ubr� ��jx�=�#����g��Y:�D���j2�R�2t�A)�����Sߙ[8��M���l�^v"�
Ͳ�䕢T|��LH��ठ_�i�R:��>6����ʯ�O�u�p���A�8cV�
5$���0������C	���FK�e�	��
�oW?D�j�b=�Ԧ�Mct$ zKk�Ɉrb��WV14_z'	�K�s�6rq�ç�7�3�4�����k����� �)��	j��\ׅ)�s�s�� �y�s����5	8�K~M=y<)��N�A���Ǎ���4�6F��ۖ&�&�5�K�}c�K<\������F*��"���t��:O��!�	�R2����	���G}20�b�yˈs��1��LU��/j*�z[�7�N���T@$�9u%��j �^@��.��s�G6`qK'�+�;�݄��3��a���������dn�@Ѧ�����oA���~��6���dA��_j+d�J[��S=ܘ�峫tO���xV3�n�����>6���)ߖ�PT����q~�u���d�nӃ�����օ�V��v�O�O�J��ܬb�
Ŵ}�Y `��YZ�2��0L�5���%�Q���t�����H�t7��$;.8Pe��Q�eؚܸ��qDΏB�cx�Z/	�������AoA����c������N��^gk���_| �
/Z�����y�B�����R�@I�l+�Yiu�n*��bk�����%#\؈` �w!
�(-X6q*�)���q���#�����U�W��0���
b��*&�[LWR՞exT
���|1.夨��(�Ț0��{�nf1L�~ �0��b���H"D!�7�����ˊY�E�f�1	��U\L8�vu���w�S�YQ!�Y��^�w�%���ܻ��ѱ��Nu6)s����/�����r�Fm̀J�~��.��c��^�u+���s�oN�pZFs�_����)d��U����'6���Z&�T=�ũ.[E�����O�T�S-R6��}L��?���ƴ>J��%sB�?lT�tX����+�\�3�OeI�y'�3I��p��Q7��{�;��P��CD�w����^����lّ۫@��)@wT0�U�ۑ~2k�<��-)�jM9�����b���w�$jM�4�|��g�Ql�}|=��� 0Ǎsȃpg�2��J6:��4k���^�0�l�0�?��h�ʲ�~=�$&Eiv����l�+��y�NK�q��z+K�lv'G|����k����%%��)����L�Yg]�O�.���7�u�ÏZ6�\����e��A���rp�����Z h���\��=HYd�t�9���X%ؔ�^H:<�>)�$g���5[5�i��=��1��.Ӹ�l�YE����zR�~A��H�*�^,�j��%NS��⸁������>�@�KR��~*�����_N$ϔ�wm7���\ʄ���J4r�vLJ/��\ G2$�sŮ��5yҶa#H�F��w>�k/��p��1NV����_����6�D�Tz9_��۫�A;4��O�/����K��m���������F�sa�����v|�x� �oX�S�.)�tҽ�Wb���*(9��s#�����@**�l�������]=� 2]��m�H��O�b#�;9i���n`0B�l^Z[\�\��P�7�)��:MʎAۂ{�`1��ʭ�@7� 'A�T0����ʀ�ƙ���{��6<���;~�����P`D޺����=�4~���<�7�
��=��K���cK����3����P�v?E�.Amw���¹�"vw�^�s36�89�(�i��ڙ��q�\��l�`���:}�ɷn�����7`�dU,���z_���>B@�1nn#�*��9��k+��+����ư'aAc�"7�3),Ӻ;uv	f�i�L T���E��C�ʍ����<Ϯ	c1X�Z�&R�]Tz�k�����1��_��u�����[����)
��ٹ<�A�D������,�9(����pd+#Q��c���IgI���C�Y��hyq)���<8�j:����uM�l]��&<�/	C�w�[�H�:�D��� �bł�T���������Ӈ	Pz�J�{�n��[K}A[��J���<4�7N���d��Q��?RI/������}���tT ��<}����G��a@j��!9��/8rxqྩ�v�!ҋ;����`����"��v	�B��+�����_���wx����F�C�砓%R'NǇ��?��ŝ��m�t��B��?ď�`��������u�[
uԺ}_�9�G�����^��R��〦��a�G��Sr��y�d�r��Ԋ�ۗ��3��t�G?�Ė���x�q�R���4�N�o-/�kV�6�vT�0��g�~,�بx�.�LC��zbRN����OJ|���r�w��}����缾��!Ұ�4(e���ԏ�g'�<g���jcLsA�<� �-駟Z��̇ZӗihG��*��Icy���⧎�!Q����e����TR	o��1��I%9GS�[K�U�К3�::+:M?���,��#灪ɸ�f��0;+G-�}�b-�x��F	�:B=JȎM�P�R(���*�b)�~�KS2�'�y���}8�Rb�1x�X�A� $
��n����[��+���%{p�e,IU��Hae?B/08��� �M�$����t�
����2EH���@�� Yà��}չ�X].5�]k��������p�QD~�H~55?�SN��7�[��� �,1��Rph�����-��'��$�qt�k
��#��l+e6k��� �hࣀ{�Oc �?Čs�f�@�w�����N��b�3��k*���䬓S�A�6\�D��2�7��Bֻ�4�d�b�7����
`^�F��6��㝻��AJ��2\t[�a�v]�(�p�SGZ�f���n�ج�D�C�"�bԺ�Z'�~�׳Dr-��t��԰'�KX F�|K����\�fR�1-<}�K�PL��e�gR"Y���`l�ϳO�Pڝ�-�uNf,e�v�jgY��c�{���֡��'�'e"�]�$�_%k�@=�h���Ma�j�����&��㞴��,�����țT��I.CJ��±v��T���X���RP�;��5u�ؗ����+�/��"��=�|��+r?f�ȟ���HTD:�Ԩ�~k�fM�b�1y��S���m���yx� ��-Ap���s�ҟ`4��{��N��-���sA��d-ͯB��)�o�VgQ�M�6���濲(�|�7l 3[�nb/��(���ij�[��aU2H��ո|2������ښA��x�	 �����Nz��ϱI��*���)�N*���!�ڏ�.�1����z�f��,_���+Oi[�[���!42ii��"�o���ř��Ͱ�4�e	�(vC��-S3��M�1,ǉ�'mf��o����N+��� �^�(���WIS�+\���d�s��!I�("�
��6Z,�S��c�&��ʗPb�=���R)�!ip얨����Z4�@�3��(��a��W��\1�/�u꯷���4�	_�g�N��bq�3M���E[�$J/GUq��>2������j�3�	�����3�E:N��eN�t@/����q��m��Ԕ�p���H�ˊ�"s��FF{�d��C��?�ޑJ���Fq�;Ѕ-+��X�b���F�
�ې�����o7n_-�x�xB,�M�ٳa�p�El�t�O1+ou ��-�-�͎7j2˜@G���������Ƿz���%�D��G����m�:_Q�pBw =�)�_Ѐ�$�T�oTju����M.@��H�v ��)xC��C��S�?df1�q�NI��	:=������b�����1/+9�(��&�ά�r�M���F�K��8Dr�Rz�OO=T�a��N-o���~��ާ�\��tJ�	
*�z��Z��lf�0_
"�A<L!^�݋��oQ��ES]�y��6���yT�jO\]��z���/�xў����7�r@��ʵ)&�ڔ����O%���y���e#�)��m({�ߌ�թŢ"�+F�ٜ��d�1ЌVO��p,ͫ�S�0��Z����W�9�nD�Ǖ�$�hO��9i�4a�hb��PIK�5#Dp�}�����ы���ؠ�sIGv���b��4�ߩ}-�)0O6=��C��޻�iE��#b���?D���#������(�nSd���*�FV�q�k�j2wv�n�m3�yI��>�-t��n&P0�@1�Y5�#�ҧ��O���N�~��V�AB��	��G�B�������Xi������gb��z�L�0+؎�ɼ
	�flԨfH݀rg%U�K���"�Q"�$�xig��z�����tPAֿ�s�۝�hq]��0=.,i�L���U%��P=>�/d~�H_�P��B��M��a�7���tsW��wnF��e���\���1O�)�EP�����&�0C��Ӛ��1b䥅�5�Y���m��,@Wv�T)��W��:R ���=C���o^`�'���5�6�x�T�������K�+�3!��j|��''F8�,.̴~��Pr��މ�l�	1bޟ����R�W�>�>�:��2���2>���st���Rd��.&���y-����n�$�8��h4�E�[�O��6>QZ.�q�i�a(5x��M�F�T�K� L������΢9����6Pɯ\�XG���[�0vط G+�c�+�Վ�5� �3a��e�Nsq&��1jꉑz�,�79������L���"��'���H�e�˟`{�b��ǆ�lxV;H��,� �;t>����br�F?DN���3"5 ���$ʝ��lv�O�BCr��7�P�D��|���|�5d���0�����x (X�	3NWt�(�j��pK=�SC���!'o�E�h<��k�0�m�ڱF�Ў��f�E���u�
T����_���nb�w��c��Kr���|6�Vu9Ȍ& ��X7NY��۩��o$iNi���ɻE���l�Gс΄����Asށj��p�K(�#�>�ޗ��0}����� }��x�0�W����T�N������u�[������T����lƽ�+��y$�:�WVj�(V�3C ら/���n7��J�h�E�  ��Ԁ�"l)��Z�/��cC�����.��Va9���̟<�n<C�\D��&7�4.L}��Βh'J�� 7'���#��60
��$���d����Âc�g��]_����w\9g>��N8�jh�g�Lw�9ʶ.�$ΣZ�II���Y���0��r}a��_�����6�pF:��"|�"O��	�p[�M޲�z/��^�o���Q�Cbi@�	xKWӤ�*������.�%B*2�?v���q^Pw��Q�4�3D�W.|M�B��.�αF'�Z��뛲\a�vIޛH�W��C�Z��Eb�A��:�GΦ���JIƱ�`UƏ�]D�U�xj��דY5��ج��, 5�;GsA��J���3����U�*����������l�f�|���u&��U��;٦ڑ4$?�RAv��2|�.�lYt�L�A-Y[���p�\
9�ky�+�.�IH$e[�#��kټ�ZY�j���]�L�{�}�� ��K�I�MHs�U[Ѿgc��/������C��$��m,�Z���+	R�9�۶,��x�8:7����g9�S��.Э����5�v��cD��,�8O��j_�»��x�W쳄��{�s�ez�hh!�`�Hi�h��/���LU��M�
4隞ᡤ"�����`ބ�v{�@�� e|��z��D�Th?*gr�a.�eHM���5�u�3�ȉg�qQ:[���*��t��\�ʩ�Y�����m@얮��
;�qD�1'�\��F"�jb5��j����YP���a�qN�(��1ۂ����/��T�����t�"��/'�9��,'���9�r��Lq `���R��yE��#���6~�6���S�'�/��ҶP����&��#��,'�U��v-?}G@鞸��Lo�Y���`�����$��|��L�s���v%��J����Ѓ�;��Z���}��;l�>A��\hc��>\`��?C#Y�G��p��'EW	/1�iK
���Oa�&G�1��'��mb+2n�ǒln3Ér�e�ktr9;,;}:ͯw�ذa���"�O�kWf8~ke5�<v��j��栲�ˡ�"�A9�LZ&�X6����ŝ�>�!�9��k0@L���ڤx�8�U�m�H�ؖ*{����8�>�C��k�$ޕ�D�>Ϭ���X�}�VƬs�A�a�kxe),���8�XB%ؙ?��A�(dL1H�rK'����}�~!��t��b�[�;}����Ǡ�[(��A���>m"���Xf���1O�i� �ܸ�Ű��|RH�WP�*����G�l	&.\K�op�"
�2��+;���ԫ�� ¸��eY�ݜ��R�7<[�I:柌!)��>8��#��Am���#��Æ��fl�ԯX0�����u��m#� {�-��@z;��oF��?>��G) �P'|��o��i��	/�"�������B$����<2�]l-�D�<	xIX����dܒ+`fxiȒ�^����;��46��W(,��=�!mC���F^���m�xW��* �4Ѐܜ�~��`
K׉ĝ��㴕�z��_��o�퓑�6{��DP�H�d�?����>��"0F��������K��e�71>�����RS�%`�\���)���@@?�y�J��U�xR�c�H��tm�1��[�!�����y�!����S�2I�x�=�7E�z����u�[����=a ��8��~s�A�#Q����Z������ʁ�ȹS,��|]�ـ���8��֒B��}/DCz|/�i�x�:;�Rw�/�z�î�p��h�h���L<��N+]���`5�0P{��S��� �=D�PvT���_�0?��Z���,�-A I���h^��M���O���C|���W���.����\M�c�	����R����)Y�2���c�ED��9U"wVj~J���S����N�|�G]�F��x�F@?H�$�E��=�X�(5�A%K�o��r
�N5����Ξ�6s3�!$�7@���t�3;C��`8�âػ?���c����x<+�>p���w��@:Ei�!�Zw͂쒳C�_
��(��MZPp*z�9���),ڮ�~�]�pXC����ȧZ�B#�ضK�h!�K�m3�ɥ�AYߒ8�1�f��� �L��>�譭I�o��6 vBOd���V/SLI����1$K�\��+�_�)����ߔּ���"����>�c�6��0��gi:_��2\(*ˎJ�"�J���w/��M��w]!*�Q�Y]UE k���>'!a2wO3����Zp(Ǜ��m5�d?s�<e�Ѥ�0�Z�����]�1?�S�E��Z�@Y�ɷ���T3�yjC�S���s%��i�p���9%��̉�L�� �"+��¡�z� OFc��.^�]><��`c���|n� �>��闪�1�C����y@�v&��̗=��Xj7�Ƌ<D:�������5m[�y1���j�a§����K	�hBZ��Cj�L$�I{�8-�]d{�͟����TŇ[�:P:�n@��p��Y�N����R:34������a��n��3��^^N��N,�8�r����(��cC�w��p���룟��
�QD� �?��H�+�i�����E9�J��׏ ���s�}��WMm����9��*T�yU�9C	{�z�F�q�ߩi��,$#�@p�V����D"Od����=��\>�$"�G>1�j�֕�1���u+l��9�+r�J�1�c1"�n޽�b��Wޢ�A��
����=��
�~����t��L;(��v��,���i���w��=�Ml�iH|JW<(P�����㿁C��VG7�cN�����ƀ���Y����<\,Y�^���)�� Ō<}J7,��q�V�,�����(V�BF����.J[g{��FD ɲ�����П�6-.6�}3�7�����P]\J+�H�QI�pN��;�� N��s��m��U/؁�%�
8��̀����}�L�����lcԽ��	�M�4!ʼ~0Iͮ���o~�,\M3p��+J]Ru�#�4b!g�{���4����i��((�Ԙ����Y�q�_�iq��]�@���ʑ���b W;�]p�0�3�� �Ā���$h�2+�5ɝ�!���l�7i�	M��T>�Z�=X�ES�\tq[�nY	�P�i[�x��2>��j�VT]Q���\B|��4a&�7�t����c &����\����:製�Xٗ=|6B��D>���ɔ�,Zi	Y��c1��o����說���U�˽K%�iT1�뉿�g�'h�Z��7Z/zw�H#H 6D�DoT��%���gV4��Y1 �e�d'Ӯne"u�_@AO��,�rj\�@��n6@�*����? z������ڛ��n
�G%ء��3O��Z�z��?ힸ��rRw�W�f��2RV�ތg�þ .t�׵��B�'BA�ԉ�	".+�:-{eQ`3�z���fCG�],j��Mg:Ե�X���P���W:�~�?���yiur�h�E><���0�5��$�,�:v}�P�X~n��ތ���6��R7��V��dJ�U��j	/,^\&��{YU�C��B�j��$������4�XĖU��4�i`8~�B����0�I�����y6y��� �dj�K6�ٲ'�����j1Rk��,| ϡ��U�M�+S�^��8���Ȃ�T��>xRZ-�O��'ɪ �^+I-���41�ST.�&��떌WѠ��^|m���fנ-���U�dy���A�E�c�d�y�l��*��0AB �F���=֯ݮU���_�d �0~�a�9X{�C(��Tva�=��c̨�	�\"��>�#ɂm�Ԅ�d
�LyQ�@�Em�x#�xnͧF��r�=�\Z��a���N3G|0��/I]�=+W��	Ӧ�
F�­��h����`��;��e�Ѩn32 �v)�h��������,.�^e����	ؠ�d�N��V]��	���7���������0C:�LoLgB}���P>�j����Z5�8U-���Mz�4�/�{��ͲW$={j#�A3��������|0�r`TTm	��,��kA��'��Cy��+�+���D���&NL�Ӌ��fES9H�a�����iW�f��[�r�U�!'��j�zo8V`S�	���c��] +Z���P�j9~��%6(�0���-+nځ��X���H��J
 ���R���FDtƉ�uF):%�'"��\
0�41�;��Y��ݒ�,+`ۇȇ�Ցᄩ���'��v���1���)�V�;,�R��h�jZT>mei(��Z�0�QV�"�hH�2�K�B�s�_d��F�U7�<Ø|�z���u@e��ǿ% ���� H/]��=�X�ś/��#�_l^x���ZCE��9�uޯ|�ZC�Ը/�T{���r?��3tBp��(.)gCZvٖƉicé �OGwW�䦹~�~=s�c������43��r�&}�yy���àZ����;�u9����l�-w��-䬙}�iuw&�0!k{��M�NrG�n矏h�Ԩ��QE����	�h��4]S?x_����qX�L�?�!��l R�g�C0��� �'TA���K�jm�&�Q(����^�+�����H�΄x^.�����,PM�c[k~`
��^x���>pt��GL��g��G*�����8A*�-�� VЌq��Ù]i�K�������ݬh��
�&էC���dA�0�[�e��_;�BEG觘�2w9���7�[-x�����aϋ��-@'��ؾ2 7���
R;� ���ϸ������p �[E��9�Q.���U��7s��	���^���Q �,���*K�E��J�%�V=�Q�D����ת�鴎əU����ۚ%)���`J������b������g�p8�U��u����zb�!&�|t1C�x�q�̩o�we}�s|�q����-��S�]H���SP%F�]�E��J]#E�75*�}��7	'ٸ�R#v�B���Q��bk4���̔:��2�����~�V�I����a|G�S�8��-����L���OG8D �n��X�+��ս��
�W�ᥬ,Q�`�Q���Y��QxvQ�$�͉�*{���ˇ��Hn!����m�����h]U����B~����x�����`�=w�ĳb%Xz��Y�귔��Z~���⋈�Pl��>tE��K�8�CıH�^z�Z���[���b�zom�H��Oin��0�- 2���t�F���Y��E\�i~qX��G2q���se`��Շ`<6��<&�h� K��� {�o�{�,��@8#��{�E��:3��ͨDѐ�n=��ě��c�_��+�s\Q�~	�R���r��P�;-���1�1����H0�O�!��A~3D�g{���!bX������_yb/�wG�E?:����RL8)
�)":����~L���$Ɣ�֣��Ե�s�P���M$�ӓ0��u$���@L�o`��� 6��$n�#��Q��)LB��Y�p�&5%̕+B�(��W$���K����̂���f�!��]���51�y-X�1�8~ ��5�H\	d���q�_M�����W�c�×͎=�	�Ң!!�3�τ]��z
�5����^���Z���L��hO���Zo��1�,HK��	�ٝ��ǚ��iA.��lTJ�D�xP6+�o���iá�L��6ICU%I�KA���CK��$�L�XD���k�P//�<�%)�͏�Kڎ�qy�#x�)]��4Xb������ޑ�����	�-m�{�����I��a|[�$ z�A}'j��O��bE�XwZ*;Ї⽗���֑�W��7l;4<]?�5�¼��c�'<��iM����� ]@-���]�4�~r���^��C�B��W%B߾�7X�bY�O��&�ݫ�y��.�:D^�����V��q/<��}Ks�@�r�ߑ��dD���X���U��D�j@�n�����y��q����^��c���,5��N7���p�p	�2�>���j��~����&�G�ߛD�����r�^O*ޕE��Š��b1�C"|AE<D��?�ڌ��q�_4�c +��?�
�p.�I\��Ҧ	[&K�����[���_�Q�|\m�5.yT��nFPP,����N�Æ��>���~��`�`�~�����\�3;��)'*{��J��:����������pv� ��NY=X�s
����wJ�g����c��{r�l��Pdжq��#�Qs�u�P�O�k��j�D �pO�E\�M�yu�<�˛^f��tGO<���
��vg�n��H����_���R�_�Vߒ�wث���bY���Y�KR���$M��Z��厡��m�Fӓ�^0֟4��z�(��w����@X���qԉ�K�G�����!tp�>��i�Bu5Z�M?��e�UHd"[��G̉�f�����R��Q.����d��JY��x�G\?�O�KA#r���Z��Sd�m�����c-A� ޴�mZ���+�F�T(�y�%��	E��Pv#�M��.K��7�c֍j���wi|p�������)��H����5�e�%�V5f&\�ZX��ٌ\:�*Z�㲸�B��~�\->�� ň�����0�6"��	���A�V�)��P�� �Q��:�i����YE+�Q�65j߾�!F���o�%�{��B����Ų�i�x	5�h�|��5X�!���I��X\�]B����{gl4Ú:K�#�E9�N���e��1:����k�l:V iu{L�x�Nj})���w����fB�+(؆E�Fr��F*E�<Ne���-�:B�]	m���!���^08�=��eB�S����g�-��|ܨT����6�{(�
����{}�E;��ϕX^�߻`��=q�M�*�T�-h�&b�h���Y�d��h>=]t&�����}(�����c+mRG@�R�i�,�{�3~JwPY�v�Jn�i_,qg����_�$n���0�q��ǂ.x��3J�E��W<0�M?�����|�O�&���Y5�+�U�릓	�y(%o8Uw�Xc��x
_�����qȁL�U+�zȺ'���188�
��`��ePAm��m$��-�e9�pG��cOU�#�+&5]�]S%i�����0��Gz�����s�&&�i�g�ZZ \�`e���9�Ub�� ́�����C�����V�� �*��w`D/~)��ˇ_��S�"*�]�\�SPI���(M��1b�
������+��HG�����K��\�Z�D��ؼ��"͔\�k��= s�Ϫ@��ڗI<��V���������w���z�SЀ�9�{r�1�����|pQ�2�T&8�����UD'c3��:uw�坈 �{�s��Zg�ɴ�E�5������c},	Z��$Z]��@*��F�tl����I�@l�m%7�Z�ߩfM�|Ur��-r����ˢ	��V��^M!$w�M�Q?\Q���>d�c�褫�~���\�r!��^�`��J&Ѕ_Z-���t; �{�HȤb�������ٯ�tk	q��V
������w��^� ��^.
��yC�����Ӵ�a�]�rY���9�j����p�N�j�_>0����+�X%I��S�y�+��ַO�27.7�2i����ȯ��!�����uV�-nHL�,Eů�f:��:N�� �w�P�p2�SƱ��$�УsxĂ�>�;�XU1�Nw����*aYcjA�a�ش�h��C����t"3a�C��5��������TʧkUF�E���?M޽�/O�����i$n�T�� t��#�pyw��:-�GP�7�mH�� >���QR�?����$����3�#)�����Hi�˓I?Fp���I;��ŏ�Y�]12�����m@�VޜeD��o��ũ��
�A�r\5�H�3��8�o�5�Ŧ�9�U�-���8r�کv
I�ei�K����_L2�N	�Y�(r%�����,m_ZAk4�MN�*>#q���m������4��N�l9
(x�$J�4�!`��xe�8���^�}W�]�_NaQ�ۺ�}!������ƃ���E�����|	�H�N �'�pC�=��8QE���c�w`�9v�t���(�t޼�/�����y�F˞�T���ܻ]�R�����WVg�n�Z,=1�)�k��Pl��k��1.���aQH���b����-����D�K���m(Y��9����'�B���q��5�M`��j�z�$K��{L��]"�ۘ�>v�ܴ�R�({a���]?(t���1]N���2�d�ᔝX��S��e�v�B~]�o	,DΣ!��A�FI��p����'h|����3���*VUdg�_lw �û�e5��T�%<xhq-Ux�3�I3��yT� ��5��;ߔF���� 'j���?y鵜2#��,TV��h��,�N�HR��Иo�����S��1�ɷs��@�r$�{�sE��~�E��.5M���3E&nn^%{Mm�86/��F�Q#M���u*�GGZ@�KQ�����m\ÎBl�08綊71[�{��{�q��!r�`u�ɴ�5�:cb��4��F�7�E+�n����e�f_�(����M����4�.�!�6��R���G�-� ɕ+O� ����Çy���5��ы]<K���G�4/hY�\�:���V�z��f/Mh�(�]le��`����ٚ�0��00<�����u�� Y��J�l�1���׋�-L1��i;��߅JB0dsД�Ƶ�	�%��	-� KV�,B��V�������v��$�4#���fތ������Y���j=8jr�g��Ss�@��MU�v��q�HZ��3|A��1�i`	�Z9�i�Y�������=2~@���5h@?��2��2�ò��zW�Au^q�5��hQ��2��B��}/ei���6�yU�^�9ˉ�L��5f��$�T|��KE����U*f��Kre��q�9}DT����ͺ��"N@�L#��2,�1��ܲ'�w�I����O�	�z� ��0{G1�l]��Xw.r�]�n��՛w�n ��x*�/^W�*� t���"ܛ���p�-M7za��$�����p*X9��l�2'M�Ic�;�r��`��視W�����y�����g�Ud�d�A����m&�A�#���Eٔ;+md���(^a�􎏀,@�uGn�|]�te�ATң�D�7�8N[ ���b
����`p��@��P�%�A���p���Q�3��@�p��펮��~ܲ�-�3�9`�kF�U�c��X�+�6F�3��#��Pmv����6�8�<�x1'�X��:JaI�|��80�ٻ)hTp�x��Z�*i�R�M�y�Ǭ@"LU��9�bI]$չ�ثm����O��A�cF~���&2��
Ap*���q�3�p��㘙��?�����D����J�7��?=Q3*��e���]H{9)/�F�g���+��ƽ�b�G\F�z��ɘ�m��Z*$F�߮!����<��gP.��h,"�ېX����4y�?a��U�p>����ݓf`�3�v�Q�ł,�l�nD�S���n���z�jXi��/�� _ꎏ%t+mH\Rl���#�W�������.�'V�V)�1�.�Ŕ�?Ei����y5o�mfO�W���WT�"e�v��~؃��t��F�.�o�<������ �=ç�q_,���;�N��S��TvH���8*��'g��@x7���}ٛy�lPڹ��?c9DU�N�:��A+���%:�+�Rh��u�aR�ס c��?q6�4Y�0�Y�0��}�Y�jx�F�6H{E�%J{�aHʘ*�l뙜ԋ�n:]P���N�)b�Tg��I�R���[ړ�)	,P�E$�Nؗ����:�y�-�$�g��v[�V��\kX�-��k�=/S�+���8�OAL|��7���[3C`������^�����U㘱j edOB�T�ҁT>*S�̲%���~G��o&\��s�5��S�'�&n�.	���Z��r텫|�����l�[����~չ����#y	�!��i�?�	�������m�Y0�:}
�U㐺Ĵ78�߷������4�������u����۾�bJ�q#��"�U��.0ඩ�6�>�h������K�?]�B���{_����h�UM�!ס��آi����Q��f��o����*	�Z�$1?�nu;��Q�)B����"HQy��D���/J�����ӓ8M��
'f��?"zo�)E�]:B���k�H�)Q���i]�+O��T�\6�Ǩ����Y�v3u�\�/^��'�-�������������w���kmYeͲac�\��q:{�&����A��D��%yN"��Ù�2�����N���K�O1eC7;���k�2��4�P���rۥ�X��������ߊ�z���q1�i�A��ִ�*c�~=�Vl`�-|�sm��a[GO55㲨/�z9������Jnֻ,����y��1�=�^�M����4d	(c�W%�'�ǃSIj�;'�Bͭp�=����Į45�{y���#�9�xϞ����"=\ڬf�W&��Ty��'��Q^JRy���윏�@��F��)b�x@�(j�,�6N�ۂ����傀�[y(-����/[�RQ��<6���@`t�y��0�Rv��{��9����a5+�-�FO�I���6;�\jZ29��Ԭ��v=B�<�,��!�:���j�n����N��/��z0a���?Bv���j����	Q��R���Э��O�� W��=������a� *�fb,m��L�G�W������߾��\������,L.�ټ��!:���~u�y��{x�.>�6d�-*��r%����}J<� �2�!,ث0̮�#s��vA1^U��Y���|H<3=r\?��y�<�WI>�C�mE��=�{.o�4�T"\ �@C�А�4�Y�)K�=s�?����K�^��sӠRM�v
�UXFxq^,#)������b1ބ/��%[O�*�#��K4��m\ǎ���z�88pw9-�Tt�Pi�ix�������#�x�Ƶ���|2��cwn�Ǝ���E��>n�0������FD�o&)ɦD��J��k��me�����@�1�.b��n"���{h��2o����������!��c�C��Ri�FҎ��.�gA���	W�ƩN#;Z�B��,�}�o{d��j.��z�	w��=hl�� N����1�,��H�����ǀ��c
I0��P�M*���B���\�q���ۄJ90$_��r�/9P^�c���F�`L��<ީ.J�A���F�ha&����M��b�p��r2 �|X�P|�NQ?�"�z.�XN�A���bO�V�\a��
�f!mv`{��Q�����q{��Wh�-��얁!�-2�ʉ��2[��z=b��D�>vW��Un_@�3�D;�֮��/K��HW6aѰZ�?Ͼ̈́��l�3�n#3FHa�l`qHj���,d`<>���C]��mp[(�TSF�6��Ed}��<�ū�֋@��(����������JA	q�=;L�#�2{Y�\���;�6<\y����eʲ�p}�>�x��x�S?p����(��$<�.  ��8���h�#?�i�'2�Hϸ�4i�����a�!��I�-��	kb���8����~�(VG����p��7ic P;Q{z���׊_Я�Nj�~h�/���H�%H�<��or�u�ݖ�)DO*G��H�{Ѩ�p�a1+P�NJx~Suw�����-o�'Jx��UCQ��7-�E�я��))�J�^ ��Jk���3d��7pj�ǘ��-	�pK��҃c��_����M�T|�Q˞4��]��sf)��Am�B),P+m�K@K��n�[��<\E:�S_-o�ɦ����'$������� y��	��P��jE��Ն���s�7<-�5�Ӽ:�[={U�y���1��MY�5{wI��l��%�4����l�O��)3���J�@��{�o:S��_b��κ�4�8@x���bR`p�	�
��
�Ǭ	��2���^�;@�����~�RN�5��TSb�3@=(�B +	�n���-�Ϳ�O��m���Q�R5�q?�PW:�u�WRo}Ո?8�m���^��׼j����r��:�CQ��XS��d�D�W�({UZn��Cu�~������ ]M	��߳�v$z�%( ��\�0|�t�i�1!pX0�P�\�J��a�9�F ��\�kF"��^ҷGGb��I+^����Ҁ����u��#ol�C��c��Q�u�ق���XՔ%��2T�=](4 �y�u�ޏID�H��/a�z��ܰ��4] ��wP`�3���Nz@�c��$�� P�K	4C�.檽�N���c-j��4�K���e�8;��8)K�X���V�"R�D"���<�H	�[�-��(]'lD���'E+e/s��V^S%���3��Q^Q�1��44����^&\��9�d9��w0�&u� �!4*463�4���6��_|�Je������A�_��w�����2C�g�=�&�e*�Z�������J�r">��T8��g8$v��~Ie�&j�H�I4�,ܼw�����y��U��ӻ7� Б�+�BN^%6M;��1G ���9�ԤE�l�i;ˉf�阗nzh���Q���BG��ͮ�Y�1�������7$�E*�Z�O�@��)�����yfb�)��e��)r[��P��4l�
WL�"�0W|^���V����.+�w���~�o�oׁs_A ��ꂦe�|��6Ј��/�(àą-������
ݶ�����=ksf��P��Japzs-=9h/�	-�ɣQ�Xd��UJqK��4��K�/i�UŊr�O�	L{5����gpoP��Ѧ��<�b�|�i$�X�g,�1���9�� *6r@;��,��*��+��68IR��m(���S������_Z� @�aXEYd?�Jy��aF��k���DDlp�K���F|WC*r�-G	��e�G��7*�Ūه��H��_������Ҷ-/V�FF���ӝ���,u��8wA�XpMbԷQ2�x}�=�o�=�����h�7[�Vqo�x�ZQ�t'�"�Y�#)t����ϥB����0�g`Y�5��֛)��4�,�Gԍ�7aC��3�P������i�=!����k�ݝ�_�W�C05�������ћ���%�Ó
͈vm	�f��"��.���(&�s�k��oꋬ�KOu�an�v����j8p|�eV����C��ؽ܍���lR��w���y���i����\�Q��­��� �a�"�l���l���OY=����+�P�o�0-��N�l�b푘;�kɑķ��c�>�:Ƌw��B=��i��0K�қ eӖL�����g<���Ө��jk_��
��=~���v�+$��x�h��)y�s����J���DM��Lο3^�&D-|�h�0�
Ok�O�-��:W��D�O3�۽���)��5@�_�R�£u2�Yq4ux�gI���u���G�{5V+B��-��pr�����k��Q�TddpѬ�bQ��$yޟ�q�<���x:e��i$lC��Ǧs�Ag��9��_a���J��<�@,����r�a�<;�kE��śi��M&��ݮE���˾_�����?����������׫.n@�&K\�Mғ��ץ�o��4�
cA���\�^CI�+�<�(�[/�������n�X_ ��j��L*���<�Q,�jϮ����.��z��JXY�����1'��aβ���a� 9Q�s̆Og��29tWX��z�w2U?�޽�W	R������:*ɋLL�ǩ����r���K�Z��uk<��s��a圁��ӟ���R�_z�Y�?�]֨u��F)�����,��� ��C
�<�֎,��>BR�H��f��t :�d�+�K�i�<����?��M�8m�Kp�p ��(���	�5]L��3i$�Q��+�yq-4��@m�U��fM�q�)���H�9tB�B�ph�*2�N��:	�V�2���}Rb��f����R-�ӣdL�J�Vz�h��y5��۟Z�?�-��7`�ᑬzj��|�A�)E檸#��|�qIX���,��8���f�ޥ�>K�t���#��V�$,�]����jn������*rL-An���h�QOJ=���I^�L5k\ʀ�V,!w}��M���,T�vU�4�9�6�{+	�k��J�d� �~B��F�;�[���Uz9�֞� �U���]���|����O2���(n�1�͙���\C!�3�)"u���H�G�f�:hd�r��\X�%��e#\��NRN�rA7�8?�(\�	#�\�3C��7%��g����h�j�\J����q̳n5#=�0�?z�#g�J�������ח��*��3��R�K��~���+�z��7���XaI:yskc�?���!����I�lY��QV�<�=!�y�5d��]V�D���5�Y��4p�]��ttP"�'!%;��Ѕ쌓Qp_��E��$c8�Dt�:i�C�wUy�.FS�X�?.����ϼ�f�����X�0���I=y�����!ߧ��UBJ�TW�i_X%�,��;ٲ���\¸�7<ʇl�ڼ%�7ܐ&/��]���J�&��%�@��S�]<�{q��n�\��H9�Q(���f�ޡ�����6��������{m)1;����&����;�R��7h�����)avy.S��Y�
��h��}Q,ċ���Ǝ�T�'��/q�N�;Z�¶�ZQǇ������Y�u.C�䣸��!�h��b�3����Z���Űd��W~��|e�g�����pe���ex6(.��a����D'�IxZb��\-LojY:�N�K�����	Y&%�g�4��d&d��d�Y6�w;On?b�↛f�y�K�~�q?,
{��� O��¶���Br��v�ِ���9��^n��s�fn��X�ZR/F���mKn�f��)�-��}���3J�o��T��V�ʗ��#���s?��?�̂Yk<�*E�G��"���@��l�8�M�ޕ��W�q� X��<)�	
Y�.4/��cj��Ǝ)���^�A	�j!:󡪥�5��K�Z��#�����m��H�5��P���|
����Z�Ϫ��9 ����kgʾV�X�3a�AMr�~�k��
�h[~�V����t�����oO}�vʰ�m�����k��cg�p�Wv��Jk�'�Uѷ~�?��T��P[5�u<4d�	]�D���g�\fE4b��Oɾi����"������Ïu��4��ԂB�F�$OQo
��Pb��O 0?�c����AWF�}I:y��;;�o7�1Ꮲ�/e����u$EKή�%n�b@����V	�}-n���<L/�" u\/ؼq�������/k��%`5o���a���Qs�XE%�rU�*��	K�NrJN3Y����!�(z�	�c�#�l�˅%"R����zW��A��7|i�b�%�g�84㚺�@�f�QCr<�֬�8cV��CVV5�yi���2����,�P����v]��Ԋ�`��.�W;y���h��}�Y�����?T%6�N�X5� qF ��y���Ԗ����r`���[R��|I����u�K�n[�`�6Z�;;ݹ(M�/O���D�O�Y��G�ڊ��2v��<P*�a>��w;|���}�-v���IX�5o(p=����*��-�Cw�:��w���|\���r�Tܿ�p�Z(?�Uja��
�HR�2�6�2ה�h΃���La��hG����3�r^����(�IL��Ư���˴f^a�Qy�7}����C�]A�_{e����v�tS�h[���sv-���<ӊ�P��oO�b�w�����:�J��^���M=>ɨpY^YG:�A9��<��fy(#5޸�K��u�WI���e���J�哓����Z_���k�&r�E�gp�d����M��$]��>;BѪ�]l]|7vTK�J��`��2��Jo�~����lc.��.|\K��s��t���S9%�lF#5�*߶D�{�A�u;��B��v�R���Q������erG�1<�O7g,^�]�ʧYZg�^;�t�?n�s��,%�JjH���2I_�t��	8�Ⱥ�(���_AG�X�)�	��OS3�a!�(�[�wt�  $e�B��vP��Oq���G��G�?�Ef$�k
���'����$78����*��ƅm�KI�I��%N��	��/��n�@e��I7�o�?q�oGj��-k*��~�@u��r��é���T�������X�����6���'-��z�~m�/�����~q�tm�|���a���a�w�S!l�#�(;���2ڌ����5���ִ}zM}����ۆ|}MbI��JB�F�V��9�TA �W�"Ee�&Pt��U9P��0[u�]���t�{��n=����"b��0�Ͻ�;X%�I�����oK�K���_��f_cJ	C"<�d�3>ϘNjԪ�=w/��n�=�>�=��oql�.��K����5r<Ik��%ADw�}��@�-�P��b܃��������0��B >lk�=NN�V�ԶS��m�*��?G�B�Q`L�:�Z�*�؟�2���^��)NU��֔8�� �yU���Q�h���_���6Ȥ5��5d��j��^��##=,���~O�d8��(N/۰�� 'i£l�粞kD��d�=[���̦V4i���Ƅ�^$.�|*Gƣ������i��.^��p���N ~3�]����.�ʣq�uI���sS��/n�br�^5L-q�_i.!p�HT@����6-�j���uń;c�(z�2�ʅ+��R��H2'����l�׎[P0�r����mS�S����T�P;�t����U���G����C'��X���0���u��t��(�"ݙ�Xn�6ņن:Vu��.r������砐W�,2.�(��4�zQbډBR&s8aږ^ݘ\�b�
�g&Mc)�B4)��Z���C�k|6��l����)?J&��5��[�Qk����e<u�EQ�u�j�]	�ҹ���5�C�S.m�<F���It3�-�쐗���.}�V~�eH���,����J(C&H־ߕ�o��ZΆ2`p}��|�w�]Ƥh�AM�`�%[�z��
ĸ[[�h^�!�L��Bn�*��z�â *MO�D���G��T�������J>C`��G�k�SE�K�S:�k9Lַp����f��0x��{/P���᪠�}�Bj��.����TWG���dS���ªBe�H�S�ټ��ex��Ib����&�_4߱=�ON��	���J��I�����d+�DZk�bύ�5�SL-�&-o`��.���K���X�����H�=k;�O׍�o�r�ߗ�:��7���q3�A��_�	�	����p=v�U?"ɕ�O �(��2��8���61��i\漷i	x���*��i>����!? 2H���K��^(.�b|�������,wp�՚dKw��Hy"�8_��<���g��+�o��-�i���m�(��@�Wq��&��I���d���o�AuM+C�l�"�Ā��������_�a�ok_�&��~~�������e���0L
��L�tC���@�����p�Ը�#�����Kw!�����Z��n0��\�c�fv)t�R� w��a�18Qہ+����|g�����EHF��IT���;_s���"F3��n��K��?�X0DḒ|3���2���(�E���ܮ��=�(���)kz�R�?�k)����qEK�K��mQ��uB��)�e���c��ZtJI"Ӑ؍���\��X��EP$�݄�9�s	@Ɲ�۶���qS����n@�QZo��߁3KTLG�̱��x��ơ{����l�x��nࢎ(k��;�5����)����s���^n,���5�Dp���Ǜ��i��H-&�2�H�:/��''���o���C�<X�����r(���7c%Y��J�K��T�/ǐ��TK2��j+8�5�VƮ��#N�Q;`K��#X+դ��j5�
N-NKz�!� ��-
��52�g΁�j|_A�$��3�`�^3�Ou���HW�/�&+�Bq��迀> R|:	U&�Y���#A��n ��㺿���fw�lG^�����T�&d"c�z��a��r����7Boi��W�"e��R�*�̈́I�Uxkf��tʝ���IS�*�$[ry��ϓi�Yd~����O-���6��՘�'��d(���I���:ɒ���{��0�������p�"�);J�M5�?
��ڣ|�6�
%&7f���*��ؘ@Ć�￪����W2'����T.��&���3}��j�m��W�4DÈ%�C`��d�~�q%�fY��`�<�5�y &���?{����t�W��������>�1N����}e��:��M[�9G�����P)DXE=�U�3?n�#
$J��FH`R�ؐA����y%��Z�������l�i���ΚD��.r(�Yˡ��rƫqIu�3��oKT�E:_�ISVN����νO�
�q��_9��&�:ܺ8�\�|&��Տ��8z�I �-_44����>G���	�y����P�:eU��W~�W9�V-�_�R��5N��� ԭ��P���d#��%U�7Ts1 ��PHȫ���xl�EJ����7����(Yx|-��h�޿`�;G3,�[a�����=Q}�HYU��+��ON6��Ҵ=�|���'!D����R �<$���	�G^6%ɘ&�$�3b��T)����+�յ� ��ɬ�	�}j�3�d�/�T���җ�|F�ċ��O����n�O�8t��<�1.wY�KA��b�PW�58w��r=�6��!�o���킊����e�Z�7ֿ���/��31�q5ӕ��o����(���e��_���6�̬
����}s�7h�|�jW�*���D{�,]_��&�����;T��k��/>6�}߆��NӨ��j�l�{��Z�c<E��b�š��j1i�3d��峾��z^�O�O�y�J���4p�)�;������ߏEoI�ht��vt�ҫgS�z����=���l{���$��=E�H[�5���3�Vr�A�2��5�wF_���싑�w=3�3��I(�qS5P}��g�ou~�i;�%f��yx̤OT�|�ta�o���+��G��x!�̏|%�$9sX��>��jƶ�#��_�W�����J���z���n�v�-�HŚ��Y�Rs�Z�)gu�LB� ���+�@�kj�A�)���{��z��53f/�j ?z�-�]|��S�_Ԁ��*�K5���#�r��]���	/5�AG�.��\�1"V`��	 `��Ӌݵ��,���c�:3t�32�Y�D�F�L��IH�c�w�
�:�G'1���>�!�ڷ�T@Xr�䱼=N-�%sR���XK��ۗ��� �}�d��t�J�J�s�Q=lΆ�ڔ҉�EJCB�!Ź}2hM"�!����D^I��hV�D�> ���T4���醎�l�ơ�x1L��-�<��|J�l�e8���B�2U��;��ȮZ;=yl�oK�ɀq;���9�d�VdF�ۅ�$7��/e�;���]��>>�g��VE�,����7�Y�a��X�z�o�C�^1��� ��)�Mb36+�Q��X���5t�~��xOf����p=y/�sr���x�Ji�(Dyv:4¨� z��J�������J,������?1�Z��mg/3.��ߔ���Qwu�2�Jح�M�,�is��pT|�g��6*?d�=��S��Tp�-uj&/�i��3�?DmIL�˃���6Ff=+>g\�?�����,z����
-�@�p�`ڗ#U�W�I��N�K�{;<�2ٹl�&T_��3ɥ۫���neɠ���K��`\D15J�-����'�2��6��Q���N,���n���Vx���[��< �����|�?U��@{��<gq�Ȑ��C�yU�ge�����E׃z���֓I8'���p�VS0;���h-g���tV�K�(��Qw�e+�2q��W0���g¸��m
�!Kz`�V~�4v��q�PGT��TQ�?_�R�0ɼ�e����V�f�؅�i���E�o����&!e3�6ڛ\�%#R{���'�kf��i"��I���i���ȕ4�%2�	�k���*<��E���S����L���m���-��%z�Q��6��s��u=#�����{Yۼ�V�Z�rlE�F�&I�j�O���ʇ9��o�D�b|<F��M����������������N3S�V���eSܩO&��u�P��ƫ���@˰sb[!�\m_ND#�I,��J��t�WV�Sj�����Y*k�Sg�a��m���R����YYD��|���P�a4_��{���F3��:�gf�����΢��D���� ��ӹ�Der��p��*�f������%�b��l1�е��
��4�w��}������	Jt,>vR�s�Z�ı�C^B�, k8��%O��&�M��zʅ8�����#>iAf챇�	��?BV��T��5����fb���c�r�p8�;��0g�H��Z߉�>O���CV12B�>�5Ek2��!��!:�����������_}�l��Cc��ɡ���p���)��9��w.?����⭮��`��/^�����~�2����cMN#����ќ�X���},e|���;-��	D���ݛ�1��̺�rY��҂`)���&��9n�e؛6����$ �J��/.��\�W�N,es
1«�Շ�`�3�~�y��;!�W�~��ݲ�8CK,˧��oI+�4�K��� ��Q9��?e z3�q�=mR�ռh��;IyWV�5tOB��Z���1����)��	�����"���t�g�Vж��.�YS�d��vy#�S\��J���a��u���;E���	i�`h���(of�u��o��Ǌؘ:��p����A�a�c�ʧ������/�B�(dx����'�����$�_"�/����_a[;0BФ��ƅ�����~�Q�U�ﲺlYQw��>�)�X 1TTސ�+����i&1Zi�̤�����@������iF�q͕z/�4��w�h�`�d?�)� ����<i������#��"h�:�0
Q�*�i���g������8�ZM�4���>��@_�M(����n���z�^�Q�IuȪ�ү�,c�0\�P.��к�VղՉf�s��=J�éG�ܿ�x��� ���3l5��(1��HC6��I�x��ƹ�ח�R1���<L7gK�y�ʨ���?�`^I��s+�XI����p�k�W�j��	�S7e�N�RGIsn�+7��1p%u���#������1�o��*�*�X��qx_q�L>+b��0�����:eЩ��[F��W���yJj��jJ��zea{��ڍ��q�׬��RМ3��{�vZ��/�zVg�o"��:�P�8ֲ��k�n���?Y
��o�**�q:Zn,�ݡ�	6{�Ǘr$����N����h/V�uHI�2���
�p��zD��h� �d�]��L����K��-/͝��d'[��o'f]�G�k�R�K��#���΀~�����o�v������;�<�qe��Tsuezɛ
�+A�g�%���׼L�eֱͦh"��e������K�N_A��G�#b��I8w)f��J��%F��߶>��4A�U�8n�C�>��~E�N��a��jO�[\>܆N(�%h,r�js]Z��t��}�78�y���C=�Y/���h�u�SN�����k�N�Z����[1>P�*��AS�v�z1�VqZX͞!�貲�s�X��{��n�yEq�q@c�g��$Q��.:�9J�>뇽\��y ��Xi6M�8�d�Kv "k
�_���A9�Q=��	�Xw��A�)]�N�΂d=i$d�P��<M|<�'8���3�o�At���p�[Ǣ��v�H��O��f��L�����'�|_B�H�W�1��30ՠ7�&��jQ�?ңڛ�zl�z� ��+A�M�/ӈ�@�4w$�ǐ�U�/�!G:�?H�3��{_@%�W=�Q] �F���DFO|ۡ�I�Yx(�����P�(��a�O�㌝�Z����v��_��TPÜ] *]G'��$�D�~�Ǽ9v�f�b��ڊ�QW&�@�@�0;l������l�(O���+���w�4�3�۔�կ��2n=�/[O�����|�5���$�I�P�j�z�ٵ]�{0ܘ���)��
��]؅q�k�Tj�,�1mL�"L>�ވ�|�������R���H:�})ieQ��W���3�����#PhR�!"�ξ@�s����Q?��흋*t�4֤��(��$�����8O�a�}�[��y���u_h�6W������:��m�*!o.6�n�����%���J=:��zZ�!���
F�I�$�Y�^)Y��t��E"?>�3t�s��:d�É�XF%-�G+����[Q�����/ty��ۄa�kJ'Ӻ��=�m��xi�.ͫ��H++d�䣅o���E+-���QQ�\�� ���Q���� vx�H�F��X��6_�����0��1�_���q
��9��� �~�*F8�'�0��B��k�.�U�k[*z�j��x��=�"�L��	$��gHX�7���^e�c#,���5��IO�����q���B@$��`Uy��4F��8����=�^e5Z�.�����:O���mi�Ƿ�AC�ɬ��dr�Xu&�D�����{ՃkSv�~0���>�b%��!Sn�it7!t��p�����͞���Z��w�������������K��mb��!���·Z�@��>�n��װLC��T���tJ��5���p��~�;A f�����V%�/�S��	D�ISdz���r�z=��x�������=5\�"U���p����<^)�KoBBz��р�k,5�@kH��R�K��_�c7��'�!;);����(!+D��+a0��TjMR��D�{W�J2X��������/hkL+ �+��]ڥ.�D&�᪁�x]�J��{���Ua��O�v�"
��dj������4��a�?Y�9��ۮ3��"h�x:7���$�M�f�sC���\���!�^�i�63-9�:�a���r�	t��jc���q7��Jn�z�&�~FĚ�ё'���Y7Ø�Lg$��U%�b:Q:�IQ�s�r.�?��t$��~�Pg�TG�v/6��+~$�E������ojMZdAɥ�>�q?��C�f?P"��H�ȱ.���|���yo91��(�H�M��OsTj�����&^C���S��1O :��*cn��;fr<�D�"%v�-���윒Yv���_��?��1���m��f1Џ=a�
����FP�>�����V�!ȱ

�����gĢ9x(�]��z������F�k�����C����$�H]m>�?��y�D�c�.�{ A�F,-#���Ð'��� }��w�Z���/1(��A�EDLs*���������2�e�
ٸD�t���b��S��3��v&�枥b<��\ξ�;h�$,�`�y��s�9�xvC�c�أ�-r�!��0E��7����S�5��$*H�n_%���ab��1�l�/z����t��C5I�^�����I��&���5cH������
�7%�f8���^	h�I���R�2ҧ��x�pI�AtͬU��rU%���򃾍�����C�^�V%�:��YA�ĩ9�Y$�]����)����-�5Bt��LLE)ā�\ow&��ͷko�9��5����X��)@aǾ��È�/'�3W��9��ҭeQ��
8pL�8�VE��Dc�ί���fx0I��Ҩ3��;��Hi"h�!��*JQ#g���֐�tsq��R�� ��x���N��m�T�B�'1����+����?b˝.��8��DV��Ivsw�%s
����t����I�B_qSʘ([��$����>͢��ۻV�EQ����/�|�uӊ�gq>�lXc���9�_��#��$�������L9���NQ�
=H]ՑTh�j�E\���"�^�,�H\(�lj���)����݄����^�˖�6Y�����k�}��	!r�\��:#�� i� ������#�(1q�b#o�$��;2u��0�R�{ץ>��'������V>ULRҒ*v+BS���Z?���Du�e�4��mL�r�����84��F���k���\!���<!G����H��,������?_��ïP��}������ �4�wC��4��������X��}�̓� �=�!.��Y4��5Ě���22�s*|Ѣ%s�W?of-��>��_�4���^��y�Qpa Z�$�0�~����y�k�Z]]�Z%�&�t����@#p,=>�R�m���s�v{�5s�f�yӪD�&���|R��_���LI��)ܾ�ry��8�<�Al���2�k|,�&Y�&����l��T�#7�����_�iP"��馷6�b9h��=\t�Q&r㊭�U%tx�HUM�!vD
=}�F!�3���8L��
#~f�ڗw���Fh ��w�V9�]�~Dh��U>1^g��Rl|g�c�ϖ�X�6b#`|WF�]��I�%�v�qT9���7¥��+�*��N%�`����Ŷ�Rh�ި�@�y\�g��8X��Y���D�	D_z2#���T�
v$I�Ȏw׫����2L���7�W�ƹ�0PX����g	O4 s����H����5q1D���wtr� �c�O��ꣶW5n�pt�9x�L!���:l^o��5�E���#"����Z�T@�H������.F1��C��=�j)e���c8�v&ơN�x���  t�r��Ӄ������	*2���<9��$y�tAP|k�Q2U��t�mRS��Ϳ����	o���`p3'�QB�i+����7��AW|VO6<�G�?;�h6Nk�d�r8TQR�~{(I9d�������핐Ut��;5s��u���͝�i��囇�MVϣvq�f�׋^�Q��&�T���F*��A�]�G���-O�5��d�0�Nk \D�	�]ۛ��T4�5��eP��+pZ|�!��j�]��;�G*�d?�u"v��nJ�(�j�N�C�0%9zXk�������z���)-�&�aUÚO�C�c�~��\f5�}�E�E�aA @�"�O��߭���F ��=5-p-��}~3���K�}�O�*�I��)@�ν��>�+���f}�t�`�������U�hs
5��#����ؽ�䜪�3�gt�����������}�����!%6���!L�v��db��.��1� �-�^��YȖ��'��C���j}ª��y�e�&�t�󙾁q���	�3m\ƸN4�t����CP>8�t�)�^�44���Mϫ�^Z�I�5Ώ��P4����c���)���Oox�1P����m��=���2�Kr���?D��p���z�IN�X�X�-�~�1ښ�b/{B�j��@PC V�/�pT�=�\S.K��>��iѢԸ��b��.e��q6������?��SZC�n˲��̺��*�E	z�����[? ���(�o���ұ{�)����>�Q���S�Bxx�>�|s�6�N��������*�e�h�.&D��
"���J�[<�"..49�r(�Fu�N9��5�d�:i3ڗ�yi&�ڳ�!�'�����d<�K�6�U�AH�Qy�A��F�����/�(cm$�V���5w�}z�l��	��/�<9"�2^��A��HE�^��ꃕ�$��[n�����Jw��e1�t��i�10�j����*�)m�W���	~[��F�C��M�����K�v���&�t�h�_X	�o,XJ���~��h4���oT�̻z��ݖ��1Գ�ܕ�#3�֮%�����6�>���/ h \�nO�W6�2v�v4�$��q���K��,;;񔮟�����#���|Mһ���Q {�V�ξ�!0�)xdo�I9�ۏzN�E#p�jy�x��jx��q<����q)�Ԡ��4�Z��2p����܆���}P#kJ!hbl5�-=J�(5N`����ͻ��~'r�@:�"���=��XΫN^����0�:k�Uo!	�s?`H7҆�Q��ޓ-E�;�Ɗ2���� �d"�+nc���_�`����gC��n�;ηeM�2�������]�*,L� j& �|����@|�p_��mX���y��s��=n���rePO�r�/~�P&�.<-!��{���~�	�d8���6�A����������y�b��m��if�Am��v��Y݃�� �.��3���|C
���|YCK�#q=T5!�O�&����Byk��v�e�y���c�C�T\_f�[�ެ�r�R
�')�+ P!��%b�ܗ�;�\+�f�m����ݡ���ӈF��*��a_�T�bA�vK�#�^��ft����w���mW9�(��IH���S�AF[^r)Z��9���a]�,ů�8)��7��|�:)��|5���Cb�2��q}�~s1b)2���W�D��������[C�T ���q�5	�ūI	y�'S��v�W��E���X��)�W(��7�hO2�:s �g7k�ܺ��qg]����^r.�����t���j�G�PR��u�)\uĕ�!���%1�����d�E��cf�����/�#Ѐ7��Mѓ:�#��h�&XJ&X6�w���oL���r�Y��	�#�o]�D�6y�XScrǩS��0+� />Fg
oC^q�� �6�Y|�1s�k�?CGR���o�g��`���!���H�������Y^��a�Q��jQ$WU=�����;wU�GCT	rV����S����(Ep���V%^X� :���)���	)=ᝏ�?*���l�Ķ������˧F�ɝ�OA�ٴ��,�kdR��T�J�VW'
��
vjd*(@�l��]Vi3#���;8��������m�0=L[e�Q|�`��j�o������(
���`,f�jgW���NR��s,Y�ǈ�>�'2��/���k/;��A>X�L�d��D�=�n�D��
T�z�i��8�7}ыr�Ncq�q����F`fC�����k�1�(���>>j�Rk@L�#��`>z
���!0�2NX~�d�<bim4]^��v� a���B�I�n�����ΐP$�'�=��CtM��j��Z\ʫ\M�rE�0���$%ݽ���uJ57�>�EM�Iׁ���1��?���#��I� �e�ƺ�%y�:��IJ�.$\��������/��Ri$$@.:9?Bm���e\%@�р�L�B�0��xBf/�����!�%-*����h��(:!��.3L�*չtҦGgWM������*�9t����|���N�|,&Ξ����Y���*,�s6W��Q^[�0>��<2�֊��޼��,��LD"�/��d��o������"}��M�-t'�Ҵrh����=��x�2��S�G�2 �/�&s9�EQ��뛍y��A�-
�TC��"���x���w;��F��ٴݓ�.2XW2��D�!�Q�LꚀ�H�a,9���mm*��9�o^�aED}�p�|���맡ɞ'��nxy&Ě�^6Ncywt���K���&�d�/ObK]_$�ykr��^������]���+(9`@0�kOx��W�Pls����p�޾��V��qB��T�3I�,�ڿ�0�f��6��Da�2�Oq5�_�nhi�
)�H�����&�Ǡ"��+�?�u��G4f_Vٰpj�/	�L���l�`rT��#�ߋ�^I�[P�o���Q�q�S^;w��5�ȟ[ǵ�崟z��/��X����D�`��@d�#w�t��UE�F�wGo4N!"������i\�N�X�ٗ�(\��_��`���?�n��>e�������z�U�	oa&���|qJ�wm(����� ~��ICk{�?_�,�����q`F���Wnx'X2��_V�`S�����}oٝ�y�l<_�h��p�v،"����l)^��Y��AN�'������	�g���˗���E�� yz�؎|��W�ufM��Q�N�x�y�A+��c��G��)
<���6���W�������	4��(1J�;]:&�i��Y(k�i�8��p��������i�8"��~c=$Y8�Ds�$R���Um+����N9����"�R��Cp�B�+z�<�Bz��0�j$A�H���H{g�Ң �P�c�,���q