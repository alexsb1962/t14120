��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�Ȱ���<�`��/�*r�L\�|��>��)�Z!�y��AVd�.�r����E��2��n/����a��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)����$�a<��d�6�q��tӏ�ˡ\s�$�L���Ÿ|^*��g�@U�*2�X���2��^�:9��D<��;�h��É}����a$;��몬g��>��W��iv���o�ăN�G\\�[�4�������W4xl��0�;O���V^��@��l5f+��\�&�7F�CqϮ�Y"�� C�T���/��Ƹg"���l ����~G�_y�kIe�+E�9�>Ǹ=�oWS�|���WV��P����������L��΋I2�G�r	y�i&�l��vЦ5�o�#����T�WrkV#��+�ڛ����C��ɀeG31>�����k�\�%�̶�@J�%A-�@�'2�}�0�΋ha���RN;zy�Q}N��5Z��}L���Z��¼�1<}M�����g�) $�8��Ρ�g���}E����G�@).�b���L��<�1�~:�~"�S��Y�p*-��^(Yj�����k��=98VK�ϲ�=�Zhy��� �#��_���c���~���YƯXrh"� Sao�%��Ƭ�;���cE��:�<:���6��E����Mr`2C���L�g.�T�"/)(dAX �B\\�xG�� ����	��r=�ى��x�⿐�z{�&��!�$�ȠC���}���?pEp�����p���р�e��Tu�M�@(���v6�ɥ.D�{(��Ķ)B0�h.ˢ�ا--��I�OtQ��I�ǧ�b:�ot����'�� �AvY��ɲ��c�Q��h�v�z�Fo�6$�ǧA��h�;�X��?F�4�E���j���X�Qd�i�� �C���¤T&=Ò�z#������z?��:�]q�����j.J�~�FH�/�ڽ@_)�f�&��[Ces�Aش�Wۛ���/�"��m���砼G� X��r糣@�mS�f^U*�x����{���3!<���5#	��[����X����7X�1
��r��;$�g���m�:$�,��CLXwcIp�RW��*���E
Y��5 �)��¯��W��)�]�'�n(k��ı����	�)�%��!b�{���!����,'Z�/�n/|pnf�O�F}ξX�^����6��e�RF�j�u�H�SS�蚺%���n�lV+��K9y�.}���؛5E�����W�h��o$C���p��`�y������%9��)�H���9H���pZ�����_�[�[d �[��;�DN�#K�X�5+��<�6TH�����f�Π�(xk�0�{"5h�B�_>��yʡ>C����6|�b��^X���)���
�����b���R�v9�Cxt�_rf�u��֛l,='ps$�2K��W2��>	gj"�#��yM-ێ�Ϛ��h%���h�h:Xx�<���!Ÿ�@I��������*�a�4��&>	�ւ�'��~�����I��E޿�?׊�&x:K�~���?�4�d�[A�#�����t��9.�v�|��}��?��F����ET����y�B&}K���.4���٠�fFJA	5g-O�fme��(/J�-�N[�A^��}��{�d�@�Y<�[�j��RY�U;���R�	?��.0�E��C'�߬$�(�ˏ��8�b�@yh>&�O��}����4"�X?&#	��Q�է*���<b�I}�^�@�w4��6w�$\}=���M ��X�f9���P������$ұ��Òs��0%��^SG1�� U���C�N�S���`�ژC9�D[u��hh�4����Uïm�M���O�����/
����޽	S�2^]��ŹN9�~���+�@˟�H�L	��E�i������Ac�$�.�u�s5cF�r�U�qB��M��mٻ�H Y�V�l��$��X�D[��f���U_�Ks;�Mi�����U< ӯp�(˞���a������x���f0w�rM���"*
�q�u�>�0�JL�ȍ���s�ގ:�*n��^���߄�����$��6n�N��y�'}0�n	������-J��F]$��1��{��l>��;BX�Iy��l��Ԗ��&��Ĳk�Ý���Ŝw
Z���hOy�Uɦ����-qC�_/Z���>��$Q�-I7�U�e��ܼ��
6c ������`�E�1�`�������QT��s���`d�7r�X���r�'y��G�����/M2�G�9cfX#��ܞ�1�T�����vQ��zy��.g�L�5��E4�����T�vθْ�~��<��V�LL�����/��	n��.�I�,�ׂ4`01����:^ӰcK��O��;��y��r0ݖ'�~=^;4v���k>�G0M�ۤV-���U��[�y�h�}NWm��r({��~ٗ�,��4�_]����z]�E���L4����Y��Gdl��A.~+�Cm���Xw��z�ݪ^
���.�qҗq��c�c4�� \R�
&k�5	����6)����i\�r�g������܇}����W	�|>/V�T�+^�F�T�f^�0+�~җeؑ`�� &���gq��9����im��Q�����x'(S�LH4S��O�߰�RP�2�I )��X	"j�L��^^"^ k��a�i���̦.��s�k�п
�ind��ځ�3�/u�����\�N�~�U��"�,:��JoG̅�	{��Zt���UC8]�p�G�50���N�S}��%���|_.����%5��:DsQS�ۨ��z�m�bY�O,��sc�a����\��y.7��@q���T��8����Ndդ�1E���҄�s?!��;�V���k'\�1~w��dͭ b����������2�������E�Wk�%��:����]K���2�QЯ�q����s�,������L�;	���U������Ԓte�\4�WȦ(9���TjR/Zh[Q�G��Ֆ*���s/��bR��	��⊸gV|���J/�A���\���{O��q��>b6E4����jl�ΐT k�q�頺���=>��AT������^���Y}���}��Y�1E�ט6 ��t��:���d���I�wE�~��U�īc*�&�j1D������[9D<�	��v�˶{����� ����b-��T�R d�-�#m�4@T}�ۧ�i��4#���m�?���[@`�ĥ��g�%DKsk�2��K�R����/{A��/V4�B���n/_&A��Z�bDE���L�CH�wl��v��Q�q��^e
�{�w�k{#d��7径�Jd�(M�CY%^���}e���2��(}�+��#�R�;�eͶ�� ��]UC��0V EK=�I��j�T��^� �o����2�xţI���]���n�^e'�mT[7g>+�:p;۱n��w���g��Nr�����Z�
u~�93nAS�VO0"�ynNʀ�����ה}&�ū�l��8}����G-*'2��*�ض�{��Rh�D<�";��`�KJ������Ms�T�[x-dL�>�
�ӴvR�t��8IǢ҃)�r[�*�)(˝��c����<�\�Ǽ4��X���������V�1�8��I����yLR�QR��?�ņ�vAv=׸FyD�{ō)��B�P[3����|z����f�ț���Ehמ������ǵ9�����m���o��ף��{o�9�y�s(VMg[�{�H1���Ăy�=ɜ�!-�xI����h�a��'�c}�������I̞�� ��a'��v0��(cl��շ�[�޲.8���e:�`xg��E�z�ད�sC�4�qdѩ0v��8�}2�p�zކݸ9��g�֖�/햤1���]YBa.:P��k�Gm�b�]�2`�K�ɉ�81*So�JjM��*���]��z������}QLA�[�Pg�(�$v
�'|����<\.(�:���K7�F�
@p3�!^�kc5�`��	-D�\(����O0�z�~S��������fN ��e"_�GQ��b�J� ����m�ު�b��,B��TI�S����� ��^�oB߇�t,ô<*�\���E���
��`�A%#�%�P���S�x��?�y<�,ZX�pB��fk��2Wg�I��"�F�L<�$�_1BH���2����L̎N��p�ju&-L;t���/#�I�]7,+��ă�0�| >iy��p�	n�k�l5I�0�d~��٭e���p��>��9�諐|�SU�(��<�z��Ćt�a"�=����U�e��49���{%O�Ip8����l�]��2V0�*�mІPf��eZ����#} �ژ�<�j<�'^��)����Me�ف�Ģ!6F�x���_�`�VӔ{M���1�T=Z��V͠�%�l l�P���]�G�=ʵ]_x1ǃkcO�'ԂI൨~F8:��[AB����'&��(ֱz�9�J�ҷ\"��3�� ��%N
�DA�+E�8�>vJK�0㫌��W� 
�:���oe������N����;��B&g�����7ҭ(��@�>b([���=HH��u��gc���v��sley�3�S�k.��(�Y�k�<�Ƣ�
�̞cB�Ze&�s�S��#�5x<�e�Y�gJP�oT��g���4�� ��އ�n\��_+���V:�֤rJ��� �_��	��5�h����?IH83��<� �����m7��n#��*5�쟃W�@)L�ʯ�wH�W�a����^����&_aJ�*2�݉e�oCچ��DJ�>2�ԏ��L���4ՠB�2�[�9�9A�6�g%{��mY�Bᗆ��S�a�kb���^-��SH�?"�ۼ�yfʸ��{�Ъ��."�����
��yr^�?�1r�,�U��Bd�v�4K��b�HW�q/cnۭ>��J�G�����t�*oV��t��oz�y��h^�}�k,��VD-H� ϏP���gF8mB�	�/@ӯ� ��^J��xÕ�Z������+)V.ޘ�	�S\�)�@2�(�����'�z������gY����3��wri*�v�JKl�e
7��kNB�3u[�v�& �t��8�f[��&�T䕤�n�\��4L�Bc��[�Ͳ����D:�v�XM��
~����Fz�������NUvP��f@j=�
����]��w�n�����=g-tS'ʠ-RM���04���"�-��!V�B��T5���&R� s:?�R�E#1�_�WD(���^s����n��d0��^+b�)�>��b�F�v����"� �夾([^�P�Z??O����pf�8��T��O8-����R��c ���2=>q��|�p\�`��_�̘�/Ibj6�G��V�$�
}�؏����g��������Z�v���XL9�Ȱ��`,�f8��oSB J��w-��­�1�>�J�蟚��ʉ������;}����3���lD"��t.f2�2tz��ݷ0�Q�d~����J�	��̭�O*/Msњ .OW^�,n���[_�Ijb��k\Y�R����X�?�h�r1}�;Y���ɇ(2A%������{�+綇�#���I�6��{�%��ύÊ�o�pQ���~��n{���)�V4�sEM2��Ď^�2�(2H�MJ������91�1/���5�+ۣ�]Lx��QJ$� ,Wmk�wSZ��>�$	�h��������0: